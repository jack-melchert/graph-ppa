// Module `global_controller` defined externally
module tile_en_unq1 (
    input [26:0] I,
    output [0:0] O
);
assign O = I[26:26];
endmodule

module tile_en (
    input [0:0] I,
    output [0:0] O
);
assign O = I;
endmodule

module rf_write_sched_0_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module rf_write_sched_0_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module rf_write_sched_0_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module rf_write_sched_0_sched_addr_gen_starting_addr (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module rf_write_sched_0_enable (
    input [16:0] I,
    output [0:0] O
);
assign O = I[16:16];
endmodule

module rf_write_iter_0_ranges_2 (
    input [16:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module rf_write_iter_0_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module rf_write_iter_0_ranges_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module rf_write_iter_0_dimensionality (
    input [22:0] I,
    output [2:0] O
);
assign O = I[22:20];
endmodule

module rf_write_addr_0_strides_2 (
    input [22:0] I,
    output [4:0] O
);
assign O = I[19:15];
endmodule

module rf_write_addr_0_strides_1 (
    input [22:0] I,
    output [4:0] O
);
assign O = I[14:10];
endmodule

module rf_write_addr_0_strides_0 (
    input [22:0] I,
    output [4:0] O
);
assign O = I[9:5];
endmodule

module rf_write_addr_0_starting_addr (
    input [22:0] I,
    output [4:0] O
);
assign O = I[4:0];
endmodule

module rf_read_sched_0_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module rf_read_sched_0_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module rf_read_sched_0_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module rf_read_sched_0_sched_addr_gen_starting_addr (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module rf_read_sched_0_enable (
    input [16:0] I,
    output [0:0] O
);
assign O = I[16:16];
endmodule

module rf_read_iter_0_ranges_2 (
    input [16:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module rf_read_iter_0_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module rf_read_iter_0_ranges_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module rf_read_iter_0_dimensionality (
    input [23:0] I,
    output [2:0] O
);
assign O = I[23:21];
endmodule

module rf_read_addr_0_strides_2 (
    input [23:0] I,
    output [4:0] O
);
assign O = I[20:16];
endmodule

module rf_read_addr_0_strides_1 (
    input [23:0] I,
    output [4:0] O
);
assign O = I[15:11];
endmodule

module rf_read_addr_0_strides_0 (
    input [23:0] I,
    output [4:0] O
);
assign O = I[10:6];
endmodule

module rf_read_addr_0_starting_addr (
    input [23:0] I,
    output [4:0] O
);
assign O = I[5:1];
endmodule

module ps_en (
    input [0:0] I,
    output [0:0] O
);
assign O = I;
endmodule

module addr_gen_3_16 (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [1:0] mux_sel,
  input logic restart,
  input logic rst_n,
  input logic [15:0] starting_addr,
  input logic step,
  input logic [2:0] [15:0] strides,
  output logic [15:0] addr_out
);

logic [15:0] calc_addr;
logic [15:0] current_addr;
logic [15:0] strt_addr;
assign strt_addr = starting_addr;
assign addr_out = calc_addr;
assign calc_addr = strt_addr + current_addr;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    current_addr <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      current_addr <= 16'h0;
    end
    else if (step) begin
      if (restart) begin
        current_addr <= 16'h0;
      end
      else current_addr <= current_addr + strides[mux_sel];
    end
  end
end
endmodule   // addr_gen_3_16

module addr_gen_3_5 (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [1:0] mux_sel,
  input logic restart,
  input logic rst_n,
  input logic [4:0] starting_addr,
  input logic step,
  input logic [2:0] [4:0] strides,
  output logic [4:0] addr_out
);

logic [4:0] calc_addr;
logic [4:0] current_addr;
logic [4:0] strt_addr;
assign strt_addr = starting_addr;
assign addr_out = calc_addr;
assign calc_addr = strt_addr + current_addr;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    current_addr <= 5'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      current_addr <= 5'h0;
    end
    else if (step) begin
      if (restart) begin
        current_addr <= 5'h0;
      end
      else current_addr <= current_addr + strides[mux_sel];
    end
  end
end
endmodule   // addr_gen_3_5

module for_loop_3_16 #(
  parameter CONFIG_WIDTH = 5'h10,
  parameter ITERATOR_SUPPORT = 3'h3
)
(
  input logic clk,
  input logic clk_en,
  input logic [2:0] dimensionality,
  input logic flush,
  input logic [2:0] [15:0] ranges,
  input logic rst_n,
  input logic step,
  output logic [1:0] mux_sel_out,
  output logic restart
);

logic [2:0] clear;
logic [2:0][15:0] dim_counter;
logic done;
logic [2:0] inc;
logic [15:0] inced_cnt;
logic [2:0] max_value;
logic maxed_value;
logic [1:0] mux_sel;
assign mux_sel_out = mux_sel;
assign inced_cnt = dim_counter[mux_sel] + 16'h1;
assign maxed_value = (dim_counter[mux_sel] == ranges[mux_sel]) & inc[mux_sel];
always_comb begin
  mux_sel = 2'h0;
  done = 1'h0;
  if (~done) begin
    if ((~max_value[0]) & (dimensionality > 3'h0)) begin
      mux_sel = 2'h0;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[1]) & (dimensionality > 3'h1)) begin
      mux_sel = 2'h1;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[2]) & (dimensionality > 3'h2)) begin
      mux_sel = 2'h2;
      done = 1'h1;
    end
  end
end
always_comb begin
  clear[0] = 1'h0;
  if (((mux_sel > 2'h0) | (~done)) & step) begin
    clear[0] = 1'h1;
  end
end
always_comb begin
  inc[0] = 1'h0;
  if ((5'h0 == 5'h0) & step & (dimensionality > 3'h0)) begin
    inc[0] = 1'h1;
  end
  else if ((mux_sel == 2'h0) & step & (dimensionality > 3'h0)) begin
    inc[0] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[0] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[0] <= 16'h0;
    end
    else if (clear[0]) begin
      dim_counter[0] <= 16'h0;
    end
    else if (inc[0]) begin
      dim_counter[0] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[0] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[0] <= 1'h0;
    end
    else if (clear[0]) begin
      max_value[0] <= 1'h0;
    end
    else if (inc[0]) begin
      max_value[0] <= maxed_value;
    end
  end
end
always_comb begin
  clear[1] = 1'h0;
  if (((mux_sel > 2'h1) | (~done)) & step) begin
    clear[1] = 1'h1;
  end
end
always_comb begin
  inc[1] = 1'h0;
  if ((5'h1 == 5'h0) & step & (dimensionality > 3'h1)) begin
    inc[1] = 1'h1;
  end
  else if ((mux_sel == 2'h1) & step & (dimensionality > 3'h1)) begin
    inc[1] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[1] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[1] <= 16'h0;
    end
    else if (clear[1]) begin
      dim_counter[1] <= 16'h0;
    end
    else if (inc[1]) begin
      dim_counter[1] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[1] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[1] <= 1'h0;
    end
    else if (clear[1]) begin
      max_value[1] <= 1'h0;
    end
    else if (inc[1]) begin
      max_value[1] <= maxed_value;
    end
  end
end
always_comb begin
  clear[2] = 1'h0;
  if (((mux_sel > 2'h2) | (~done)) & step) begin
    clear[2] = 1'h1;
  end
end
always_comb begin
  inc[2] = 1'h0;
  if ((5'h2 == 5'h0) & step & (dimensionality > 3'h2)) begin
    inc[2] = 1'h1;
  end
  else if ((mux_sel == 2'h2) & step & (dimensionality > 3'h2)) begin
    inc[2] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[2] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[2] <= 16'h0;
    end
    else if (clear[2]) begin
      dim_counter[2] <= 16'h0;
    end
    else if (inc[2]) begin
      dim_counter[2] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[2] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[2] <= 1'h0;
    end
    else if (clear[2]) begin
      max_value[2] <= 1'h0;
    end
    else if (inc[2]) begin
      max_value[2] <= maxed_value;
    end
  end
end
assign restart = step & (~done);
endmodule   // for_loop_3_16

module pond (
  input logic clk,
  input logic clk_en,
  input logic [7:0] config_addr_in,
  input logic [31:0] config_data_in,
  input logic config_en,
  input logic config_read,
  input logic config_write,
  input logic [0:0] [15:0] data_in_pond,
  input logic flush,
  input logic [4:0] rf_read_addr_0_starting_addr,
  input logic [2:0] [4:0] rf_read_addr_0_strides,
  input logic [2:0] rf_read_iter_0_dimensionality,
  input logic [2:0] [15:0] rf_read_iter_0_ranges,
  input logic rf_read_sched_0_enable,
  input logic [15:0] rf_read_sched_0_sched_addr_gen_starting_addr,
  input logic [2:0] [15:0] rf_read_sched_0_sched_addr_gen_strides,
  input logic [4:0] rf_write_addr_0_starting_addr,
  input logic [2:0] [4:0] rf_write_addr_0_strides,
  input logic [2:0] rf_write_iter_0_dimensionality,
  input logic [2:0] [15:0] rf_write_iter_0_ranges,
  input logic rf_write_sched_0_enable,
  input logic [15:0] rf_write_sched_0_sched_addr_gen_starting_addr,
  input logic [2:0] [15:0] rf_write_sched_0_sched_addr_gen_strides,
  input logic rst_n,
  input logic tile_en,
  output logic [0:0] [31:0] config_data_out,
  output logic [0:0] [15:0] data_out_pond,
  output logic valid_out_pond
);

logic cfg_seq_clk;
logic [15:0] config_data_in_shrt;
logic [0:0][15:0] config_data_out_shrt;
logic config_seq_clk;
logic config_seq_clk_en;
logic [15:0] cycle_count;
logic gclk;
logic [4:0] mem_addr_cfg;
logic [0:0][15:0] mem_data_cfg;
logic [0:0][15:0] mem_data_in;
logic [0:0][15:0] mem_data_out;
logic [0:0][4:0] mem_read_addr;
logic [0:0][4:0] mem_write_addr;
logic read;
logic [0:0][4:0] read_addr;
logic rf_clk;
logic [4:0] rf_read_addr_0_addr_out;
logic rf_read_addr_0_clk;
logic rf_read_iter_0_clk;
logic [1:0] rf_read_iter_0_mux_sel_out;
logic rf_read_iter_0_restart;
logic rf_read_sched_0_clk;
logic rf_read_sched_0_valid_output;
logic [4:0] rf_write_addr_0_addr_out;
logic rf_write_addr_0_clk;
logic rf_write_iter_0_clk;
logic [1:0] rf_write_iter_0_mux_sel_out;
logic rf_write_iter_0_restart;
logic rf_write_sched_0_clk;
logic rf_write_sched_0_valid_output;
logic [0:0][15:0] s_mem_data_in;
logic [0:0][4:0] s_mem_read_addr;
logic [0:0][4:0] s_mem_write_addr;
logic t_read;
logic t_write;
logic write;
logic [0:0][4:0] write_addr;
logic write_rf;
assign gclk = clk & tile_en;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    cycle_count <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      cycle_count <= 16'h0;
    end
    else if (1'h1) begin
      cycle_count <= cycle_count + 16'h1;
    end
  end
end
assign data_out_pond[0] = mem_data_out[0];
assign valid_out_pond = t_read;
assign rf_write_iter_0_clk = gclk;
assign rf_write_addr_0_clk = gclk;
assign write_addr[0] = rf_write_addr_0_addr_out;
assign rf_write_sched_0_clk = gclk;
assign t_write = rf_write_sched_0_valid_output;
assign rf_read_iter_0_clk = gclk;
assign rf_read_addr_0_clk = gclk;
assign read_addr[0] = rf_read_addr_0_addr_out;
assign rf_read_sched_0_clk = gclk;
assign t_read = rf_read_sched_0_valid_output;
assign write = |t_write;
assign mem_write_addr[0] = s_mem_write_addr[0];
assign mem_data_in[0] = s_mem_data_in[0];
assign read = |t_read;
assign mem_read_addr[0] = s_mem_read_addr[0];
assign config_data_in_shrt = config_data_in[15:0];
assign config_data_out[0] = 32'(config_data_out_shrt[0]);
assign cfg_seq_clk = gclk;
assign config_seq_clk = cfg_seq_clk;
assign config_seq_clk_en = clk_en | (|config_en);
assign rf_clk = gclk;
assign write_rf = (|config_en) ? config_write: write;
assign s_mem_data_in[0] = (|config_en) ? mem_data_cfg: data_in_pond[0];
assign s_mem_write_addr[0] = (|config_en) ? mem_addr_cfg: write_addr[0];
assign s_mem_read_addr[0] = (|config_en) ? mem_addr_cfg: read_addr[0];
for_loop_3_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(3'h3))
rf_write_iter_0 (
  .clk(rf_write_iter_0_clk),
  .clk_en(clk_en),
  .dimensionality(rf_write_iter_0_dimensionality),
  .flush(flush),
  .ranges(rf_write_iter_0_ranges),
  .rst_n(rst_n),
  .step(t_write),
  .mux_sel_out(rf_write_iter_0_mux_sel_out),
  .restart(rf_write_iter_0_restart)
);

addr_gen_3_5 rf_write_addr_0 (
  .clk(rf_write_addr_0_clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(rf_write_iter_0_mux_sel_out),
  .restart(rf_write_iter_0_restart),
  .rst_n(rst_n),
  .starting_addr(rf_write_addr_0_starting_addr),
  .step(t_write),
  .strides(rf_write_addr_0_strides),
  .addr_out(rf_write_addr_0_addr_out)
);

sched_gen_3_16 rf_write_sched_0 (
  .clk(rf_write_sched_0_clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(rf_write_sched_0_enable),
  .finished(rf_write_iter_0_restart),
  .flush(flush),
  .mux_sel(rf_write_iter_0_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(rf_write_sched_0_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(rf_write_sched_0_sched_addr_gen_strides),
  .valid_output(rf_write_sched_0_valid_output)
);

for_loop_3_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(3'h3))
rf_read_iter_0 (
  .clk(rf_read_iter_0_clk),
  .clk_en(clk_en),
  .dimensionality(rf_read_iter_0_dimensionality),
  .flush(flush),
  .ranges(rf_read_iter_0_ranges),
  .rst_n(rst_n),
  .step(t_read),
  .mux_sel_out(rf_read_iter_0_mux_sel_out),
  .restart(rf_read_iter_0_restart)
);

addr_gen_3_5 rf_read_addr_0 (
  .clk(rf_read_addr_0_clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(rf_read_iter_0_mux_sel_out),
  .restart(rf_read_iter_0_restart),
  .rst_n(rst_n),
  .starting_addr(rf_read_addr_0_starting_addr),
  .step(t_read),
  .strides(rf_read_addr_0_strides),
  .addr_out(rf_read_addr_0_addr_out)
);

sched_gen_3_16 rf_read_sched_0 (
  .clk(rf_read_sched_0_clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(rf_read_sched_0_enable),
  .finished(rf_read_iter_0_restart),
  .flush(flush),
  .mux_sel(rf_read_iter_0_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(rf_read_sched_0_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(rf_read_sched_0_sched_addr_gen_strides),
  .valid_output(rf_read_sched_0_valid_output)
);

storage_config_seq config_seq (
  .clk(config_seq_clk),
  .clk_en(config_seq_clk_en),
  .config_addr_in(config_addr_in),
  .config_data_in(config_data_in_shrt),
  .config_en(config_en),
  .config_rd(config_read),
  .config_wr(config_write),
  .flush(flush),
  .rd_data_stg(mem_data_out),
  .rst_n(rst_n),
  .addr_out(mem_addr_cfg),
  .rd_data_out(config_data_out_shrt),
  .wr_data(mem_data_cfg)
);

register_file rf (
  .clk(rf_clk),
  .clk_en(clk_en),
  .data_in(mem_data_in),
  .flush(flush),
  .rd_addr(mem_read_addr[0]),
  .rst_n(rst_n),
  .wen(write_rf),
  .wr_addr(mem_write_addr[0]),
  .data_out(mem_data_out)
);

endmodule   // pond

module pond_W (
  input logic clk,
  input logic clk_en,
  input logic [7:0] config_addr_in,
  input logic [31:0] config_data_in,
  input logic config_en,
  input logic config_read,
  input logic config_write,
  input logic [0:0] [15:0] data_in_pond,
  input logic flush,
  input logic [4:0] rf_read_addr_0_starting_addr,
  input logic [4:0] rf_read_addr_0_strides_0,
  input logic [4:0] rf_read_addr_0_strides_1,
  input logic [4:0] rf_read_addr_0_strides_2,
  input logic [2:0] rf_read_iter_0_dimensionality,
  input logic [15:0] rf_read_iter_0_ranges_0,
  input logic [15:0] rf_read_iter_0_ranges_1,
  input logic [15:0] rf_read_iter_0_ranges_2,
  input logic rf_read_sched_0_enable,
  input logic [15:0] rf_read_sched_0_sched_addr_gen_starting_addr,
  input logic [15:0] rf_read_sched_0_sched_addr_gen_strides_0,
  input logic [15:0] rf_read_sched_0_sched_addr_gen_strides_1,
  input logic [15:0] rf_read_sched_0_sched_addr_gen_strides_2,
  input logic [4:0] rf_write_addr_0_starting_addr,
  input logic [4:0] rf_write_addr_0_strides_0,
  input logic [4:0] rf_write_addr_0_strides_1,
  input logic [4:0] rf_write_addr_0_strides_2,
  input logic [2:0] rf_write_iter_0_dimensionality,
  input logic [15:0] rf_write_iter_0_ranges_0,
  input logic [15:0] rf_write_iter_0_ranges_1,
  input logic [15:0] rf_write_iter_0_ranges_2,
  input logic rf_write_sched_0_enable,
  input logic [15:0] rf_write_sched_0_sched_addr_gen_starting_addr,
  input logic [15:0] rf_write_sched_0_sched_addr_gen_strides_0,
  input logic [15:0] rf_write_sched_0_sched_addr_gen_strides_1,
  input logic [15:0] rf_write_sched_0_sched_addr_gen_strides_2,
  input logic rst_n,
  input logic tile_en,
  output logic [0:0] [31:0] config_data_out,
  output logic [0:0] [15:0] data_out_pond,
  output logic valid_out_pond
);

logic [2:0][4:0] pond_rf_read_addr_0_strides;
logic [2:0][15:0] pond_rf_read_iter_0_ranges;
logic [2:0][15:0] pond_rf_read_sched_0_sched_addr_gen_strides;
logic [2:0][4:0] pond_rf_write_addr_0_strides;
logic [2:0][15:0] pond_rf_write_iter_0_ranges;
logic [2:0][15:0] pond_rf_write_sched_0_sched_addr_gen_strides;
assign pond_rf_read_addr_0_strides[0] = rf_read_addr_0_strides_0;
assign pond_rf_read_addr_0_strides[1] = rf_read_addr_0_strides_1;
assign pond_rf_read_addr_0_strides[2] = rf_read_addr_0_strides_2;
assign pond_rf_read_iter_0_ranges[0] = rf_read_iter_0_ranges_0;
assign pond_rf_read_iter_0_ranges[1] = rf_read_iter_0_ranges_1;
assign pond_rf_read_iter_0_ranges[2] = rf_read_iter_0_ranges_2;
assign pond_rf_read_sched_0_sched_addr_gen_strides[0] = rf_read_sched_0_sched_addr_gen_strides_0;
assign pond_rf_read_sched_0_sched_addr_gen_strides[1] = rf_read_sched_0_sched_addr_gen_strides_1;
assign pond_rf_read_sched_0_sched_addr_gen_strides[2] = rf_read_sched_0_sched_addr_gen_strides_2;
assign pond_rf_write_addr_0_strides[0] = rf_write_addr_0_strides_0;
assign pond_rf_write_addr_0_strides[1] = rf_write_addr_0_strides_1;
assign pond_rf_write_addr_0_strides[2] = rf_write_addr_0_strides_2;
assign pond_rf_write_iter_0_ranges[0] = rf_write_iter_0_ranges_0;
assign pond_rf_write_iter_0_ranges[1] = rf_write_iter_0_ranges_1;
assign pond_rf_write_iter_0_ranges[2] = rf_write_iter_0_ranges_2;
assign pond_rf_write_sched_0_sched_addr_gen_strides[0] = rf_write_sched_0_sched_addr_gen_strides_0;
assign pond_rf_write_sched_0_sched_addr_gen_strides[1] = rf_write_sched_0_sched_addr_gen_strides_1;
assign pond_rf_write_sched_0_sched_addr_gen_strides[2] = rf_write_sched_0_sched_addr_gen_strides_2;
pond pond (
  .clk(clk),
  .clk_en(clk_en),
  .config_addr_in(config_addr_in),
  .config_data_in(config_data_in),
  .config_en(config_en),
  .config_read(config_read),
  .config_write(config_write),
  .data_in_pond(data_in_pond),
  .flush(flush),
  .rf_read_addr_0_starting_addr(rf_read_addr_0_starting_addr),
  .rf_read_addr_0_strides(pond_rf_read_addr_0_strides),
  .rf_read_iter_0_dimensionality(rf_read_iter_0_dimensionality),
  .rf_read_iter_0_ranges(pond_rf_read_iter_0_ranges),
  .rf_read_sched_0_enable(rf_read_sched_0_enable),
  .rf_read_sched_0_sched_addr_gen_starting_addr(rf_read_sched_0_sched_addr_gen_starting_addr),
  .rf_read_sched_0_sched_addr_gen_strides(pond_rf_read_sched_0_sched_addr_gen_strides),
  .rf_write_addr_0_starting_addr(rf_write_addr_0_starting_addr),
  .rf_write_addr_0_strides(pond_rf_write_addr_0_strides),
  .rf_write_iter_0_dimensionality(rf_write_iter_0_dimensionality),
  .rf_write_iter_0_ranges(pond_rf_write_iter_0_ranges),
  .rf_write_sched_0_enable(rf_write_sched_0_enable),
  .rf_write_sched_0_sched_addr_gen_starting_addr(rf_write_sched_0_sched_addr_gen_starting_addr),
  .rf_write_sched_0_sched_addr_gen_strides(pond_rf_write_sched_0_sched_addr_gen_strides),
  .rst_n(rst_n),
  .tile_en(tile_en),
  .config_data_out(config_data_out),
  .data_out_pond(data_out_pond),
  .valid_out_pond(valid_out_pond)
);

endmodule   // pond_W

module register_file (
  input logic clk,
  input logic clk_en,
  input logic [0:0] [15:0] data_in,
  input logic flush,
  input logic [4:0] rd_addr,
  input logic rst_n,
  input logic wen,
  input logic [4:0] wr_addr,
  output logic [0:0] [15:0] data_out
);

logic [31:0][0:0][15:0] data_array;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    data_array <= 512'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      data_array <= 512'h0;
    end
    else if (wen) begin
      data_array[wr_addr] <= data_in;
    end
  end
end
always_comb begin
  data_out = data_array[rd_addr];
end
endmodule   // register_file

module sched_gen_3_16 (
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic enable,
  input logic finished,
  input logic flush,
  input logic [1:0] mux_sel,
  input logic rst_n,
  input logic [15:0] sched_addr_gen_starting_addr,
  input logic [2:0] [15:0] sched_addr_gen_strides,
  output logic valid_output
);

logic [15:0] addr_out;
logic valid_gate;
logic valid_gate_inv;
logic valid_out;
assign valid_gate = ~valid_gate_inv;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    valid_gate_inv <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      valid_gate_inv <= 1'h0;
    end
    else if (finished) begin
      valid_gate_inv <= 1'h1;
    end
  end
end
always_comb begin
  valid_out = (cycle_count == addr_out) & valid_gate & enable;
end
always_comb begin
  valid_output = valid_out;
end
addr_gen_3_16 sched_addr_gen (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(mux_sel),
  .restart(1'h0),
  .rst_n(rst_n),
  .starting_addr(sched_addr_gen_starting_addr),
  .step(valid_out),
  .strides(sched_addr_gen_strides),
  .addr_out(addr_out)
);

endmodule   // sched_gen_3_16

module storage_config_seq (
  input logic clk,
  input logic clk_en,
  input logic [7:0] config_addr_in,
  input logic [15:0] config_data_in,
  input logic config_en,
  input logic config_rd,
  input logic config_wr,
  input logic flush,
  input logic [0:0][0:0] [15:0] rd_data_stg,
  input logic rst_n,
  output logic [4:0] addr_out,
  output logic [0:0] [15:0] rd_data_out,
  output logic ren_out,
  output logic wen_out,
  output logic [0:0] [15:0] wr_data
);

assign addr_out = config_addr_in[4:0];
assign wr_data[0] = config_data_in;
assign rd_data_out[0] = rd_data_stg[0];
assign wen_out = config_wr;
assign ren_out = config_rd;
endmodule   // storage_config_seq


module mux_aoi_const_20_16 ( 
	input logic  [15 : 0] I0, 
	input logic  [15 : 0] I1, 
	input logic  [15 : 0] I2, 
	input logic  [15 : 0] I3, 
	input logic  [15 : 0] I4, 
	input logic  [15 : 0] I5, 
	input logic  [15 : 0] I6, 
	input logic  [15 : 0] I7, 
	input logic  [15 : 0] I8, 
	input logic  [15 : 0] I9, 
	input logic  [15 : 0] I10, 
	input logic  [15 : 0] I11, 
	input logic  [15 : 0] I12, 
	input logic  [15 : 0] I13, 
	input logic  [15 : 0] I14, 
	input logic  [15 : 0] I15, 
	input logic  [15 : 0] I16, 
	input logic  [15 : 0] I17, 
	input logic  [15 : 0] I18, 
	input logic  [15 : 0] I19, 
	input logic  [4 : 0] S ,
	output logic [15 : 0] O); 

	logic  [31 : 0] out_sel;
	logic  [15 : 0] O_int0;
	logic  [15 : 0] O_int1;
	logic  [15 : 0] O_int2;
	logic  [15 : 0] O_int3;
	logic  [15 : 0] O_int4;
	logic  [15 : 0] O_int5;
	logic  [15 : 0] O_int6;
	logic  [15 : 0] O_int7;
	logic  [15 : 0] O_int8;
	logic  [15 : 0] O_int9;
	logic  [15 : 0] O_int10;

precoder_16_20 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_16_20 u_mux_logic ( 
	.I0 (I0),
	.I1 (I1),
	.I2 (I2),
	.I3 (I3),
	.I4 (I4),
	.I5 (I5),
	.I6 (I6),
	.I7 (I7),
	.I8 (I8),
	.I9 (I9),
	.I10 (I10),
	.I11 (I11),
	.I12 (I12),
	.I13 (I13),
	.I14 (I14),
	.I15 (I15),
	.I16 (I16),
	.I17 (I17),
	.I18 (I18),
	.I19 (I19),
	.out_sel(out_sel), 
	.O0(O_int0), 
	.O1(O_int1), 
	.O2(O_int2), 
	.O3(O_int3), 
	.O4(O_int4), 
	.O5(O_int5), 
	.O6(O_int6), 
	.O7(O_int7), 
	.O8(O_int8), 
	.O9(O_int9), 
	.O10(O_int10)); 
	assign O = (  	O_int0 | 	O_int1 | 	O_int2 | 	O_int3 | 	O_int4 | 	O_int5 | 	O_int6 | 	O_int7 | 	O_int8 | 	O_int9 | 	O_int10 	); 

endmodule 

module precoder_16_20 (
	input logic  [4 : 0] S ,
	output logic  [31 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		5'd0    :   out_sel = 32'b00000000000000000000000000000001;
		5'd1    :   out_sel = 32'b00000000000000000000000000000010;
		5'd2    :   out_sel = 32'b00000000000000000000000000000100;
		5'd3    :   out_sel = 32'b00000000000000000000000000001000;
		5'd4    :   out_sel = 32'b00000000000000000000000000010000;
		5'd5    :   out_sel = 32'b00000000000000000000000000100000;
		5'd6    :   out_sel = 32'b00000000000000000000000001000000;
		5'd7    :   out_sel = 32'b00000000000000000000000010000000;
		5'd8    :   out_sel = 32'b00000000000000000000000100000000;
		5'd9    :   out_sel = 32'b00000000000000000000001000000000;
		5'd10    :   out_sel = 32'b00000000000000000000010000000000;
		5'd11    :   out_sel = 32'b00000000000000000000100000000000;
		5'd12    :   out_sel = 32'b00000000000000000001000000000000;
		5'd13    :   out_sel = 32'b00000000000000000010000000000000;
		5'd14    :   out_sel = 32'b00000000000000000100000000000000;
		5'd15    :   out_sel = 32'b00000000000000001000000000000000;
		5'd16    :   out_sel = 32'b00000000000000010000000000000000;
		5'd17    :   out_sel = 32'b00000000000000100000000000000000;
		5'd18    :   out_sel = 32'b00000000000001000000000000000000;
		5'd19    :   out_sel = 32'b00000000000010000000000000000000;
		5'd20    :   out_sel = 32'b00000000000100000000000000000000;
		default :   out_sel = 32'b0;
	endcase 
end 

endmodule 

module mux_logic_16_20 ( 
	input logic  [31 : 0] out_sel,
	input logic  [15 : 0] I0, 
	input logic  [15 : 0] I1, 
	input logic  [15 : 0] I2, 
	input logic  [15 : 0] I3, 
	input logic  [15 : 0] I4, 
	input logic  [15 : 0] I5, 
	input logic  [15 : 0] I6, 
	input logic  [15 : 0] I7, 
	input logic  [15 : 0] I8, 
	input logic  [15 : 0] I9, 
	input logic  [15 : 0] I10, 
	input logic  [15 : 0] I11, 
	input logic  [15 : 0] I12, 
	input logic  [15 : 0] I13, 
	input logic  [15 : 0] I14, 
	input logic  [15 : 0] I15, 
	input logic  [15 : 0] I16, 
	input logic  [15 : 0] I17, 
	input logic  [15 : 0] I18, 
	input logic  [15 : 0] I19, 
	output logic  [15 : 0] O0, 
	output logic  [15 : 0] O1, 
	output logic  [15 : 0] O2, 
	output logic  [15 : 0] O3, 
	output logic  [15 : 0] O4, 
	output logic  [15 : 0] O5, 
	output logic  [15 : 0] O6, 
	output logic  [15 : 0] O7, 
	output logic  [15 : 0] O8, 
	output logic  [15 : 0] O9, 
	output logic  [15 : 0] O10); 
	SC7P5T_AO22X0P5_SSC14R inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_0 ( 
	.A1(out_sel[2]), 
	.A2(I2[0]), 
	.B1(out_sel[3]), 
	.B2(I3[0]), 
	.Z(O1[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_2_0 ( 
	.A1(out_sel[4]), 
	.A2(I4[0]), 
	.B1(out_sel[5]), 
	.B2(I5[0]), 
	.Z(O2[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_3_0 ( 
	.A1(out_sel[6]), 
	.A2(I6[0]), 
	.B1(out_sel[7]), 
	.B2(I7[0]), 
	.Z(O3[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_4_0 ( 
	.A1(out_sel[8]), 
	.A2(I8[0]), 
	.B1(out_sel[9]), 
	.B2(I9[0]), 
	.Z(O4[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_5_0 ( 
	.A1(out_sel[10]), 
	.A2(I10[0]), 
	.B1(out_sel[11]), 
	.B2(I11[0]), 
	.Z(O5[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_6_0 ( 
	.A1(out_sel[12]), 
	.A2(I12[0]), 
	.B1(out_sel[13]), 
	.B2(I13[0]), 
	.Z(O6[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_7_0 ( 
	.A1(out_sel[14]), 
	.A2(I14[0]), 
	.B1(out_sel[15]), 
	.B2(I15[0]), 
	.Z(O7[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_8_0 ( 
	.A1(out_sel[16]), 
	.A2(I16[0]), 
	.B1(out_sel[17]), 
	.B2(I17[0]), 
	.Z(O8[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_9_0 ( 
	.A1(out_sel[18]), 
	.A2(I18[0]), 
	.B1(out_sel[19]), 
	.B2(I19[0]), 
	.Z(O9[0])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_0 ( 
	.A(out_sel[20]), 
	.B(1'b0), 
	.Z(O10[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_1 ( 
	.A1(out_sel[0]), 
	.A2(I0[1]), 
	.B1(out_sel[1]), 
	.B2(I1[1]), 
	.Z(O0[1])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_1 ( 
	.A1(out_sel[2]), 
	.A2(I2[1]), 
	.B1(out_sel[3]), 
	.B2(I3[1]), 
	.Z(O1[1])); 
	SC7P5T_AO22X0P5_SSC14R inst_2_1 ( 
	.A1(out_sel[4]), 
	.A2(I4[1]), 
	.B1(out_sel[5]), 
	.B2(I5[1]), 
	.Z(O2[1])); 
	SC7P5T_AO22X0P5_SSC14R inst_3_1 ( 
	.A1(out_sel[6]), 
	.A2(I6[1]), 
	.B1(out_sel[7]), 
	.B2(I7[1]), 
	.Z(O3[1])); 
	SC7P5T_AO22X0P5_SSC14R inst_4_1 ( 
	.A1(out_sel[8]), 
	.A2(I8[1]), 
	.B1(out_sel[9]), 
	.B2(I9[1]), 
	.Z(O4[1])); 
	SC7P5T_AO22X0P5_SSC14R inst_5_1 ( 
	.A1(out_sel[10]), 
	.A2(I10[1]), 
	.B1(out_sel[11]), 
	.B2(I11[1]), 
	.Z(O5[1])); 
	SC7P5T_AO22X0P5_SSC14R inst_6_1 ( 
	.A1(out_sel[12]), 
	.A2(I12[1]), 
	.B1(out_sel[13]), 
	.B2(I13[1]), 
	.Z(O6[1])); 
	SC7P5T_AO22X0P5_SSC14R inst_7_1 ( 
	.A1(out_sel[14]), 
	.A2(I14[1]), 
	.B1(out_sel[15]), 
	.B2(I15[1]), 
	.Z(O7[1])); 
	SC7P5T_AO22X0P5_SSC14R inst_8_1 ( 
	.A1(out_sel[16]), 
	.A2(I16[1]), 
	.B1(out_sel[17]), 
	.B2(I17[1]), 
	.Z(O8[1])); 
	SC7P5T_AO22X0P5_SSC14R inst_9_1 ( 
	.A1(out_sel[18]), 
	.A2(I18[1]), 
	.B1(out_sel[19]), 
	.B2(I19[1]), 
	.Z(O9[1])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_1 ( 
	.A(out_sel[20]), 
	.B(1'b0), 
	.Z(O10[1])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_2 ( 
	.A1(out_sel[0]), 
	.A2(I0[2]), 
	.B1(out_sel[1]), 
	.B2(I1[2]), 
	.Z(O0[2])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_2 ( 
	.A1(out_sel[2]), 
	.A2(I2[2]), 
	.B1(out_sel[3]), 
	.B2(I3[2]), 
	.Z(O1[2])); 
	SC7P5T_AO22X0P5_SSC14R inst_2_2 ( 
	.A1(out_sel[4]), 
	.A2(I4[2]), 
	.B1(out_sel[5]), 
	.B2(I5[2]), 
	.Z(O2[2])); 
	SC7P5T_AO22X0P5_SSC14R inst_3_2 ( 
	.A1(out_sel[6]), 
	.A2(I6[2]), 
	.B1(out_sel[7]), 
	.B2(I7[2]), 
	.Z(O3[2])); 
	SC7P5T_AO22X0P5_SSC14R inst_4_2 ( 
	.A1(out_sel[8]), 
	.A2(I8[2]), 
	.B1(out_sel[9]), 
	.B2(I9[2]), 
	.Z(O4[2])); 
	SC7P5T_AO22X0P5_SSC14R inst_5_2 ( 
	.A1(out_sel[10]), 
	.A2(I10[2]), 
	.B1(out_sel[11]), 
	.B2(I11[2]), 
	.Z(O5[2])); 
	SC7P5T_AO22X0P5_SSC14R inst_6_2 ( 
	.A1(out_sel[12]), 
	.A2(I12[2]), 
	.B1(out_sel[13]), 
	.B2(I13[2]), 
	.Z(O6[2])); 
	SC7P5T_AO22X0P5_SSC14R inst_7_2 ( 
	.A1(out_sel[14]), 
	.A2(I14[2]), 
	.B1(out_sel[15]), 
	.B2(I15[2]), 
	.Z(O7[2])); 
	SC7P5T_AO22X0P5_SSC14R inst_8_2 ( 
	.A1(out_sel[16]), 
	.A2(I16[2]), 
	.B1(out_sel[17]), 
	.B2(I17[2]), 
	.Z(O8[2])); 
	SC7P5T_AO22X0P5_SSC14R inst_9_2 ( 
	.A1(out_sel[18]), 
	.A2(I18[2]), 
	.B1(out_sel[19]), 
	.B2(I19[2]), 
	.Z(O9[2])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_2 ( 
	.A(out_sel[20]), 
	.B(1'b0), 
	.Z(O10[2])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_3 ( 
	.A1(out_sel[0]), 
	.A2(I0[3]), 
	.B1(out_sel[1]), 
	.B2(I1[3]), 
	.Z(O0[3])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_3 ( 
	.A1(out_sel[2]), 
	.A2(I2[3]), 
	.B1(out_sel[3]), 
	.B2(I3[3]), 
	.Z(O1[3])); 
	SC7P5T_AO22X0P5_SSC14R inst_2_3 ( 
	.A1(out_sel[4]), 
	.A2(I4[3]), 
	.B1(out_sel[5]), 
	.B2(I5[3]), 
	.Z(O2[3])); 
	SC7P5T_AO22X0P5_SSC14R inst_3_3 ( 
	.A1(out_sel[6]), 
	.A2(I6[3]), 
	.B1(out_sel[7]), 
	.B2(I7[3]), 
	.Z(O3[3])); 
	SC7P5T_AO22X0P5_SSC14R inst_4_3 ( 
	.A1(out_sel[8]), 
	.A2(I8[3]), 
	.B1(out_sel[9]), 
	.B2(I9[3]), 
	.Z(O4[3])); 
	SC7P5T_AO22X0P5_SSC14R inst_5_3 ( 
	.A1(out_sel[10]), 
	.A2(I10[3]), 
	.B1(out_sel[11]), 
	.B2(I11[3]), 
	.Z(O5[3])); 
	SC7P5T_AO22X0P5_SSC14R inst_6_3 ( 
	.A1(out_sel[12]), 
	.A2(I12[3]), 
	.B1(out_sel[13]), 
	.B2(I13[3]), 
	.Z(O6[3])); 
	SC7P5T_AO22X0P5_SSC14R inst_7_3 ( 
	.A1(out_sel[14]), 
	.A2(I14[3]), 
	.B1(out_sel[15]), 
	.B2(I15[3]), 
	.Z(O7[3])); 
	SC7P5T_AO22X0P5_SSC14R inst_8_3 ( 
	.A1(out_sel[16]), 
	.A2(I16[3]), 
	.B1(out_sel[17]), 
	.B2(I17[3]), 
	.Z(O8[3])); 
	SC7P5T_AO22X0P5_SSC14R inst_9_3 ( 
	.A1(out_sel[18]), 
	.A2(I18[3]), 
	.B1(out_sel[19]), 
	.B2(I19[3]), 
	.Z(O9[3])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_3 ( 
	.A(out_sel[20]), 
	.B(1'b0), 
	.Z(O10[3])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_4 ( 
	.A1(out_sel[0]), 
	.A2(I0[4]), 
	.B1(out_sel[1]), 
	.B2(I1[4]), 
	.Z(O0[4])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_4 ( 
	.A1(out_sel[2]), 
	.A2(I2[4]), 
	.B1(out_sel[3]), 
	.B2(I3[4]), 
	.Z(O1[4])); 
	SC7P5T_AO22X0P5_SSC14R inst_2_4 ( 
	.A1(out_sel[4]), 
	.A2(I4[4]), 
	.B1(out_sel[5]), 
	.B2(I5[4]), 
	.Z(O2[4])); 
	SC7P5T_AO22X0P5_SSC14R inst_3_4 ( 
	.A1(out_sel[6]), 
	.A2(I6[4]), 
	.B1(out_sel[7]), 
	.B2(I7[4]), 
	.Z(O3[4])); 
	SC7P5T_AO22X0P5_SSC14R inst_4_4 ( 
	.A1(out_sel[8]), 
	.A2(I8[4]), 
	.B1(out_sel[9]), 
	.B2(I9[4]), 
	.Z(O4[4])); 
	SC7P5T_AO22X0P5_SSC14R inst_5_4 ( 
	.A1(out_sel[10]), 
	.A2(I10[4]), 
	.B1(out_sel[11]), 
	.B2(I11[4]), 
	.Z(O5[4])); 
	SC7P5T_AO22X0P5_SSC14R inst_6_4 ( 
	.A1(out_sel[12]), 
	.A2(I12[4]), 
	.B1(out_sel[13]), 
	.B2(I13[4]), 
	.Z(O6[4])); 
	SC7P5T_AO22X0P5_SSC14R inst_7_4 ( 
	.A1(out_sel[14]), 
	.A2(I14[4]), 
	.B1(out_sel[15]), 
	.B2(I15[4]), 
	.Z(O7[4])); 
	SC7P5T_AO22X0P5_SSC14R inst_8_4 ( 
	.A1(out_sel[16]), 
	.A2(I16[4]), 
	.B1(out_sel[17]), 
	.B2(I17[4]), 
	.Z(O8[4])); 
	SC7P5T_AO22X0P5_SSC14R inst_9_4 ( 
	.A1(out_sel[18]), 
	.A2(I18[4]), 
	.B1(out_sel[19]), 
	.B2(I19[4]), 
	.Z(O9[4])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_4 ( 
	.A(out_sel[20]), 
	.B(1'b0), 
	.Z(O10[4])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_5 ( 
	.A1(out_sel[0]), 
	.A2(I0[5]), 
	.B1(out_sel[1]), 
	.B2(I1[5]), 
	.Z(O0[5])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_5 ( 
	.A1(out_sel[2]), 
	.A2(I2[5]), 
	.B1(out_sel[3]), 
	.B2(I3[5]), 
	.Z(O1[5])); 
	SC7P5T_AO22X0P5_SSC14R inst_2_5 ( 
	.A1(out_sel[4]), 
	.A2(I4[5]), 
	.B1(out_sel[5]), 
	.B2(I5[5]), 
	.Z(O2[5])); 
	SC7P5T_AO22X0P5_SSC14R inst_3_5 ( 
	.A1(out_sel[6]), 
	.A2(I6[5]), 
	.B1(out_sel[7]), 
	.B2(I7[5]), 
	.Z(O3[5])); 
	SC7P5T_AO22X0P5_SSC14R inst_4_5 ( 
	.A1(out_sel[8]), 
	.A2(I8[5]), 
	.B1(out_sel[9]), 
	.B2(I9[5]), 
	.Z(O4[5])); 
	SC7P5T_AO22X0P5_SSC14R inst_5_5 ( 
	.A1(out_sel[10]), 
	.A2(I10[5]), 
	.B1(out_sel[11]), 
	.B2(I11[5]), 
	.Z(O5[5])); 
	SC7P5T_AO22X0P5_SSC14R inst_6_5 ( 
	.A1(out_sel[12]), 
	.A2(I12[5]), 
	.B1(out_sel[13]), 
	.B2(I13[5]), 
	.Z(O6[5])); 
	SC7P5T_AO22X0P5_SSC14R inst_7_5 ( 
	.A1(out_sel[14]), 
	.A2(I14[5]), 
	.B1(out_sel[15]), 
	.B2(I15[5]), 
	.Z(O7[5])); 
	SC7P5T_AO22X0P5_SSC14R inst_8_5 ( 
	.A1(out_sel[16]), 
	.A2(I16[5]), 
	.B1(out_sel[17]), 
	.B2(I17[5]), 
	.Z(O8[5])); 
	SC7P5T_AO22X0P5_SSC14R inst_9_5 ( 
	.A1(out_sel[18]), 
	.A2(I18[5]), 
	.B1(out_sel[19]), 
	.B2(I19[5]), 
	.Z(O9[5])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_5 ( 
	.A(out_sel[20]), 
	.B(1'b0), 
	.Z(O10[5])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_6 ( 
	.A1(out_sel[0]), 
	.A2(I0[6]), 
	.B1(out_sel[1]), 
	.B2(I1[6]), 
	.Z(O0[6])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_6 ( 
	.A1(out_sel[2]), 
	.A2(I2[6]), 
	.B1(out_sel[3]), 
	.B2(I3[6]), 
	.Z(O1[6])); 
	SC7P5T_AO22X0P5_SSC14R inst_2_6 ( 
	.A1(out_sel[4]), 
	.A2(I4[6]), 
	.B1(out_sel[5]), 
	.B2(I5[6]), 
	.Z(O2[6])); 
	SC7P5T_AO22X0P5_SSC14R inst_3_6 ( 
	.A1(out_sel[6]), 
	.A2(I6[6]), 
	.B1(out_sel[7]), 
	.B2(I7[6]), 
	.Z(O3[6])); 
	SC7P5T_AO22X0P5_SSC14R inst_4_6 ( 
	.A1(out_sel[8]), 
	.A2(I8[6]), 
	.B1(out_sel[9]), 
	.B2(I9[6]), 
	.Z(O4[6])); 
	SC7P5T_AO22X0P5_SSC14R inst_5_6 ( 
	.A1(out_sel[10]), 
	.A2(I10[6]), 
	.B1(out_sel[11]), 
	.B2(I11[6]), 
	.Z(O5[6])); 
	SC7P5T_AO22X0P5_SSC14R inst_6_6 ( 
	.A1(out_sel[12]), 
	.A2(I12[6]), 
	.B1(out_sel[13]), 
	.B2(I13[6]), 
	.Z(O6[6])); 
	SC7P5T_AO22X0P5_SSC14R inst_7_6 ( 
	.A1(out_sel[14]), 
	.A2(I14[6]), 
	.B1(out_sel[15]), 
	.B2(I15[6]), 
	.Z(O7[6])); 
	SC7P5T_AO22X0P5_SSC14R inst_8_6 ( 
	.A1(out_sel[16]), 
	.A2(I16[6]), 
	.B1(out_sel[17]), 
	.B2(I17[6]), 
	.Z(O8[6])); 
	SC7P5T_AO22X0P5_SSC14R inst_9_6 ( 
	.A1(out_sel[18]), 
	.A2(I18[6]), 
	.B1(out_sel[19]), 
	.B2(I19[6]), 
	.Z(O9[6])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_6 ( 
	.A(out_sel[20]), 
	.B(1'b0), 
	.Z(O10[6])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_7 ( 
	.A1(out_sel[0]), 
	.A2(I0[7]), 
	.B1(out_sel[1]), 
	.B2(I1[7]), 
	.Z(O0[7])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_7 ( 
	.A1(out_sel[2]), 
	.A2(I2[7]), 
	.B1(out_sel[3]), 
	.B2(I3[7]), 
	.Z(O1[7])); 
	SC7P5T_AO22X0P5_SSC14R inst_2_7 ( 
	.A1(out_sel[4]), 
	.A2(I4[7]), 
	.B1(out_sel[5]), 
	.B2(I5[7]), 
	.Z(O2[7])); 
	SC7P5T_AO22X0P5_SSC14R inst_3_7 ( 
	.A1(out_sel[6]), 
	.A2(I6[7]), 
	.B1(out_sel[7]), 
	.B2(I7[7]), 
	.Z(O3[7])); 
	SC7P5T_AO22X0P5_SSC14R inst_4_7 ( 
	.A1(out_sel[8]), 
	.A2(I8[7]), 
	.B1(out_sel[9]), 
	.B2(I9[7]), 
	.Z(O4[7])); 
	SC7P5T_AO22X0P5_SSC14R inst_5_7 ( 
	.A1(out_sel[10]), 
	.A2(I10[7]), 
	.B1(out_sel[11]), 
	.B2(I11[7]), 
	.Z(O5[7])); 
	SC7P5T_AO22X0P5_SSC14R inst_6_7 ( 
	.A1(out_sel[12]), 
	.A2(I12[7]), 
	.B1(out_sel[13]), 
	.B2(I13[7]), 
	.Z(O6[7])); 
	SC7P5T_AO22X0P5_SSC14R inst_7_7 ( 
	.A1(out_sel[14]), 
	.A2(I14[7]), 
	.B1(out_sel[15]), 
	.B2(I15[7]), 
	.Z(O7[7])); 
	SC7P5T_AO22X0P5_SSC14R inst_8_7 ( 
	.A1(out_sel[16]), 
	.A2(I16[7]), 
	.B1(out_sel[17]), 
	.B2(I17[7]), 
	.Z(O8[7])); 
	SC7P5T_AO22X0P5_SSC14R inst_9_7 ( 
	.A1(out_sel[18]), 
	.A2(I18[7]), 
	.B1(out_sel[19]), 
	.B2(I19[7]), 
	.Z(O9[7])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_7 ( 
	.A(out_sel[20]), 
	.B(1'b0), 
	.Z(O10[7])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_8 ( 
	.A1(out_sel[0]), 
	.A2(I0[8]), 
	.B1(out_sel[1]), 
	.B2(I1[8]), 
	.Z(O0[8])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_8 ( 
	.A1(out_sel[2]), 
	.A2(I2[8]), 
	.B1(out_sel[3]), 
	.B2(I3[8]), 
	.Z(O1[8])); 
	SC7P5T_AO22X0P5_SSC14R inst_2_8 ( 
	.A1(out_sel[4]), 
	.A2(I4[8]), 
	.B1(out_sel[5]), 
	.B2(I5[8]), 
	.Z(O2[8])); 
	SC7P5T_AO22X0P5_SSC14R inst_3_8 ( 
	.A1(out_sel[6]), 
	.A2(I6[8]), 
	.B1(out_sel[7]), 
	.B2(I7[8]), 
	.Z(O3[8])); 
	SC7P5T_AO22X0P5_SSC14R inst_4_8 ( 
	.A1(out_sel[8]), 
	.A2(I8[8]), 
	.B1(out_sel[9]), 
	.B2(I9[8]), 
	.Z(O4[8])); 
	SC7P5T_AO22X0P5_SSC14R inst_5_8 ( 
	.A1(out_sel[10]), 
	.A2(I10[8]), 
	.B1(out_sel[11]), 
	.B2(I11[8]), 
	.Z(O5[8])); 
	SC7P5T_AO22X0P5_SSC14R inst_6_8 ( 
	.A1(out_sel[12]), 
	.A2(I12[8]), 
	.B1(out_sel[13]), 
	.B2(I13[8]), 
	.Z(O6[8])); 
	SC7P5T_AO22X0P5_SSC14R inst_7_8 ( 
	.A1(out_sel[14]), 
	.A2(I14[8]), 
	.B1(out_sel[15]), 
	.B2(I15[8]), 
	.Z(O7[8])); 
	SC7P5T_AO22X0P5_SSC14R inst_8_8 ( 
	.A1(out_sel[16]), 
	.A2(I16[8]), 
	.B1(out_sel[17]), 
	.B2(I17[8]), 
	.Z(O8[8])); 
	SC7P5T_AO22X0P5_SSC14R inst_9_8 ( 
	.A1(out_sel[18]), 
	.A2(I18[8]), 
	.B1(out_sel[19]), 
	.B2(I19[8]), 
	.Z(O9[8])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_8 ( 
	.A(out_sel[20]), 
	.B(1'b0), 
	.Z(O10[8])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_9 ( 
	.A1(out_sel[0]), 
	.A2(I0[9]), 
	.B1(out_sel[1]), 
	.B2(I1[9]), 
	.Z(O0[9])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_9 ( 
	.A1(out_sel[2]), 
	.A2(I2[9]), 
	.B1(out_sel[3]), 
	.B2(I3[9]), 
	.Z(O1[9])); 
	SC7P5T_AO22X0P5_SSC14R inst_2_9 ( 
	.A1(out_sel[4]), 
	.A2(I4[9]), 
	.B1(out_sel[5]), 
	.B2(I5[9]), 
	.Z(O2[9])); 
	SC7P5T_AO22X0P5_SSC14R inst_3_9 ( 
	.A1(out_sel[6]), 
	.A2(I6[9]), 
	.B1(out_sel[7]), 
	.B2(I7[9]), 
	.Z(O3[9])); 
	SC7P5T_AO22X0P5_SSC14R inst_4_9 ( 
	.A1(out_sel[8]), 
	.A2(I8[9]), 
	.B1(out_sel[9]), 
	.B2(I9[9]), 
	.Z(O4[9])); 
	SC7P5T_AO22X0P5_SSC14R inst_5_9 ( 
	.A1(out_sel[10]), 
	.A2(I10[9]), 
	.B1(out_sel[11]), 
	.B2(I11[9]), 
	.Z(O5[9])); 
	SC7P5T_AO22X0P5_SSC14R inst_6_9 ( 
	.A1(out_sel[12]), 
	.A2(I12[9]), 
	.B1(out_sel[13]), 
	.B2(I13[9]), 
	.Z(O6[9])); 
	SC7P5T_AO22X0P5_SSC14R inst_7_9 ( 
	.A1(out_sel[14]), 
	.A2(I14[9]), 
	.B1(out_sel[15]), 
	.B2(I15[9]), 
	.Z(O7[9])); 
	SC7P5T_AO22X0P5_SSC14R inst_8_9 ( 
	.A1(out_sel[16]), 
	.A2(I16[9]), 
	.B1(out_sel[17]), 
	.B2(I17[9]), 
	.Z(O8[9])); 
	SC7P5T_AO22X0P5_SSC14R inst_9_9 ( 
	.A1(out_sel[18]), 
	.A2(I18[9]), 
	.B1(out_sel[19]), 
	.B2(I19[9]), 
	.Z(O9[9])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_9 ( 
	.A(out_sel[20]), 
	.B(1'b0), 
	.Z(O10[9])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_10 ( 
	.A1(out_sel[0]), 
	.A2(I0[10]), 
	.B1(out_sel[1]), 
	.B2(I1[10]), 
	.Z(O0[10])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_10 ( 
	.A1(out_sel[2]), 
	.A2(I2[10]), 
	.B1(out_sel[3]), 
	.B2(I3[10]), 
	.Z(O1[10])); 
	SC7P5T_AO22X0P5_SSC14R inst_2_10 ( 
	.A1(out_sel[4]), 
	.A2(I4[10]), 
	.B1(out_sel[5]), 
	.B2(I5[10]), 
	.Z(O2[10])); 
	SC7P5T_AO22X0P5_SSC14R inst_3_10 ( 
	.A1(out_sel[6]), 
	.A2(I6[10]), 
	.B1(out_sel[7]), 
	.B2(I7[10]), 
	.Z(O3[10])); 
	SC7P5T_AO22X0P5_SSC14R inst_4_10 ( 
	.A1(out_sel[8]), 
	.A2(I8[10]), 
	.B1(out_sel[9]), 
	.B2(I9[10]), 
	.Z(O4[10])); 
	SC7P5T_AO22X0P5_SSC14R inst_5_10 ( 
	.A1(out_sel[10]), 
	.A2(I10[10]), 
	.B1(out_sel[11]), 
	.B2(I11[10]), 
	.Z(O5[10])); 
	SC7P5T_AO22X0P5_SSC14R inst_6_10 ( 
	.A1(out_sel[12]), 
	.A2(I12[10]), 
	.B1(out_sel[13]), 
	.B2(I13[10]), 
	.Z(O6[10])); 
	SC7P5T_AO22X0P5_SSC14R inst_7_10 ( 
	.A1(out_sel[14]), 
	.A2(I14[10]), 
	.B1(out_sel[15]), 
	.B2(I15[10]), 
	.Z(O7[10])); 
	SC7P5T_AO22X0P5_SSC14R inst_8_10 ( 
	.A1(out_sel[16]), 
	.A2(I16[10]), 
	.B1(out_sel[17]), 
	.B2(I17[10]), 
	.Z(O8[10])); 
	SC7P5T_AO22X0P5_SSC14R inst_9_10 ( 
	.A1(out_sel[18]), 
	.A2(I18[10]), 
	.B1(out_sel[19]), 
	.B2(I19[10]), 
	.Z(O9[10])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_10 ( 
	.A(out_sel[20]), 
	.B(1'b0), 
	.Z(O10[10])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_11 ( 
	.A1(out_sel[0]), 
	.A2(I0[11]), 
	.B1(out_sel[1]), 
	.B2(I1[11]), 
	.Z(O0[11])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_11 ( 
	.A1(out_sel[2]), 
	.A2(I2[11]), 
	.B1(out_sel[3]), 
	.B2(I3[11]), 
	.Z(O1[11])); 
	SC7P5T_AO22X0P5_SSC14R inst_2_11 ( 
	.A1(out_sel[4]), 
	.A2(I4[11]), 
	.B1(out_sel[5]), 
	.B2(I5[11]), 
	.Z(O2[11])); 
	SC7P5T_AO22X0P5_SSC14R inst_3_11 ( 
	.A1(out_sel[6]), 
	.A2(I6[11]), 
	.B1(out_sel[7]), 
	.B2(I7[11]), 
	.Z(O3[11])); 
	SC7P5T_AO22X0P5_SSC14R inst_4_11 ( 
	.A1(out_sel[8]), 
	.A2(I8[11]), 
	.B1(out_sel[9]), 
	.B2(I9[11]), 
	.Z(O4[11])); 
	SC7P5T_AO22X0P5_SSC14R inst_5_11 ( 
	.A1(out_sel[10]), 
	.A2(I10[11]), 
	.B1(out_sel[11]), 
	.B2(I11[11]), 
	.Z(O5[11])); 
	SC7P5T_AO22X0P5_SSC14R inst_6_11 ( 
	.A1(out_sel[12]), 
	.A2(I12[11]), 
	.B1(out_sel[13]), 
	.B2(I13[11]), 
	.Z(O6[11])); 
	SC7P5T_AO22X0P5_SSC14R inst_7_11 ( 
	.A1(out_sel[14]), 
	.A2(I14[11]), 
	.B1(out_sel[15]), 
	.B2(I15[11]), 
	.Z(O7[11])); 
	SC7P5T_AO22X0P5_SSC14R inst_8_11 ( 
	.A1(out_sel[16]), 
	.A2(I16[11]), 
	.B1(out_sel[17]), 
	.B2(I17[11]), 
	.Z(O8[11])); 
	SC7P5T_AO22X0P5_SSC14R inst_9_11 ( 
	.A1(out_sel[18]), 
	.A2(I18[11]), 
	.B1(out_sel[19]), 
	.B2(I19[11]), 
	.Z(O9[11])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_11 ( 
	.A(out_sel[20]), 
	.B(1'b0), 
	.Z(O10[11])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_12 ( 
	.A1(out_sel[0]), 
	.A2(I0[12]), 
	.B1(out_sel[1]), 
	.B2(I1[12]), 
	.Z(O0[12])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_12 ( 
	.A1(out_sel[2]), 
	.A2(I2[12]), 
	.B1(out_sel[3]), 
	.B2(I3[12]), 
	.Z(O1[12])); 
	SC7P5T_AO22X0P5_SSC14R inst_2_12 ( 
	.A1(out_sel[4]), 
	.A2(I4[12]), 
	.B1(out_sel[5]), 
	.B2(I5[12]), 
	.Z(O2[12])); 
	SC7P5T_AO22X0P5_SSC14R inst_3_12 ( 
	.A1(out_sel[6]), 
	.A2(I6[12]), 
	.B1(out_sel[7]), 
	.B2(I7[12]), 
	.Z(O3[12])); 
	SC7P5T_AO22X0P5_SSC14R inst_4_12 ( 
	.A1(out_sel[8]), 
	.A2(I8[12]), 
	.B1(out_sel[9]), 
	.B2(I9[12]), 
	.Z(O4[12])); 
	SC7P5T_AO22X0P5_SSC14R inst_5_12 ( 
	.A1(out_sel[10]), 
	.A2(I10[12]), 
	.B1(out_sel[11]), 
	.B2(I11[12]), 
	.Z(O5[12])); 
	SC7P5T_AO22X0P5_SSC14R inst_6_12 ( 
	.A1(out_sel[12]), 
	.A2(I12[12]), 
	.B1(out_sel[13]), 
	.B2(I13[12]), 
	.Z(O6[12])); 
	SC7P5T_AO22X0P5_SSC14R inst_7_12 ( 
	.A1(out_sel[14]), 
	.A2(I14[12]), 
	.B1(out_sel[15]), 
	.B2(I15[12]), 
	.Z(O7[12])); 
	SC7P5T_AO22X0P5_SSC14R inst_8_12 ( 
	.A1(out_sel[16]), 
	.A2(I16[12]), 
	.B1(out_sel[17]), 
	.B2(I17[12]), 
	.Z(O8[12])); 
	SC7P5T_AO22X0P5_SSC14R inst_9_12 ( 
	.A1(out_sel[18]), 
	.A2(I18[12]), 
	.B1(out_sel[19]), 
	.B2(I19[12]), 
	.Z(O9[12])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_12 ( 
	.A(out_sel[20]), 
	.B(1'b0), 
	.Z(O10[12])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_13 ( 
	.A1(out_sel[0]), 
	.A2(I0[13]), 
	.B1(out_sel[1]), 
	.B2(I1[13]), 
	.Z(O0[13])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_13 ( 
	.A1(out_sel[2]), 
	.A2(I2[13]), 
	.B1(out_sel[3]), 
	.B2(I3[13]), 
	.Z(O1[13])); 
	SC7P5T_AO22X0P5_SSC14R inst_2_13 ( 
	.A1(out_sel[4]), 
	.A2(I4[13]), 
	.B1(out_sel[5]), 
	.B2(I5[13]), 
	.Z(O2[13])); 
	SC7P5T_AO22X0P5_SSC14R inst_3_13 ( 
	.A1(out_sel[6]), 
	.A2(I6[13]), 
	.B1(out_sel[7]), 
	.B2(I7[13]), 
	.Z(O3[13])); 
	SC7P5T_AO22X0P5_SSC14R inst_4_13 ( 
	.A1(out_sel[8]), 
	.A2(I8[13]), 
	.B1(out_sel[9]), 
	.B2(I9[13]), 
	.Z(O4[13])); 
	SC7P5T_AO22X0P5_SSC14R inst_5_13 ( 
	.A1(out_sel[10]), 
	.A2(I10[13]), 
	.B1(out_sel[11]), 
	.B2(I11[13]), 
	.Z(O5[13])); 
	SC7P5T_AO22X0P5_SSC14R inst_6_13 ( 
	.A1(out_sel[12]), 
	.A2(I12[13]), 
	.B1(out_sel[13]), 
	.B2(I13[13]), 
	.Z(O6[13])); 
	SC7P5T_AO22X0P5_SSC14R inst_7_13 ( 
	.A1(out_sel[14]), 
	.A2(I14[13]), 
	.B1(out_sel[15]), 
	.B2(I15[13]), 
	.Z(O7[13])); 
	SC7P5T_AO22X0P5_SSC14R inst_8_13 ( 
	.A1(out_sel[16]), 
	.A2(I16[13]), 
	.B1(out_sel[17]), 
	.B2(I17[13]), 
	.Z(O8[13])); 
	SC7P5T_AO22X0P5_SSC14R inst_9_13 ( 
	.A1(out_sel[18]), 
	.A2(I18[13]), 
	.B1(out_sel[19]), 
	.B2(I19[13]), 
	.Z(O9[13])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_13 ( 
	.A(out_sel[20]), 
	.B(1'b0), 
	.Z(O10[13])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_14 ( 
	.A1(out_sel[0]), 
	.A2(I0[14]), 
	.B1(out_sel[1]), 
	.B2(I1[14]), 
	.Z(O0[14])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_14 ( 
	.A1(out_sel[2]), 
	.A2(I2[14]), 
	.B1(out_sel[3]), 
	.B2(I3[14]), 
	.Z(O1[14])); 
	SC7P5T_AO22X0P5_SSC14R inst_2_14 ( 
	.A1(out_sel[4]), 
	.A2(I4[14]), 
	.B1(out_sel[5]), 
	.B2(I5[14]), 
	.Z(O2[14])); 
	SC7P5T_AO22X0P5_SSC14R inst_3_14 ( 
	.A1(out_sel[6]), 
	.A2(I6[14]), 
	.B1(out_sel[7]), 
	.B2(I7[14]), 
	.Z(O3[14])); 
	SC7P5T_AO22X0P5_SSC14R inst_4_14 ( 
	.A1(out_sel[8]), 
	.A2(I8[14]), 
	.B1(out_sel[9]), 
	.B2(I9[14]), 
	.Z(O4[14])); 
	SC7P5T_AO22X0P5_SSC14R inst_5_14 ( 
	.A1(out_sel[10]), 
	.A2(I10[14]), 
	.B1(out_sel[11]), 
	.B2(I11[14]), 
	.Z(O5[14])); 
	SC7P5T_AO22X0P5_SSC14R inst_6_14 ( 
	.A1(out_sel[12]), 
	.A2(I12[14]), 
	.B1(out_sel[13]), 
	.B2(I13[14]), 
	.Z(O6[14])); 
	SC7P5T_AO22X0P5_SSC14R inst_7_14 ( 
	.A1(out_sel[14]), 
	.A2(I14[14]), 
	.B1(out_sel[15]), 
	.B2(I15[14]), 
	.Z(O7[14])); 
	SC7P5T_AO22X0P5_SSC14R inst_8_14 ( 
	.A1(out_sel[16]), 
	.A2(I16[14]), 
	.B1(out_sel[17]), 
	.B2(I17[14]), 
	.Z(O8[14])); 
	SC7P5T_AO22X0P5_SSC14R inst_9_14 ( 
	.A1(out_sel[18]), 
	.A2(I18[14]), 
	.B1(out_sel[19]), 
	.B2(I19[14]), 
	.Z(O9[14])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_14 ( 
	.A(out_sel[20]), 
	.B(1'b0), 
	.Z(O10[14])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_15 ( 
	.A1(out_sel[0]), 
	.A2(I0[15]), 
	.B1(out_sel[1]), 
	.B2(I1[15]), 
	.Z(O0[15])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_15 ( 
	.A1(out_sel[2]), 
	.A2(I2[15]), 
	.B1(out_sel[3]), 
	.B2(I3[15]), 
	.Z(O1[15])); 
	SC7P5T_AO22X0P5_SSC14R inst_2_15 ( 
	.A1(out_sel[4]), 
	.A2(I4[15]), 
	.B1(out_sel[5]), 
	.B2(I5[15]), 
	.Z(O2[15])); 
	SC7P5T_AO22X0P5_SSC14R inst_3_15 ( 
	.A1(out_sel[6]), 
	.A2(I6[15]), 
	.B1(out_sel[7]), 
	.B2(I7[15]), 
	.Z(O3[15])); 
	SC7P5T_AO22X0P5_SSC14R inst_4_15 ( 
	.A1(out_sel[8]), 
	.A2(I8[15]), 
	.B1(out_sel[9]), 
	.B2(I9[15]), 
	.Z(O4[15])); 
	SC7P5T_AO22X0P5_SSC14R inst_5_15 ( 
	.A1(out_sel[10]), 
	.A2(I10[15]), 
	.B1(out_sel[11]), 
	.B2(I11[15]), 
	.Z(O5[15])); 
	SC7P5T_AO22X0P5_SSC14R inst_6_15 ( 
	.A1(out_sel[12]), 
	.A2(I12[15]), 
	.B1(out_sel[13]), 
	.B2(I13[15]), 
	.Z(O6[15])); 
	SC7P5T_AO22X0P5_SSC14R inst_7_15 ( 
	.A1(out_sel[14]), 
	.A2(I14[15]), 
	.B1(out_sel[15]), 
	.B2(I15[15]), 
	.Z(O7[15])); 
	SC7P5T_AO22X0P5_SSC14R inst_8_15 ( 
	.A1(out_sel[16]), 
	.A2(I16[15]), 
	.B1(out_sel[17]), 
	.B2(I17[15]), 
	.Z(O8[15])); 
	SC7P5T_AO22X0P5_SSC14R inst_9_15 ( 
	.A1(out_sel[18]), 
	.A2(I18[15]), 
	.B1(out_sel[19]), 
	.B2(I19[15]), 
	.Z(O9[15])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_15 ( 
	.A(out_sel[20]), 
	.B(1'b0), 
	.Z(O10[15])); 
endmodule 

module mux_aoi_const_20_1 ( 
	input logic  [0 : 0] I0, 
	input logic  [0 : 0] I1, 
	input logic  [0 : 0] I2, 
	input logic  [0 : 0] I3, 
	input logic  [0 : 0] I4, 
	input logic  [0 : 0] I5, 
	input logic  [0 : 0] I6, 
	input logic  [0 : 0] I7, 
	input logic  [0 : 0] I8, 
	input logic  [0 : 0] I9, 
	input logic  [0 : 0] I10, 
	input logic  [0 : 0] I11, 
	input logic  [0 : 0] I12, 
	input logic  [0 : 0] I13, 
	input logic  [0 : 0] I14, 
	input logic  [0 : 0] I15, 
	input logic  [0 : 0] I16, 
	input logic  [0 : 0] I17, 
	input logic  [0 : 0] I18, 
	input logic  [0 : 0] I19, 
	input logic  [4 : 0] S ,
	output logic [0 : 0] O); 

	logic  [31 : 0] out_sel;
	logic  [0 : 0] O_int0;
	logic  [0 : 0] O_int1;
	logic  [0 : 0] O_int2;
	logic  [0 : 0] O_int3;
	logic  [0 : 0] O_int4;
	logic  [0 : 0] O_int5;
	logic  [0 : 0] O_int6;
	logic  [0 : 0] O_int7;
	logic  [0 : 0] O_int8;
	logic  [0 : 0] O_int9;
	logic  [0 : 0] O_int10;

precoder_1_20 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_1_20 u_mux_logic ( 
	.I0 (I0),
	.I1 (I1),
	.I2 (I2),
	.I3 (I3),
	.I4 (I4),
	.I5 (I5),
	.I6 (I6),
	.I7 (I7),
	.I8 (I8),
	.I9 (I9),
	.I10 (I10),
	.I11 (I11),
	.I12 (I12),
	.I13 (I13),
	.I14 (I14),
	.I15 (I15),
	.I16 (I16),
	.I17 (I17),
	.I18 (I18),
	.I19 (I19),
	.out_sel(out_sel), 
	.O0(O_int0), 
	.O1(O_int1), 
	.O2(O_int2), 
	.O3(O_int3), 
	.O4(O_int4), 
	.O5(O_int5), 
	.O6(O_int6), 
	.O7(O_int7), 
	.O8(O_int8), 
	.O9(O_int9), 
	.O10(O_int10)); 
	assign O = (  	O_int0 | 	O_int1 | 	O_int2 | 	O_int3 | 	O_int4 | 	O_int5 | 	O_int6 | 	O_int7 | 	O_int8 | 	O_int9 | 	O_int10 	); 

endmodule 

module precoder_1_20 (
	input logic  [4 : 0] S ,
	output logic  [31 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		5'd0    :   out_sel = 32'b00000000000000000000000000000001;
		5'd1    :   out_sel = 32'b00000000000000000000000000000010;
		5'd2    :   out_sel = 32'b00000000000000000000000000000100;
		5'd3    :   out_sel = 32'b00000000000000000000000000001000;
		5'd4    :   out_sel = 32'b00000000000000000000000000010000;
		5'd5    :   out_sel = 32'b00000000000000000000000000100000;
		5'd6    :   out_sel = 32'b00000000000000000000000001000000;
		5'd7    :   out_sel = 32'b00000000000000000000000010000000;
		5'd8    :   out_sel = 32'b00000000000000000000000100000000;
		5'd9    :   out_sel = 32'b00000000000000000000001000000000;
		5'd10    :   out_sel = 32'b00000000000000000000010000000000;
		5'd11    :   out_sel = 32'b00000000000000000000100000000000;
		5'd12    :   out_sel = 32'b00000000000000000001000000000000;
		5'd13    :   out_sel = 32'b00000000000000000010000000000000;
		5'd14    :   out_sel = 32'b00000000000000000100000000000000;
		5'd15    :   out_sel = 32'b00000000000000001000000000000000;
		5'd16    :   out_sel = 32'b00000000000000010000000000000000;
		5'd17    :   out_sel = 32'b00000000000000100000000000000000;
		5'd18    :   out_sel = 32'b00000000000001000000000000000000;
		5'd19    :   out_sel = 32'b00000000000010000000000000000000;
		5'd20    :   out_sel = 32'b00000000000100000000000000000000;
		default :   out_sel = 32'b0;
	endcase 
end 

endmodule 

module mux_logic_1_20 ( 
	input logic  [31 : 0] out_sel,
	input logic  [0 : 0] I0, 
	input logic  [0 : 0] I1, 
	input logic  [0 : 0] I2, 
	input logic  [0 : 0] I3, 
	input logic  [0 : 0] I4, 
	input logic  [0 : 0] I5, 
	input logic  [0 : 0] I6, 
	input logic  [0 : 0] I7, 
	input logic  [0 : 0] I8, 
	input logic  [0 : 0] I9, 
	input logic  [0 : 0] I10, 
	input logic  [0 : 0] I11, 
	input logic  [0 : 0] I12, 
	input logic  [0 : 0] I13, 
	input logic  [0 : 0] I14, 
	input logic  [0 : 0] I15, 
	input logic  [0 : 0] I16, 
	input logic  [0 : 0] I17, 
	input logic  [0 : 0] I18, 
	input logic  [0 : 0] I19, 
	output logic  [0 : 0] O0, 
	output logic  [0 : 0] O1, 
	output logic  [0 : 0] O2, 
	output logic  [0 : 0] O3, 
	output logic  [0 : 0] O4, 
	output logic  [0 : 0] O5, 
	output logic  [0 : 0] O6, 
	output logic  [0 : 0] O7, 
	output logic  [0 : 0] O8, 
	output logic  [0 : 0] O9, 
	output logic  [0 : 0] O10); 
	SC7P5T_AO22X0P5_SSC14R inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_0 ( 
	.A1(out_sel[2]), 
	.A2(I2[0]), 
	.B1(out_sel[3]), 
	.B2(I3[0]), 
	.Z(O1[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_2_0 ( 
	.A1(out_sel[4]), 
	.A2(I4[0]), 
	.B1(out_sel[5]), 
	.B2(I5[0]), 
	.Z(O2[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_3_0 ( 
	.A1(out_sel[6]), 
	.A2(I6[0]), 
	.B1(out_sel[7]), 
	.B2(I7[0]), 
	.Z(O3[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_4_0 ( 
	.A1(out_sel[8]), 
	.A2(I8[0]), 
	.B1(out_sel[9]), 
	.B2(I9[0]), 
	.Z(O4[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_5_0 ( 
	.A1(out_sel[10]), 
	.A2(I10[0]), 
	.B1(out_sel[11]), 
	.B2(I11[0]), 
	.Z(O5[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_6_0 ( 
	.A1(out_sel[12]), 
	.A2(I12[0]), 
	.B1(out_sel[13]), 
	.B2(I13[0]), 
	.Z(O6[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_7_0 ( 
	.A1(out_sel[14]), 
	.A2(I14[0]), 
	.B1(out_sel[15]), 
	.B2(I15[0]), 
	.Z(O7[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_8_0 ( 
	.A1(out_sel[16]), 
	.A2(I16[0]), 
	.B1(out_sel[17]), 
	.B2(I17[0]), 
	.Z(O8[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_9_0 ( 
	.A1(out_sel[18]), 
	.A2(I18[0]), 
	.B1(out_sel[19]), 
	.B2(I19[0]), 
	.Z(O9[0])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_0 ( 
	.A(out_sel[20]), 
	.B(1'b0), 
	.Z(O10[0])); 
endmodule 

module mux_aoi_7_1 ( 
	input logic  [0 : 0] I0, 
	input logic  [0 : 0] I1, 
	input logic  [0 : 0] I2, 
	input logic  [0 : 0] I3, 
	input logic  [0 : 0] I4, 
	input logic  [0 : 0] I5, 
	input logic  [0 : 0] I6, 
	input logic  [2 : 0] S ,
	output logic [0 : 0] O); 

	logic  [7 : 0] out_sel;
	logic  [0 : 0] O_int0;
	logic  [0 : 0] O_int1;
	logic  [0 : 0] O_int2;
	logic  [0 : 0] O_int3;

precoder_1_7 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_1_7 u_mux_logic ( 
	.I0 (I0),
	.I1 (I1),
	.I2 (I2),
	.I3 (I3),
	.I4 (I4),
	.I5 (I5),
	.I6 (I6),
	.out_sel(out_sel), 
	.O0(O_int0), 
	.O1(O_int1), 
	.O2(O_int2), 
	.O3(O_int3)); 
	assign O = (  	O_int0 | 	O_int1 | 	O_int2 | 	O_int3 	); 

endmodule 

module precoder_1_7 (
	input logic  [2 : 0] S ,
	output logic  [7 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		3'd0    :   out_sel = 8'b00000001;
		3'd1    :   out_sel = 8'b00000010;
		3'd2    :   out_sel = 8'b00000100;
		3'd3    :   out_sel = 8'b00001000;
		3'd4    :   out_sel = 8'b00010000;
		3'd5    :   out_sel = 8'b00100000;
		3'd6    :   out_sel = 8'b01000000;
		default :   out_sel = 8'b0;
	endcase 
end 

endmodule 

module mux_logic_1_7 ( 
	input logic  [7 : 0] out_sel,
	input logic  [0 : 0] I0, 
	input logic  [0 : 0] I1, 
	input logic  [0 : 0] I2, 
	input logic  [0 : 0] I3, 
	input logic  [0 : 0] I4, 
	input logic  [0 : 0] I5, 
	input logic  [0 : 0] I6, 
	output logic  [0 : 0] O0, 
	output logic  [0 : 0] O1, 
	output logic  [0 : 0] O2, 
	output logic  [0 : 0] O3); 
	SC7P5T_AO22X0P5_SSC14R inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_0 ( 
	.A1(out_sel[2]), 
	.A2(I2[0]), 
	.B1(out_sel[3]), 
	.B2(I3[0]), 
	.Z(O1[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_2_0 ( 
	.A1(out_sel[4]), 
	.A2(I4[0]), 
	.B1(out_sel[5]), 
	.B2(I5[0]), 
	.Z(O2[0])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_0 ( 
	.A(out_sel[6]), 
	.B(I6[0]), 
	.Z(O3[0])); 
endmodule 

module mux_aoi_5_16 ( 
	input logic  [15 : 0] I0, 
	input logic  [15 : 0] I1, 
	input logic  [15 : 0] I2, 
	input logic  [15 : 0] I3, 
	input logic  [15 : 0] I4, 
	input logic  [2 : 0] S ,
	output logic [15 : 0] O); 

	logic  [7 : 0] out_sel;
	logic  [15 : 0] O_int0;
	logic  [15 : 0] O_int1;
	logic  [15 : 0] O_int2;

precoder_16_5 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_16_5 u_mux_logic ( 
	.I0 (I0),
	.I1 (I1),
	.I2 (I2),
	.I3 (I3),
	.I4 (I4),
	.out_sel(out_sel), 
	.O0(O_int0), 
	.O1(O_int1), 
	.O2(O_int2)); 
	assign O = (  	O_int0 | 	O_int1 | 	O_int2 	); 

endmodule 

module precoder_16_5 (
	input logic  [2 : 0] S ,
	output logic  [7 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		3'd0    :   out_sel = 8'b00000001;
		3'd1    :   out_sel = 8'b00000010;
		3'd2    :   out_sel = 8'b00000100;
		3'd3    :   out_sel = 8'b00001000;
		3'd4    :   out_sel = 8'b00010000;
		default :   out_sel = 8'b0;
	endcase 
end 

endmodule 

module mux_logic_16_5 ( 
	input logic  [7 : 0] out_sel,
	input logic  [15 : 0] I0, 
	input logic  [15 : 0] I1, 
	input logic  [15 : 0] I2, 
	input logic  [15 : 0] I3, 
	input logic  [15 : 0] I4, 
	output logic  [15 : 0] O0, 
	output logic  [15 : 0] O1, 
	output logic  [15 : 0] O2); 
	SC7P5T_AO22X0P5_SSC14R inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_0 ( 
	.A1(out_sel[2]), 
	.A2(I2[0]), 
	.B1(out_sel[3]), 
	.B2(I3[0]), 
	.Z(O1[0])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_0 ( 
	.A(out_sel[4]), 
	.B(I4[0]), 
	.Z(O2[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_1 ( 
	.A1(out_sel[0]), 
	.A2(I0[1]), 
	.B1(out_sel[1]), 
	.B2(I1[1]), 
	.Z(O0[1])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_1 ( 
	.A1(out_sel[2]), 
	.A2(I2[1]), 
	.B1(out_sel[3]), 
	.B2(I3[1]), 
	.Z(O1[1])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_1 ( 
	.A(out_sel[4]), 
	.B(I4[1]), 
	.Z(O2[1])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_2 ( 
	.A1(out_sel[0]), 
	.A2(I0[2]), 
	.B1(out_sel[1]), 
	.B2(I1[2]), 
	.Z(O0[2])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_2 ( 
	.A1(out_sel[2]), 
	.A2(I2[2]), 
	.B1(out_sel[3]), 
	.B2(I3[2]), 
	.Z(O1[2])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_2 ( 
	.A(out_sel[4]), 
	.B(I4[2]), 
	.Z(O2[2])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_3 ( 
	.A1(out_sel[0]), 
	.A2(I0[3]), 
	.B1(out_sel[1]), 
	.B2(I1[3]), 
	.Z(O0[3])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_3 ( 
	.A1(out_sel[2]), 
	.A2(I2[3]), 
	.B1(out_sel[3]), 
	.B2(I3[3]), 
	.Z(O1[3])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_3 ( 
	.A(out_sel[4]), 
	.B(I4[3]), 
	.Z(O2[3])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_4 ( 
	.A1(out_sel[0]), 
	.A2(I0[4]), 
	.B1(out_sel[1]), 
	.B2(I1[4]), 
	.Z(O0[4])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_4 ( 
	.A1(out_sel[2]), 
	.A2(I2[4]), 
	.B1(out_sel[3]), 
	.B2(I3[4]), 
	.Z(O1[4])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_4 ( 
	.A(out_sel[4]), 
	.B(I4[4]), 
	.Z(O2[4])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_5 ( 
	.A1(out_sel[0]), 
	.A2(I0[5]), 
	.B1(out_sel[1]), 
	.B2(I1[5]), 
	.Z(O0[5])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_5 ( 
	.A1(out_sel[2]), 
	.A2(I2[5]), 
	.B1(out_sel[3]), 
	.B2(I3[5]), 
	.Z(O1[5])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_5 ( 
	.A(out_sel[4]), 
	.B(I4[5]), 
	.Z(O2[5])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_6 ( 
	.A1(out_sel[0]), 
	.A2(I0[6]), 
	.B1(out_sel[1]), 
	.B2(I1[6]), 
	.Z(O0[6])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_6 ( 
	.A1(out_sel[2]), 
	.A2(I2[6]), 
	.B1(out_sel[3]), 
	.B2(I3[6]), 
	.Z(O1[6])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_6 ( 
	.A(out_sel[4]), 
	.B(I4[6]), 
	.Z(O2[6])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_7 ( 
	.A1(out_sel[0]), 
	.A2(I0[7]), 
	.B1(out_sel[1]), 
	.B2(I1[7]), 
	.Z(O0[7])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_7 ( 
	.A1(out_sel[2]), 
	.A2(I2[7]), 
	.B1(out_sel[3]), 
	.B2(I3[7]), 
	.Z(O1[7])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_7 ( 
	.A(out_sel[4]), 
	.B(I4[7]), 
	.Z(O2[7])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_8 ( 
	.A1(out_sel[0]), 
	.A2(I0[8]), 
	.B1(out_sel[1]), 
	.B2(I1[8]), 
	.Z(O0[8])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_8 ( 
	.A1(out_sel[2]), 
	.A2(I2[8]), 
	.B1(out_sel[3]), 
	.B2(I3[8]), 
	.Z(O1[8])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_8 ( 
	.A(out_sel[4]), 
	.B(I4[8]), 
	.Z(O2[8])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_9 ( 
	.A1(out_sel[0]), 
	.A2(I0[9]), 
	.B1(out_sel[1]), 
	.B2(I1[9]), 
	.Z(O0[9])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_9 ( 
	.A1(out_sel[2]), 
	.A2(I2[9]), 
	.B1(out_sel[3]), 
	.B2(I3[9]), 
	.Z(O1[9])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_9 ( 
	.A(out_sel[4]), 
	.B(I4[9]), 
	.Z(O2[9])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_10 ( 
	.A1(out_sel[0]), 
	.A2(I0[10]), 
	.B1(out_sel[1]), 
	.B2(I1[10]), 
	.Z(O0[10])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_10 ( 
	.A1(out_sel[2]), 
	.A2(I2[10]), 
	.B1(out_sel[3]), 
	.B2(I3[10]), 
	.Z(O1[10])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_10 ( 
	.A(out_sel[4]), 
	.B(I4[10]), 
	.Z(O2[10])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_11 ( 
	.A1(out_sel[0]), 
	.A2(I0[11]), 
	.B1(out_sel[1]), 
	.B2(I1[11]), 
	.Z(O0[11])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_11 ( 
	.A1(out_sel[2]), 
	.A2(I2[11]), 
	.B1(out_sel[3]), 
	.B2(I3[11]), 
	.Z(O1[11])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_11 ( 
	.A(out_sel[4]), 
	.B(I4[11]), 
	.Z(O2[11])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_12 ( 
	.A1(out_sel[0]), 
	.A2(I0[12]), 
	.B1(out_sel[1]), 
	.B2(I1[12]), 
	.Z(O0[12])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_12 ( 
	.A1(out_sel[2]), 
	.A2(I2[12]), 
	.B1(out_sel[3]), 
	.B2(I3[12]), 
	.Z(O1[12])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_12 ( 
	.A(out_sel[4]), 
	.B(I4[12]), 
	.Z(O2[12])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_13 ( 
	.A1(out_sel[0]), 
	.A2(I0[13]), 
	.B1(out_sel[1]), 
	.B2(I1[13]), 
	.Z(O0[13])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_13 ( 
	.A1(out_sel[2]), 
	.A2(I2[13]), 
	.B1(out_sel[3]), 
	.B2(I3[13]), 
	.Z(O1[13])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_13 ( 
	.A(out_sel[4]), 
	.B(I4[13]), 
	.Z(O2[13])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_14 ( 
	.A1(out_sel[0]), 
	.A2(I0[14]), 
	.B1(out_sel[1]), 
	.B2(I1[14]), 
	.Z(O0[14])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_14 ( 
	.A1(out_sel[2]), 
	.A2(I2[14]), 
	.B1(out_sel[3]), 
	.B2(I3[14]), 
	.Z(O1[14])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_14 ( 
	.A(out_sel[4]), 
	.B(I4[14]), 
	.Z(O2[14])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_15 ( 
	.A1(out_sel[0]), 
	.A2(I0[15]), 
	.B1(out_sel[1]), 
	.B2(I1[15]), 
	.Z(O0[15])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_15 ( 
	.A1(out_sel[2]), 
	.A2(I2[15]), 
	.B1(out_sel[3]), 
	.B2(I3[15]), 
	.Z(O1[15])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_15 ( 
	.A(out_sel[4]), 
	.B(I4[15]), 
	.Z(O2[15])); 
endmodule 

module mux_aoi_5_1 ( 
	input logic  [0 : 0] I0, 
	input logic  [0 : 0] I1, 
	input logic  [0 : 0] I2, 
	input logic  [0 : 0] I3, 
	input logic  [0 : 0] I4, 
	input logic  [2 : 0] S ,
	output logic [0 : 0] O); 

	logic  [7 : 0] out_sel;
	logic  [0 : 0] O_int0;
	logic  [0 : 0] O_int1;
	logic  [0 : 0] O_int2;

precoder_1_5 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_1_5 u_mux_logic ( 
	.I0 (I0),
	.I1 (I1),
	.I2 (I2),
	.I3 (I3),
	.I4 (I4),
	.out_sel(out_sel), 
	.O0(O_int0), 
	.O1(O_int1), 
	.O2(O_int2)); 
	assign O = (  	O_int0 | 	O_int1 | 	O_int2 	); 

endmodule 

module precoder_1_5 (
	input logic  [2 : 0] S ,
	output logic  [7 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		3'd0    :   out_sel = 8'b00000001;
		3'd1    :   out_sel = 8'b00000010;
		3'd2    :   out_sel = 8'b00000100;
		3'd3    :   out_sel = 8'b00001000;
		3'd4    :   out_sel = 8'b00010000;
		default :   out_sel = 8'b0;
	endcase 
end 

endmodule 

module mux_logic_1_5 ( 
	input logic  [7 : 0] out_sel,
	input logic  [0 : 0] I0, 
	input logic  [0 : 0] I1, 
	input logic  [0 : 0] I2, 
	input logic  [0 : 0] I3, 
	input logic  [0 : 0] I4, 
	output logic  [0 : 0] O0, 
	output logic  [0 : 0] O1, 
	output logic  [0 : 0] O2); 
	SC7P5T_AO22X0P5_SSC14R inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_1_0 ( 
	.A1(out_sel[2]), 
	.A2(I2[0]), 
	.B1(out_sel[3]), 
	.B2(I3[0]), 
	.Z(O1[0])); 
	SC7P5T_AN2X0P5_SSC14R inst_and_0 ( 
	.A(out_sel[4]), 
	.B(I4[0]), 
	.Z(O2[0])); 
endmodule 

module mux_aoi_2_16 ( 
	input logic  [15 : 0] I0, 
	input logic  [15 : 0] I1, 
input logic S, 
	output logic [15 : 0] O); 

	logic  [1 : 0] out_sel;
	logic  [15 : 0] O_int0;

precoder_16_2 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_16_2 u_mux_logic ( 
	.I0 (I0),
	.I1 (I1),
	.out_sel(out_sel), 
	.O0(O_int0)); 
	assign O = (  	O_int0 	); 

endmodule 

module precoder_16_2 (
	input logic  [0 : 0] S ,
	output logic  [1 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		1'd0    :   out_sel = 2'b01;
		1'd1    :   out_sel = 2'b10;
		default :   out_sel = 2'b0;
	endcase 
end 

endmodule 

module mux_logic_16_2 ( 
	input logic  [1 : 0] out_sel,
	input logic  [15 : 0] I0, 
	input logic  [15 : 0] I1, 
	output logic  [15 : 0] O0); 
	SC7P5T_AO22X0P5_SSC14R inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_1 ( 
	.A1(out_sel[0]), 
	.A2(I0[1]), 
	.B1(out_sel[1]), 
	.B2(I1[1]), 
	.Z(O0[1])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_2 ( 
	.A1(out_sel[0]), 
	.A2(I0[2]), 
	.B1(out_sel[1]), 
	.B2(I1[2]), 
	.Z(O0[2])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_3 ( 
	.A1(out_sel[0]), 
	.A2(I0[3]), 
	.B1(out_sel[1]), 
	.B2(I1[3]), 
	.Z(O0[3])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_4 ( 
	.A1(out_sel[0]), 
	.A2(I0[4]), 
	.B1(out_sel[1]), 
	.B2(I1[4]), 
	.Z(O0[4])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_5 ( 
	.A1(out_sel[0]), 
	.A2(I0[5]), 
	.B1(out_sel[1]), 
	.B2(I1[5]), 
	.Z(O0[5])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_6 ( 
	.A1(out_sel[0]), 
	.A2(I0[6]), 
	.B1(out_sel[1]), 
	.B2(I1[6]), 
	.Z(O0[6])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_7 ( 
	.A1(out_sel[0]), 
	.A2(I0[7]), 
	.B1(out_sel[1]), 
	.B2(I1[7]), 
	.Z(O0[7])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_8 ( 
	.A1(out_sel[0]), 
	.A2(I0[8]), 
	.B1(out_sel[1]), 
	.B2(I1[8]), 
	.Z(O0[8])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_9 ( 
	.A1(out_sel[0]), 
	.A2(I0[9]), 
	.B1(out_sel[1]), 
	.B2(I1[9]), 
	.Z(O0[9])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_10 ( 
	.A1(out_sel[0]), 
	.A2(I0[10]), 
	.B1(out_sel[1]), 
	.B2(I1[10]), 
	.Z(O0[10])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_11 ( 
	.A1(out_sel[0]), 
	.A2(I0[11]), 
	.B1(out_sel[1]), 
	.B2(I1[11]), 
	.Z(O0[11])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_12 ( 
	.A1(out_sel[0]), 
	.A2(I0[12]), 
	.B1(out_sel[1]), 
	.B2(I1[12]), 
	.Z(O0[12])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_13 ( 
	.A1(out_sel[0]), 
	.A2(I0[13]), 
	.B1(out_sel[1]), 
	.B2(I1[13]), 
	.Z(O0[13])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_14 ( 
	.A1(out_sel[0]), 
	.A2(I0[14]), 
	.B1(out_sel[1]), 
	.B2(I1[14]), 
	.Z(O0[14])); 
	SC7P5T_AO22X0P5_SSC14R inst_0_15 ( 
	.A1(out_sel[0]), 
	.A2(I0[15]), 
	.B1(out_sel[1]), 
	.B2(I1[15]), 
	.Z(O0[15])); 
endmodule 

module mux_aoi_2_1 ( 
	input logic  [0 : 0] I0, 
	input logic  [0 : 0] I1, 
input logic S, 
	output logic [0 : 0] O); 

	logic  [1 : 0] out_sel;
	logic  [0 : 0] O_int0;

precoder_1_2 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_1_2 u_mux_logic ( 
	.I0 (I0),
	.I1 (I1),
	.out_sel(out_sel), 
	.O0(O_int0)); 
	assign O = (  	O_int0 	); 

endmodule 

module precoder_1_2 (
	input logic  [0 : 0] S ,
	output logic  [1 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		1'd0    :   out_sel = 2'b01;
		1'd1    :   out_sel = 2'b10;
		default :   out_sel = 2'b0;
	endcase 
end 

endmodule 

module mux_logic_1_2 ( 
	input logic  [1 : 0] out_sel,
	input logic  [0 : 0] I0, 
	input logic  [0 : 0] I1, 
	output logic  [0 : 0] O0); 
	SC7P5T_AO22X0P5_SSC14R inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
endmodule 

module mode (
    input [26:0] I,
    output [1:0] O
);
assign O = I[25:24];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5 (
    input [26:0] I,
    output [3:0] O
);
assign O = I[23:20];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4 (
    input [26:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3 (
    input [26:0] I,
    output [3:0] O
);
assign O = I[15:12];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2 (
    input [26:0] I,
    output [3:0] O
);
assign O = I[11:8];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1 (
    input [26:0] I,
    output [3:0] O
);
assign O = I[7:4];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0 (
    input [26:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr (
    input [31:0] I,
    output [3:0] O
);
assign O = I[31:28];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[27:24];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[23:20];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[15:12];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[11:8];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[7:4];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr (
    input [31:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr (
    input [16:0] I,
    output [15:0] O
);
assign O = I[16:1];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable (
    input [16:0] I,
    output [0:0] O
);
assign O = I[0:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr (
    input [24:0] I,
    output [15:0] O
);
assign O = I[24:9];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable (
    input [24:0] I,
    output [0:0] O
);
assign O = I[8:8];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5 (
    input [24:0] I,
    output [3:0] O
);
assign O = I[7:4];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4 (
    input [24:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[31:28];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[27:24];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[23:20];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr (
    input [31:0] I,
    output [3:0] O
);
assign O = I[15:12];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[11:8];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[7:4];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[31:28];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[27:24];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[23:20];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr (
    input [31:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0 (
    input [19:0] I,
    output [15:0] O
);
assign O = I[19:4];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality (
    input [19:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality (
    input [19:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5 (
    input [19:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable (
    input [16:0] I,
    output [0:0] O
);
assign O = I[16:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5 (
    input [16:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable (
    input [16:0] I,
    output [0:0] O
);
assign O = I[16:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5 (
    input [16:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0 (
    input [19:0] I,
    output [15:0] O
);
assign O = I[19:4];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality (
    input [19:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality (
    input [30:0] I,
    output [3:0] O
);
assign O = I[30:27];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5 (
    input [30:0] I,
    output [8:0] O
);
assign O = I[26:18];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4 (
    input [30:0] I,
    output [8:0] O
);
assign O = I[17:9];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3 (
    input [30:0] I,
    output [8:0] O
);
assign O = I[8:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[26:18];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[17:9];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[8:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr (
    input [26:0] I,
    output [8:0] O
);
assign O = I[26:18];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[17:9];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[8:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[26:18];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[17:9];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[8:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[26:18];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr (
    input [26:0] I,
    output [8:0] O
);
assign O = I[17:9];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[8:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[26:18];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[17:9];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[8:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[26:18];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[17:9];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr (
    input [26:0] I,
    output [8:0] O
);
assign O = I[8:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[26:18];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[17:9];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[8:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[26:18];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[17:9];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[8:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr (
    input [25:0] I,
    output [8:0] O
);
assign O = I[25:17];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en (
    input [25:0] I,
    output [0:0] O
);
assign O = I[16:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5 (
    input [25:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0 (
    input [19:0] I,
    output [15:0] O
);
assign O = I[19:4];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality (
    input [19:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality (
    input [19:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5 (
    input [19:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable (
    input [16:0] I,
    output [0:0] O
);
assign O = I[16:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5 (
    input [16:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable (
    input [16:0] I,
    output [0:0] O
);
assign O = I[16:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5 (
    input [16:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0 (
    input [19:0] I,
    output [15:0] O
);
assign O = I[19:4];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality (
    input [19:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality (
    input [19:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5 (
    input [19:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable (
    input [16:0] I,
    output [0:0] O
);
assign O = I[16:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5 (
    input [16:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable (
    input [16:0] I,
    output [0:0] O
);
assign O = I[16:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5 (
    input [16:0] I,
    output [3:0] O
);
assign O = I[15:12];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4 (
    input [16:0] I,
    output [3:0] O
);
assign O = I[11:8];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3 (
    input [16:0] I,
    output [3:0] O
);
assign O = I[7:4];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2 (
    input [16:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[31:28];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[27:24];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr (
    input [31:0] I,
    output [3:0] O
);
assign O = I[23:20];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[15:12];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[11:8];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[7:4];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[31:28];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr (
    input [31:0] I,
    output [3:0] O
);
assign O = I[27:24];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[23:20];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[15:12];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[11:8];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[7:4];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr (
    input [31:0] I,
    output [3:0] O
);
assign O = I[31:28];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[27:24];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[23:20];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[15:12];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[11:8];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[7:4];
endmodule

module mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr (
    input [31:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module mem_ctrl_strg_fifo_flat_strg_fifo_inst_fifo_depth (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable (
    input [16:0] I,
    output [0:0] O
);
assign O = I[16:16];
endmodule

module mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5 (
    input [16:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0 (
    input [24:0] I,
    output [15:0] O
);
assign O = I[24:9];
endmodule

module mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality (
    input [24:0] I,
    output [3:0] O
);
assign O = I[8:5];
endmodule

module mantle_wire__typeBitIn81 (
    output [80:0] in,
    input [80:0] out
);
assign in = out;
endmodule

module mantle_wire__typeBitIn32 (
    output [31:0] in,
    input [31:0] out
);
assign in = out;
endmodule

module mantle_wire__typeBit8 (
    input [7:0] in,
    output [7:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit4 (
    input [3:0] in,
    output [3:0] out
);
assign out = in;
endmodule

module regCE_arst #(
    parameter width = 1,
    parameter init = 1
) (
    input [width-1:0] in,
    input ce,
    output [width-1:0] out,
    input clk,
    input arst
);
  reg [width-1:0] value;
  always @(posedge clk, posedge arst) begin
    if (arst) begin
      value <= init;
    end
    else if (ce) begin
      value <= in;
    end
  end
  assign out = value;
endmodule

module regCE #(
    parameter width = 1
) (
    input [width-1:0] in,
    input ce,
    output [width-1:0] out,
    input clk
);
  reg [width-1:0] value;
  always @(posedge clk) begin
    if (ce) begin
      value <= in;
    end
  end
  assign out = value;
endmodule

module io_core (
    input [15:0] glb2io_16,
    input [0:0] glb2io_1,
    output [15:0] io2glb_16,
    output [0:0] io2glb_1,
    input [15:0] f2io_16,
    input [0:0] f2io_1,
    output [15:0] io2f_16,
    output [0:0] io2f_1
);
assign io2glb_16 = f2io_16;
assign io2glb_1 = f2io_1;
assign io2f_16 = glb2io_16;
assign io2f_1 = glb2io_1;
endmodule

module inst_2 (
    input [31:0] I,
    output [31:0] O
);
assign O = I;
endmodule

module inst_1 (
    input [31:0] I,
    output [31:0] O
);
assign O = I;
endmodule

module inst_0 (
    input [31:0] I,
    output [31:0] O
);
assign O = I;
endmodule

module input_width_1_num_1_reg_value (
    input [24:0] I,
    output [0:0] O
);
assign O = I[4:4];
endmodule

module input_width_1_num_1_reg_sel (
    input [24:0] I,
    output [0:0] O
);
assign O = I[3:3];
endmodule

module input_width_1_num_0_reg_value (
    input [24:0] I,
    output [0:0] O
);
assign O = I[2:2];
endmodule

module input_width_1_num_0_reg_sel (
    input [24:0] I,
    output [0:0] O
);
assign O = I[1:1];
endmodule

typedef struct packed {
    logic mode;
    logic [15:0] relocation_value;
    logic relocation_is_msb;
} pcfg_dma_ctrl_t;

typedef struct packed {
    logic wr_en;
    logic [7:0] wr_strb;
    logic [18:0] wr_addr;
    logic [63:0] wr_data;
} wr_packet_t;

typedef struct packed {
    logic [1:0] west;
    logic [1:0] east;
    logic [1:0] south;
} pcfg_broadcast_mux_t;

typedef struct packed {
    logic [63:0] rd_data;
    logic rd_data_valid;
} rdrs_packet_t;

typedef struct packed {
    logic rd_en;
    logic [18:0] rd_addr;
} rdrq_packet_t;

typedef struct packed {
rdrq_packet_t rdrq;
rdrs_packet_t rdrs;
} rd_packet_t;

typedef struct packed {
wr_packet_t wr;
rdrq_packet_t rdrq;
rdrs_packet_t rdrs;
} packet_t;

typedef struct packed {
    logic [18:0] start_addr;
    logic [15:0] cycle_start_addr;
    logic [3:0] dim;
    logic [31:0] range_0;
    logic [19:0] stride_0;
    logic [15:0] cycle_stride_0;
    logic [31:0] range_1;
    logic [19:0] stride_1;
    logic [15:0] cycle_stride_1;
    logic [31:0] range_2;
    logic [19:0] stride_2;
    logic [15:0] cycle_stride_2;
    logic [31:0] range_3;
    logic [19:0] stride_3;
    logic [15:0] cycle_stride_3;
    logic [31:0] range_4;
    logic [19:0] stride_4;
    logic [15:0] cycle_stride_4;
    logic [31:0] range_5;
    logic [19:0] stride_5;
    logic [15:0] cycle_stride_5;
    logic [31:0] range_6;
    logic [19:0] stride_6;
    logic [15:0] cycle_stride_6;
    logic [31:0] range_7;
    logic [19:0] stride_7;
    logic [15:0] cycle_stride_7;
} dma_header_t;

typedef struct packed {
    logic [1:0] mode;
    logic use_valid;
    logic use_flush;
    logic [1:0] data_mux;
    logic num_repeat;
} load_dma_ctrl_t;

typedef struct packed {
    logic rd_en;
    logic wr_en;
    logic [31:0] addr;
    logic [31:0] data;
} cgra_cfg_t;

typedef struct packed {
    logic [18:0] start_addr;
    logic [15:0] num_cfg;
} pcfg_dma_header_t;

typedef struct packed {
    logic tile_connected;
    logic [5:0] latency;
} cfg_pcfg_network_t;

typedef struct packed {
    logic tile_connected;
    logic [5:0] latency;
} cfg_data_network_t;

typedef struct packed {
    logic rd_en;
    logic [16:0] rd_addr;
} rdrq_bank_packet_t;

typedef struct packed {
    logic [1:0] mode;
    logic use_valid;
    logic [1:0] data_mux;
    logic num_repeat;
} store_dma_ctrl_t;

typedef struct packed {
    logic wr_en;
    logic [7:0] wr_strb;
    logic [16:0] wr_addr;
    logic [63:0] wr_data;
} wr_bank_packet_t;

interface glb_tile_ifc_A_12_D_32;
  logic [11:0] rd_addr;
  logic rd_clk_en;
  logic [31:0] rd_data;
  logic rd_data_valid;
  logic rd_en;
  logic [11:0] wr_addr;
  logic wr_clk_en;
  logic [31:0] wr_data;
  logic wr_en;
  modport master(input rd_data, input rd_data_valid, output rd_addr, output rd_clk_en, output rd_en, output wr_addr, output wr_clk_en, output wr_data, output wr_en);
  modport slave(input rd_addr, input rd_clk_en, input rd_en, input wr_addr, input wr_clk_en, input wr_data, input wr_en, output rd_data, output rd_data_valid);
endinterface

interface glb_tile_ifc_A_19_D_32;
  logic [18:0] rd_addr;
  logic rd_clk_en;
  logic [31:0] rd_data;
  logic rd_data_valid;
  logic rd_en;
  logic [18:0] wr_addr;
  logic wr_clk_en;
  logic [31:0] wr_data;
  logic wr_en;
  modport master(input rd_data, input rd_data_valid, output rd_addr, output rd_clk_en, output rd_en, output wr_addr, output wr_clk_en, output wr_data, output wr_en);
  modport slave(input rd_addr, input rd_clk_en, input rd_en, input wr_addr, input wr_clk_en, input wr_data, input wr_en, output rd_data, output rd_data_valid);
endinterface

interface glb_tile_ifc_A_19_D_64;
  logic [18:0] rd_addr;
  logic rd_clk_en;
  logic [63:0] rd_data;
  logic rd_data_valid;
  logic rd_en;
  logic [18:0] wr_addr;
  logic wr_clk_en;
  logic [63:0] wr_data;
  logic wr_en;
  logic [7:0] wr_strb;
  modport master(input rd_data, input rd_data_valid, output rd_addr, output rd_clk_en, output rd_en, output wr_addr, output wr_clk_en, output wr_data, output wr_en, output wr_strb);
  modport slave(input rd_addr, input rd_clk_en, input rd_en, input wr_addr, input wr_clk_en, input wr_data, input wr_en, input wr_strb, output rd_data, output rd_data_valid);
endinterface

module IN12LP_S1DB_W04096B064M08S2_HB (
  input logic [11:0] A,
  input logic [63:0] BW,
  input logic CEN,
  input logic CLK,
  input logic [63:0] D,
  input logic MA_SAWL0,
  input logic MA_SAWL1,
  input logic MA_STABAS0,
  input logic MA_STABAS1,
  input logic MA_VD0,
  input logic MA_VD1,
  input logic MA_WL0,
  input logic MA_WL1,
  input logic MA_WRAS0,
  input logic MA_WRAS1,
  input logic MA_WRT,
  input logic RDWEN,
  input logic T_LOGIC,
  input logic T_Q_RST,
  output logic [63:0] Q
);

logic [63:0] data_array [4095:0];

always_ff @(posedge CLK) begin
  if (CEN == 1'h0) begin
    Q <= data_array[A];
    if (RDWEN == 1'h0) begin
      for (int unsigned i = 0; i < 64; i += 1) begin
          if (BW[6'(i)]) begin
            data_array[A][6'(i)] <= D[6'(i)];
          end
        end
    end
  end
end
endmodule   // IN12LP_S1DB_W04096B064M08S2_HB

module SC7P5T_CKGPRELATNX1_SSC14R (
  input logic CLK,
  input logic E,
  input logic TE,
  output logic Z
);

logic enable_latch;
always_latch begin
  if (~CLK) begin
    enable_latch = E;
  end
end
assign Z = CLK & enable_latch;
endmodule   // SC7P5T_CKGPRELATNX1_SSC14R

module clk_gate (
  input logic clk,
  input logic enable,
  output logic gclk
);

SC7P5T_CKGPRELATNX1_SSC14R CG_CELL (
  .CLK(clk),
  .E(enable),
  .TE(1'h0),
  .Z(gclk)
);

endmodule   // clk_gate

module glb_addr_gen #(
  parameter addr_width = 32'h10
)
(
  input logic clk,
  input logic clk_en,
  input logic [2:0] mux_sel,
  input logic reset,
  input logic restart,
  input logic [addr_width-1:0] start_addr,
  input logic step,
  input logic [7:0] [addr_width-1:0] strides,
  output logic [addr_width-1:0] addr_out
);

logic [addr_width-1:0] current_addr;
assign addr_out = start_addr + current_addr;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    current_addr <= 16'h0;
  end
  else if (clk_en) begin
    if (restart) begin
      current_addr <= 16'h0;
    end
    else if (step) begin
      current_addr <= current_addr + strides[mux_sel];
    end
  end
end
endmodule   // glb_addr_gen

module glb_bank (
  input logic clk,
  input rdrq_bank_packet_t rdrq_packet,
  input logic reset,
  input wr_bank_packet_t wr_packet,
  output rdrs_packet_t rdrs_packet
);

logic [16:0] mem_addr;
logic [63:0] mem_data_in;
logic [63:0] mem_data_in_bit_sel;
logic [63:0] mem_data_out;
logic mem_rd_en;
logic mem_wr_en;
logic [63:0] packet_rd_data_r;
logic packet_rd_en_d;
logic [63:0] wr_data_bit_sel;
assign wr_data_bit_sel[0] = wr_packet.wr_strb[0];
assign wr_data_bit_sel[1] = wr_packet.wr_strb[0];
assign wr_data_bit_sel[2] = wr_packet.wr_strb[0];
assign wr_data_bit_sel[3] = wr_packet.wr_strb[0];
assign wr_data_bit_sel[4] = wr_packet.wr_strb[0];
assign wr_data_bit_sel[5] = wr_packet.wr_strb[0];
assign wr_data_bit_sel[6] = wr_packet.wr_strb[0];
assign wr_data_bit_sel[7] = wr_packet.wr_strb[0];
assign wr_data_bit_sel[8] = wr_packet.wr_strb[1];
assign wr_data_bit_sel[9] = wr_packet.wr_strb[1];
assign wr_data_bit_sel[10] = wr_packet.wr_strb[1];
assign wr_data_bit_sel[11] = wr_packet.wr_strb[1];
assign wr_data_bit_sel[12] = wr_packet.wr_strb[1];
assign wr_data_bit_sel[13] = wr_packet.wr_strb[1];
assign wr_data_bit_sel[14] = wr_packet.wr_strb[1];
assign wr_data_bit_sel[15] = wr_packet.wr_strb[1];
assign wr_data_bit_sel[16] = wr_packet.wr_strb[2];
assign wr_data_bit_sel[17] = wr_packet.wr_strb[2];
assign wr_data_bit_sel[18] = wr_packet.wr_strb[2];
assign wr_data_bit_sel[19] = wr_packet.wr_strb[2];
assign wr_data_bit_sel[20] = wr_packet.wr_strb[2];
assign wr_data_bit_sel[21] = wr_packet.wr_strb[2];
assign wr_data_bit_sel[22] = wr_packet.wr_strb[2];
assign wr_data_bit_sel[23] = wr_packet.wr_strb[2];
assign wr_data_bit_sel[24] = wr_packet.wr_strb[3];
assign wr_data_bit_sel[25] = wr_packet.wr_strb[3];
assign wr_data_bit_sel[26] = wr_packet.wr_strb[3];
assign wr_data_bit_sel[27] = wr_packet.wr_strb[3];
assign wr_data_bit_sel[28] = wr_packet.wr_strb[3];
assign wr_data_bit_sel[29] = wr_packet.wr_strb[3];
assign wr_data_bit_sel[30] = wr_packet.wr_strb[3];
assign wr_data_bit_sel[31] = wr_packet.wr_strb[3];
assign wr_data_bit_sel[32] = wr_packet.wr_strb[4];
assign wr_data_bit_sel[33] = wr_packet.wr_strb[4];
assign wr_data_bit_sel[34] = wr_packet.wr_strb[4];
assign wr_data_bit_sel[35] = wr_packet.wr_strb[4];
assign wr_data_bit_sel[36] = wr_packet.wr_strb[4];
assign wr_data_bit_sel[37] = wr_packet.wr_strb[4];
assign wr_data_bit_sel[38] = wr_packet.wr_strb[4];
assign wr_data_bit_sel[39] = wr_packet.wr_strb[4];
assign wr_data_bit_sel[40] = wr_packet.wr_strb[5];
assign wr_data_bit_sel[41] = wr_packet.wr_strb[5];
assign wr_data_bit_sel[42] = wr_packet.wr_strb[5];
assign wr_data_bit_sel[43] = wr_packet.wr_strb[5];
assign wr_data_bit_sel[44] = wr_packet.wr_strb[5];
assign wr_data_bit_sel[45] = wr_packet.wr_strb[5];
assign wr_data_bit_sel[46] = wr_packet.wr_strb[5];
assign wr_data_bit_sel[47] = wr_packet.wr_strb[5];
assign wr_data_bit_sel[48] = wr_packet.wr_strb[6];
assign wr_data_bit_sel[49] = wr_packet.wr_strb[6];
assign wr_data_bit_sel[50] = wr_packet.wr_strb[6];
assign wr_data_bit_sel[51] = wr_packet.wr_strb[6];
assign wr_data_bit_sel[52] = wr_packet.wr_strb[6];
assign wr_data_bit_sel[53] = wr_packet.wr_strb[6];
assign wr_data_bit_sel[54] = wr_packet.wr_strb[6];
assign wr_data_bit_sel[55] = wr_packet.wr_strb[6];
assign wr_data_bit_sel[56] = wr_packet.wr_strb[7];
assign wr_data_bit_sel[57] = wr_packet.wr_strb[7];
assign wr_data_bit_sel[58] = wr_packet.wr_strb[7];
assign wr_data_bit_sel[59] = wr_packet.wr_strb[7];
assign wr_data_bit_sel[60] = wr_packet.wr_strb[7];
assign wr_data_bit_sel[61] = wr_packet.wr_strb[7];
assign wr_data_bit_sel[62] = wr_packet.wr_strb[7];
assign wr_data_bit_sel[63] = wr_packet.wr_strb[7];
always_comb begin
  if (wr_packet.wr_en) begin
    mem_wr_en = 1'h1;
    mem_rd_en = 1'h0;
    mem_addr = wr_packet.wr_addr;
    mem_data_in = wr_packet.wr_data;
    mem_data_in_bit_sel = wr_data_bit_sel;
  end
  else if (rdrq_packet.rd_en) begin
    mem_wr_en = 1'h0;
    mem_rd_en = 1'h1;
    mem_addr = rdrq_packet.rd_addr;
    mem_data_in = 64'h0;
    mem_data_in_bit_sel = 64'h0;
  end
  else begin
    mem_wr_en = 1'h0;
    mem_rd_en = 1'h0;
    mem_addr = 17'h0;
    mem_data_in = 64'h0;
    mem_data_in_bit_sel = 64'h0;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    packet_rd_data_r <= 64'h0;
  end
  else packet_rd_data_r <= rdrs_packet.rd_data;
end
always_comb begin
  if (packet_rd_en_d) begin
    rdrs_packet.rd_data = mem_data_out;
  end
  else rdrs_packet.rd_data = packet_rd_data_r;
  rdrs_packet.rd_data_valid = packet_rd_en_d;
end
glb_bank_memory glb_bank_memory (
  .addr(mem_addr),
  .clk(clk),
  .data_in(mem_data_in),
  .data_in_bit_sel(mem_data_in_bit_sel),
  .ren(mem_rd_en),
  .reset(reset),
  .wen(mem_wr_en),
  .data_out(mem_data_out)
);

pipeline_w_1_d_1 packet_rdrq_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(rdrq_packet.rd_en),
  .reset(reset),
  .out_(packet_rd_en_d)
);

endmodule   // glb_bank

module glb_bank_memory (
  input logic [16:0] addr,
  input logic clk,
  input logic [63:0] data_in,
  input logic [63:0] data_in_bit_sel,
  input logic ren,
  input logic reset,
  input logic wen,
  output logic [63:0] data_out
);

logic glb_bank_sram_gen_CEB;
logic glb_bank_sram_gen_WEB;
logic [13:0] sram_addr;
logic [13:0] sram_addr_d;
logic sram_cen;
logic sram_cen_d;
logic [63:0] sram_data_in;
logic [63:0] sram_data_in_bit_sel;
logic [63:0] sram_data_in_bit_sel_d;
logic [63:0] sram_data_in_d;
logic [63:0] sram_data_out;
logic [143:0] sram_signals_pipeline_in_;
logic [143:0] sram_signals_pipeline_out_;
logic sram_wen;
logic sram_wen_d;
assign sram_signals_pipeline_in_ = {sram_wen, sram_cen, sram_addr, sram_data_in, sram_data_in_bit_sel};
assign {sram_wen_d, sram_cen_d, sram_addr_d, sram_data_in_d, sram_data_in_bit_sel_d} = sram_signals_pipeline_out_;
assign glb_bank_sram_gen_CEB = ~sram_cen_d;
assign glb_bank_sram_gen_WEB = ~sram_wen_d;
always_comb begin
  sram_wen = wen;
  sram_cen = wen | ren;
  sram_addr = addr[16:3];
  sram_data_in = data_in;
  sram_data_in_bit_sel = data_in_bit_sel;
  data_out = sram_data_out;
end
pipeline_w_144_d_0 sram_signals_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(sram_signals_pipeline_in_),
  .reset(reset),
  .out_(sram_signals_pipeline_out_)
);

glb_bank_sram_gen glb_bank_sram_gen (
  .A(sram_addr_d),
  .BW(sram_data_in_bit_sel_d),
  .CEB(glb_bank_sram_gen_CEB),
  .CLK(clk),
  .D(sram_data_in_d),
  .RESET(reset),
  .WEB(glb_bank_sram_gen_WEB),
  .Q(sram_data_out)
);

endmodule   // glb_bank_memory

module glb_bank_mux (
  input logic cfg_pcfg_tile_connected_next,
  input logic cfg_pcfg_tile_connected_prev,
  input logic cfg_tile_connected_next,
  input logic cfg_tile_connected_prev,
  input logic clk,
  input logic glb_tile_id,
  input rdrq_packet_t rdrq_packet_dma2bank,
  input rdrq_packet_t rdrq_packet_pcfgdma2bank,
  input rdrq_packet_t rdrq_packet_pcfgring2bank,
  input rdrq_packet_t rdrq_packet_procsw2bank,
  input rdrq_packet_t rdrq_packet_ring2bank,
  input rdrs_packet_t [1:0] rdrs_packet_bankarr2sw,
  input logic reset,
  input wr_packet_t wr_packet_dma2bank,
  input wr_packet_t wr_packet_procsw2bank,
  input wr_packet_t wr_packet_ring2bank,
  output rdrq_bank_packet_t [1:0] rdrq_packet_sw2bankarr,
  output rdrs_packet_t rdrs_packet_bank2dma,
  output rdrs_packet_t rdrs_packet_bank2pcfgdma,
  output rdrs_packet_t rdrs_packet_bank2pcfgring,
  output rdrs_packet_t rdrs_packet_bank2procsw,
  output rdrs_packet_t rdrs_packet_bank2ring,
  output wr_bank_packet_t [1:0] wr_packet_sw2bankarr
);

typedef enum logic[1:0] {
  none = 2'h0,
  proc = 2'h1,
  strm = 2'h2,
  pcfg = 2'h3
} rd_type_e;
rd_type_e rd_type_0;
rd_type_e rd_type_1;
rd_type_e rd_type_d_0;
rd_type_e rd_type_d_1;
logic [3:0] rd_type_pipeline_1_in_;
logic [3:0] rd_type_pipeline_1_out_;
rdrq_bank_packet_t [1:0] rdrq_packet_sw2bankarr_w;
logic [17:0] rdrq_sw2bank_pipeline_0_out_;
logic [17:0] rdrq_sw2bank_pipeline_1_out_;
logic [64:0] rdrs_bank2sw_pipeline_0_out_;
logic [64:0] rdrs_bank2sw_pipeline_1_out_;
rdrs_packet_t [1:0] rdrs_packet_bankarr2sw_d;
wr_bank_packet_t [1:0] wr_packet_sw2bankarr_w;
logic [89:0] wr_sw2bank_pipeline_0_out_;
logic [89:0] wr_sw2bank_pipeline_1_out_;
assign wr_packet_sw2bankarr[0] = wr_sw2bank_pipeline_0_out_;
assign wr_packet_sw2bankarr[1] = wr_sw2bank_pipeline_1_out_;
assign rdrq_packet_sw2bankarr[0] = rdrq_sw2bank_pipeline_0_out_;
assign rdrq_packet_sw2bankarr[1] = rdrq_sw2bank_pipeline_1_out_;
assign rd_type_pipeline_1_in_ = {rd_type_0, rd_type_1};
assign {rd_type_d_0, rd_type_d_1} = rd_type_pipeline_1_out_;
assign rdrs_packet_bankarr2sw_d[0] = rdrs_bank2sw_pipeline_0_out_;
assign rdrs_packet_bankarr2sw_d[1] = rdrs_bank2sw_pipeline_1_out_;
always_comb begin
  if ((wr_packet_procsw2bank.wr_en == 1'h1) & (wr_packet_procsw2bank.wr_addr[18] == glb_tile_id) & (wr_packet_procsw2bank.wr_addr[17] == 1'h0)) begin
    wr_packet_sw2bankarr_w[0].wr_en = wr_packet_procsw2bank.wr_en;
    wr_packet_sw2bankarr_w[0].wr_addr = wr_packet_procsw2bank.wr_addr[16:0];
    wr_packet_sw2bankarr_w[0].wr_strb = wr_packet_procsw2bank.wr_strb;
    wr_packet_sw2bankarr_w[0].wr_data = wr_packet_procsw2bank.wr_data;
  end
  else if ((wr_packet_dma2bank.wr_en == 1'h1) & (~cfg_tile_connected_prev) & (~cfg_tile_connected_next) & (wr_packet_dma2bank.wr_addr[18] == glb_tile_id) & (wr_packet_dma2bank.wr_addr[17] == 1'h0)) begin
    wr_packet_sw2bankarr_w[0].wr_en = wr_packet_dma2bank.wr_en;
    wr_packet_sw2bankarr_w[0].wr_addr = wr_packet_dma2bank.wr_addr[16:0];
    wr_packet_sw2bankarr_w[0].wr_strb = wr_packet_dma2bank.wr_strb;
    wr_packet_sw2bankarr_w[0].wr_data = wr_packet_dma2bank.wr_data;
  end
  else if ((wr_packet_ring2bank.wr_en == 1'h1) & (wr_packet_ring2bank.wr_addr[18] == glb_tile_id) & (wr_packet_ring2bank.wr_addr[17] == 1'h0)) begin
    wr_packet_sw2bankarr_w[0].wr_en = wr_packet_ring2bank.wr_en;
    wr_packet_sw2bankarr_w[0].wr_addr = wr_packet_ring2bank.wr_addr[16:0];
    wr_packet_sw2bankarr_w[0].wr_strb = wr_packet_ring2bank.wr_strb;
    wr_packet_sw2bankarr_w[0].wr_data = wr_packet_ring2bank.wr_data;
  end
  else wr_packet_sw2bankarr_w[0] = 90'h0;
end
always_comb begin
  if ((wr_packet_procsw2bank.wr_en == 1'h1) & (wr_packet_procsw2bank.wr_addr[18] == glb_tile_id) & (wr_packet_procsw2bank.wr_addr[17] == 1'h1)) begin
    wr_packet_sw2bankarr_w[1].wr_en = wr_packet_procsw2bank.wr_en;
    wr_packet_sw2bankarr_w[1].wr_addr = wr_packet_procsw2bank.wr_addr[16:0];
    wr_packet_sw2bankarr_w[1].wr_strb = wr_packet_procsw2bank.wr_strb;
    wr_packet_sw2bankarr_w[1].wr_data = wr_packet_procsw2bank.wr_data;
  end
  else if ((wr_packet_dma2bank.wr_en == 1'h1) & (~cfg_tile_connected_prev) & (~cfg_tile_connected_next) & (wr_packet_dma2bank.wr_addr[18] == glb_tile_id) & (wr_packet_dma2bank.wr_addr[17] == 1'h1)) begin
    wr_packet_sw2bankarr_w[1].wr_en = wr_packet_dma2bank.wr_en;
    wr_packet_sw2bankarr_w[1].wr_addr = wr_packet_dma2bank.wr_addr[16:0];
    wr_packet_sw2bankarr_w[1].wr_strb = wr_packet_dma2bank.wr_strb;
    wr_packet_sw2bankarr_w[1].wr_data = wr_packet_dma2bank.wr_data;
  end
  else if ((wr_packet_ring2bank.wr_en == 1'h1) & (wr_packet_ring2bank.wr_addr[18] == glb_tile_id) & (wr_packet_ring2bank.wr_addr[17] == 1'h1)) begin
    wr_packet_sw2bankarr_w[1].wr_en = wr_packet_ring2bank.wr_en;
    wr_packet_sw2bankarr_w[1].wr_addr = wr_packet_ring2bank.wr_addr[16:0];
    wr_packet_sw2bankarr_w[1].wr_strb = wr_packet_ring2bank.wr_strb;
    wr_packet_sw2bankarr_w[1].wr_data = wr_packet_ring2bank.wr_data;
  end
  else wr_packet_sw2bankarr_w[1] = 90'h0;
end
always_comb begin
  if ((rdrq_packet_procsw2bank.rd_en == 1'h1) & (rdrq_packet_procsw2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_procsw2bank.rd_addr[17] == 1'h0)) begin
    rdrq_packet_sw2bankarr_w[0].rd_en = rdrq_packet_procsw2bank.rd_en;
    rdrq_packet_sw2bankarr_w[0].rd_addr = rdrq_packet_procsw2bank.rd_addr[16:0];
    rd_type_0 = proc;
  end
  else if ((rdrq_packet_pcfgdma2bank.rd_en == 1'h1) & (~cfg_pcfg_tile_connected_prev) & (~cfg_pcfg_tile_connected_next) & (rdrq_packet_pcfgdma2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_pcfgdma2bank.rd_addr[17] == 1'h0)) begin
    rdrq_packet_sw2bankarr_w[0].rd_en = rdrq_packet_pcfgdma2bank.rd_en;
    rdrq_packet_sw2bankarr_w[0].rd_addr = rdrq_packet_pcfgdma2bank.rd_addr[16:0];
    rd_type_0 = pcfg;
  end
  else if ((rdrq_packet_pcfgring2bank.rd_en == 1'h1) & (rdrq_packet_pcfgring2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_pcfgring2bank.rd_addr[17] == 1'h0)) begin
    rdrq_packet_sw2bankarr_w[0].rd_en = rdrq_packet_pcfgring2bank.rd_en;
    rdrq_packet_sw2bankarr_w[0].rd_addr = rdrq_packet_pcfgring2bank.rd_addr[16:0];
    rd_type_0 = pcfg;
  end
  else if ((rdrq_packet_dma2bank.rd_en == 1'h1) & (~cfg_tile_connected_prev) & (~cfg_tile_connected_next) & (rdrq_packet_dma2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_dma2bank.rd_addr[17] == 1'h0)) begin
    rdrq_packet_sw2bankarr_w[0].rd_en = rdrq_packet_dma2bank.rd_en;
    rdrq_packet_sw2bankarr_w[0].rd_addr = rdrq_packet_dma2bank.rd_addr[16:0];
    rd_type_0 = strm;
  end
  else if ((rdrq_packet_ring2bank.rd_en == 1'h1) & (rdrq_packet_ring2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_ring2bank.rd_addr[17] == 1'h0)) begin
    rdrq_packet_sw2bankarr_w[0].rd_en = rdrq_packet_ring2bank.rd_en;
    rdrq_packet_sw2bankarr_w[0].rd_addr = rdrq_packet_ring2bank.rd_addr[16:0];
    rd_type_0 = strm;
  end
  else begin
    rdrq_packet_sw2bankarr_w[0] = 18'h0;
    rd_type_0 = none;
  end
end
always_comb begin
  if ((rdrq_packet_procsw2bank.rd_en == 1'h1) & (rdrq_packet_procsw2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_procsw2bank.rd_addr[17] == 1'h1)) begin
    rdrq_packet_sw2bankarr_w[1].rd_en = rdrq_packet_procsw2bank.rd_en;
    rdrq_packet_sw2bankarr_w[1].rd_addr = rdrq_packet_procsw2bank.rd_addr[16:0];
    rd_type_1 = proc;
  end
  else if ((rdrq_packet_pcfgdma2bank.rd_en == 1'h1) & (~cfg_pcfg_tile_connected_prev) & (~cfg_pcfg_tile_connected_next) & (rdrq_packet_pcfgdma2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_pcfgdma2bank.rd_addr[17] == 1'h1)) begin
    rdrq_packet_sw2bankarr_w[1].rd_en = rdrq_packet_pcfgdma2bank.rd_en;
    rdrq_packet_sw2bankarr_w[1].rd_addr = rdrq_packet_pcfgdma2bank.rd_addr[16:0];
    rd_type_1 = pcfg;
  end
  else if ((rdrq_packet_pcfgring2bank.rd_en == 1'h1) & (rdrq_packet_pcfgring2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_pcfgring2bank.rd_addr[17] == 1'h1)) begin
    rdrq_packet_sw2bankarr_w[1].rd_en = rdrq_packet_pcfgring2bank.rd_en;
    rdrq_packet_sw2bankarr_w[1].rd_addr = rdrq_packet_pcfgring2bank.rd_addr[16:0];
    rd_type_1 = pcfg;
  end
  else if ((rdrq_packet_dma2bank.rd_en == 1'h1) & (~cfg_tile_connected_prev) & (~cfg_tile_connected_next) & (rdrq_packet_dma2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_dma2bank.rd_addr[17] == 1'h1)) begin
    rdrq_packet_sw2bankarr_w[1].rd_en = rdrq_packet_dma2bank.rd_en;
    rdrq_packet_sw2bankarr_w[1].rd_addr = rdrq_packet_dma2bank.rd_addr[16:0];
    rd_type_1 = strm;
  end
  else if ((rdrq_packet_ring2bank.rd_en == 1'h1) & (rdrq_packet_ring2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_ring2bank.rd_addr[17] == 1'h1)) begin
    rdrq_packet_sw2bankarr_w[1].rd_en = rdrq_packet_ring2bank.rd_en;
    rdrq_packet_sw2bankarr_w[1].rd_addr = rdrq_packet_ring2bank.rd_addr[16:0];
    rd_type_1 = strm;
  end
  else begin
    rdrq_packet_sw2bankarr_w[1] = 18'h0;
    rd_type_1 = none;
  end
end
always_comb begin
  rdrs_packet_bank2dma = 65'h0;
  if ((~cfg_tile_connected_next) & (~cfg_tile_connected_prev)) begin
    if (rd_type_d_0 == strm) begin
      rdrs_packet_bank2dma = rdrs_packet_bankarr2sw_d[0];
    end
    if (rd_type_d_1 == strm) begin
      rdrs_packet_bank2dma = rdrs_packet_bankarr2sw_d[1];
    end
  end
end
always_comb begin
  rdrs_packet_bank2ring = 65'h0;
  if (cfg_tile_connected_next | cfg_tile_connected_prev) begin
    if (rd_type_d_0 == strm) begin
      rdrs_packet_bank2ring = rdrs_packet_bankarr2sw_d[0];
    end
    if (rd_type_d_1 == strm) begin
      rdrs_packet_bank2ring = rdrs_packet_bankarr2sw_d[1];
    end
  end
end
always_comb begin
  rdrs_packet_bank2procsw = 65'h0;
  if (rd_type_d_0 == proc) begin
    rdrs_packet_bank2procsw = rdrs_packet_bankarr2sw_d[0];
  end
  if (rd_type_d_1 == proc) begin
    rdrs_packet_bank2procsw = rdrs_packet_bankarr2sw_d[1];
  end
end
always_comb begin
  rdrs_packet_bank2pcfgdma = 65'h0;
  if ((~cfg_pcfg_tile_connected_next) & (~cfg_pcfg_tile_connected_prev)) begin
    if (rd_type_d_0 == pcfg) begin
      rdrs_packet_bank2pcfgdma = rdrs_packet_bankarr2sw_d[0];
    end
    if (rd_type_d_1 == pcfg) begin
      rdrs_packet_bank2pcfgdma = rdrs_packet_bankarr2sw_d[1];
    end
  end
end
always_comb begin
  rdrs_packet_bank2pcfgring = 65'h0;
  if (cfg_pcfg_tile_connected_next | cfg_pcfg_tile_connected_prev) begin
    if (rd_type_d_0 == pcfg) begin
      rdrs_packet_bank2pcfgring = rdrs_packet_bankarr2sw_d[0];
    end
    if (rd_type_d_1 == pcfg) begin
      rdrs_packet_bank2pcfgring = rdrs_packet_bankarr2sw_d[1];
    end
  end
end
pipeline_w_90_d_0 wr_sw2bank_pipeline_0 (
  .clk(clk),
  .clk_en(1'h1),
  .in_(wr_packet_sw2bankarr_w[0]),
  .reset(reset),
  .out_(wr_sw2bank_pipeline_0_out_)
);

pipeline_w_90_d_0 wr_sw2bank_pipeline_1 (
  .clk(clk),
  .clk_en(1'h1),
  .in_(wr_packet_sw2bankarr_w[1]),
  .reset(reset),
  .out_(wr_sw2bank_pipeline_1_out_)
);

pipeline_w_18_d_0 rdrq_sw2bank_pipeline_0 (
  .clk(clk),
  .clk_en(1'h1),
  .in_(rdrq_packet_sw2bankarr_w[0]),
  .reset(reset),
  .out_(rdrq_sw2bank_pipeline_0_out_)
);

pipeline_w_18_d_0 rdrq_sw2bank_pipeline_1 (
  .clk(clk),
  .clk_en(1'h1),
  .in_(rdrq_packet_sw2bankarr_w[1]),
  .reset(reset),
  .out_(rdrq_sw2bank_pipeline_1_out_)
);

pipeline_w_4_d_2 rd_type_pipeline_1 (
  .clk(clk),
  .clk_en(1'h1),
  .in_(rd_type_pipeline_1_in_),
  .reset(reset),
  .out_(rd_type_pipeline_1_out_)
);

pipeline_w_65_d_1 rdrs_bank2sw_pipeline_0 (
  .clk(clk),
  .clk_en(1'h1),
  .in_(rdrs_packet_bankarr2sw[0]),
  .reset(reset),
  .out_(rdrs_bank2sw_pipeline_0_out_)
);

pipeline_w_65_d_1 rdrs_bank2sw_pipeline_1 (
  .clk(clk),
  .clk_en(1'h1),
  .in_(rdrs_packet_bankarr2sw[1]),
  .reset(reset),
  .out_(rdrs_bank2sw_pipeline_1_out_)
);

endmodule   // glb_bank_mux

module glb_bank_sram_gen (
  input logic [13:0] A,
  input logic [63:0] BW,
  input logic CEB,
  input logic CLK,
  input logic [63:0] D,
  input logic RESET,
  input logic WEB,
  output logic [63:0] Q
);

logic [11:0] A_SRAM;
logic [11:0] A_SRAM_d;
logic [63:0] BW_d;
logic [3:0] CEB_DEMUX;
logic [3:0] CEB_DEMUX_d;
logic CEB_d;
logic [63:0] D_d;
logic [1:0] Q_SEL;
logic [63:0] Q_SRAM2MUX [3:0];
logic [63:0] Q_w;
logic [1:0] SRAM_SEL;
logic [1:0] SRAM_SEL_d;
logic [3:0] WEB_DEMUX;
logic [3:0] WEB_DEMUX_d;
logic WEB_d;
logic [63:0] sram_array_0_Q;
logic [63:0] sram_array_1_Q;
logic [63:0] sram_array_2_Q;
logic [63:0] sram_array_3_Q;
logic [77:0] sram_signals_pipeline_in_;
logic [77:0] sram_signals_pipeline_out_;
logic [73:0] sram_signals_reset_high_pipeline_in_;
logic [73:0] sram_signals_reset_high_pipeline_out_;
assign SRAM_SEL = A[13:12];
assign A_SRAM = A[11:0];
assign sram_signals_reset_high_pipeline_in_ = {WEB, CEB, WEB_DEMUX, CEB_DEMUX, BW};
assign {WEB_d, CEB_d, WEB_DEMUX_d, CEB_DEMUX_d, BW_d} = sram_signals_reset_high_pipeline_out_;
assign sram_signals_pipeline_in_ = {A_SRAM, SRAM_SEL, D};
assign {A_SRAM_d, SRAM_SEL_d, D_d} = sram_signals_pipeline_out_;

always_ff @(posedge CLK, posedge RESET) begin
  if (RESET) begin
    Q_SEL <= 2'h0;
  end
  else if ((CEB_d == 1'h0) & (WEB_d == 1'h1)) begin
    Q_SEL <= SRAM_SEL_d;
  end
end
always_comb begin
  if (~WEB) begin
    WEB_DEMUX = ~(4'h1 << 4'(SRAM_SEL));
  end
  else WEB_DEMUX = 4'hF;
  if (~CEB) begin
    CEB_DEMUX = ~(4'h1 << 4'(SRAM_SEL));
  end
  else CEB_DEMUX = 4'hF;
end
assign Q_SRAM2MUX[0] = sram_array_0_Q;
assign Q_SRAM2MUX[1] = sram_array_1_Q;
assign Q_SRAM2MUX[2] = sram_array_2_Q;
assign Q_SRAM2MUX[3] = sram_array_3_Q;
assign Q_w = Q_SRAM2MUX[Q_SEL];
pipeline_w_74_d_0_reset_high sram_signals_reset_high_pipeline (
  .clk(CLK),
  .clk_en(1'h1),
  .in_(sram_signals_reset_high_pipeline_in_),
  .reset(RESET),
  .out_(sram_signals_reset_high_pipeline_out_)
);

pipeline_w_78_d_0 sram_signals_pipeline (
  .clk(CLK),
  .clk_en(1'h1),
  .in_(sram_signals_pipeline_in_),
  .reset(RESET),
  .out_(sram_signals_pipeline_out_)
);

pipeline_w_64_d_0 sram_signals_output_pipeline (
  .clk(CLK),
  .clk_en(1'h1),
  .in_(Q_w),
  .reset(RESET),
  .out_(Q)
);

IN12LP_S1DB_W04096B064M08S2_HB sram_array_0 (
  .A(A_SRAM_d),
  .BW(BW_d),
  .CEN(CEB_DEMUX_d[0]),
  .CLK(CLK),
  .D(D_d),
  .MA_SAWL0(1'h0),
  .MA_SAWL1(1'h0),
  .MA_STABAS0(1'h0),
  .MA_STABAS1(1'h0),
  .MA_VD0(1'h0),
  .MA_VD1(1'h0),
  .MA_WL0(1'h0),
  .MA_WL1(1'h0),
  .MA_WRAS0(1'h0),
  .MA_WRAS1(1'h0),
  .MA_WRT(1'h0),
  .RDWEN(WEB_DEMUX_d[0]),
  .T_LOGIC(1'h0),
  .T_Q_RST(1'h0),
  .Q(sram_array_0_Q)
);

IN12LP_S1DB_W04096B064M08S2_HB sram_array_1 (
  .A(A_SRAM_d),
  .BW(BW_d),
  .CEN(CEB_DEMUX_d[1]),
  .CLK(CLK),
  .D(D_d),
  .MA_SAWL0(1'h0),
  .MA_SAWL1(1'h0),
  .MA_STABAS0(1'h0),
  .MA_STABAS1(1'h0),
  .MA_VD0(1'h0),
  .MA_VD1(1'h0),
  .MA_WL0(1'h0),
  .MA_WL1(1'h0),
  .MA_WRAS0(1'h0),
  .MA_WRAS1(1'h0),
  .MA_WRT(1'h0),
  .RDWEN(WEB_DEMUX_d[1]),
  .T_LOGIC(1'h0),
  .T_Q_RST(1'h0),
  .Q(sram_array_1_Q)
);

IN12LP_S1DB_W04096B064M08S2_HB sram_array_2 (
  .A(A_SRAM_d),
  .BW(BW_d),
  .CEN(CEB_DEMUX_d[2]),
  .CLK(CLK),
  .D(D_d),
  .MA_SAWL0(1'h0),
  .MA_SAWL1(1'h0),
  .MA_STABAS0(1'h0),
  .MA_STABAS1(1'h0),
  .MA_VD0(1'h0),
  .MA_VD1(1'h0),
  .MA_WL0(1'h0),
  .MA_WL1(1'h0),
  .MA_WRAS0(1'h0),
  .MA_WRAS1(1'h0),
  .MA_WRT(1'h0),
  .RDWEN(WEB_DEMUX_d[2]),
  .T_LOGIC(1'h0),
  .T_Q_RST(1'h0),
  .Q(sram_array_2_Q)
);

IN12LP_S1DB_W04096B064M08S2_HB sram_array_3 (
  .A(A_SRAM_d),
  .BW(BW_d),
  .CEN(CEB_DEMUX_d[3]),
  .CLK(CLK),
  .D(D_d),
  .MA_SAWL0(1'h0),
  .MA_SAWL1(1'h0),
  .MA_STABAS0(1'h0),
  .MA_STABAS1(1'h0),
  .MA_VD0(1'h0),
  .MA_VD1(1'h0),
  .MA_WL0(1'h0),
  .MA_WL1(1'h0),
  .MA_WRAS0(1'h0),
  .MA_WRAS1(1'h0),
  .MA_WRT(1'h0),
  .RDWEN(WEB_DEMUX_d[3]),
  .T_LOGIC(1'h0),
  .T_Q_RST(1'h0),
  .Q(sram_array_3_Q)
);

endmodule   // glb_bank_sram_gen

module glb_cfg (
  glb_tile_ifc_A_12_D_32.master if_cfg_est_m,
  glb_tile_ifc_A_12_D_32.slave if_cfg_wst_s,
  input logic gclk,
  input logic glb_tile_id,
  input logic mclk,
  input logic reset,
  output cfg_data_network_t cfg_data_network,
  output load_dma_ctrl_t cfg_ld_dma_ctrl,
  output dma_header_t cfg_ld_dma_header,
  output pcfg_broadcast_mux_t cfg_pcfg_broadcast_mux,
  output pcfg_dma_ctrl_t cfg_pcfg_dma_ctrl,
  output pcfg_dma_header_t cfg_pcfg_dma_header,
  output cfg_pcfg_network_t cfg_pcfg_network,
  output store_dma_ctrl_t cfg_st_dma_ctrl,
  output dma_header_t cfg_st_dma_header
);

logic [8:0] glb_cfg_ctrl_h2d_pio_dec_address;
logic glb_pio_d2h_dec_pio_ack;
logic glb_pio_d2h_dec_pio_nack;
logic [31:0] glb_pio_d2h_dec_pio_read_data;
logic [5:0] glb_pio_h2d_pio_dec_address;
logic glb_pio_h2d_pio_dec_read;
logic glb_pio_h2d_pio_dec_write;
logic [31:0] glb_pio_h2d_pio_dec_write_data;
logic glb_pio_l2h_data_network_ctrl_connected_r;
logic [5:0] glb_pio_l2h_data_network_latency_value_r;
logic [1:0] glb_pio_l2h_ld_dma_ctrl_data_mux_r;
logic [1:0] glb_pio_l2h_ld_dma_ctrl_mode_r;
logic glb_pio_l2h_ld_dma_ctrl_num_repeat_r;
logic glb_pio_l2h_ld_dma_ctrl_use_flush_r;
logic glb_pio_l2h_ld_dma_ctrl_use_valid_r;
logic [15:0] glb_pio_l2h_ld_dma_header_0_cycle_start_addr_cycle_start_addr_r;
logic [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_0_cycle_stride_r;
logic [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_1_cycle_stride_r;
logic [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_2_cycle_stride_r;
logic [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_3_cycle_stride_r;
logic [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_4_cycle_stride_r;
logic [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_5_cycle_stride_r;
logic [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_6_cycle_stride_r;
logic [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_7_cycle_stride_r;
logic [3:0] glb_pio_l2h_ld_dma_header_0_dim_dim_r;
logic [31:0] glb_pio_l2h_ld_dma_header_0_range_0_range_r;
logic [31:0] glb_pio_l2h_ld_dma_header_0_range_1_range_r;
logic [31:0] glb_pio_l2h_ld_dma_header_0_range_2_range_r;
logic [31:0] glb_pio_l2h_ld_dma_header_0_range_3_range_r;
logic [31:0] glb_pio_l2h_ld_dma_header_0_range_4_range_r;
logic [31:0] glb_pio_l2h_ld_dma_header_0_range_5_range_r;
logic [31:0] glb_pio_l2h_ld_dma_header_0_range_6_range_r;
logic [31:0] glb_pio_l2h_ld_dma_header_0_range_7_range_r;
logic [18:0] glb_pio_l2h_ld_dma_header_0_start_addr_start_addr_r;
logic [19:0] glb_pio_l2h_ld_dma_header_0_stride_0_stride_r;
logic [19:0] glb_pio_l2h_ld_dma_header_0_stride_1_stride_r;
logic [19:0] glb_pio_l2h_ld_dma_header_0_stride_2_stride_r;
logic [19:0] glb_pio_l2h_ld_dma_header_0_stride_3_stride_r;
logic [19:0] glb_pio_l2h_ld_dma_header_0_stride_4_stride_r;
logic [19:0] glb_pio_l2h_ld_dma_header_0_stride_5_stride_r;
logic [19:0] glb_pio_l2h_ld_dma_header_0_stride_6_stride_r;
logic [19:0] glb_pio_l2h_ld_dma_header_0_stride_7_stride_r;
logic [1:0] glb_pio_l2h_pcfg_broadcast_mux_east_r;
logic [1:0] glb_pio_l2h_pcfg_broadcast_mux_south_r;
logic [1:0] glb_pio_l2h_pcfg_broadcast_mux_west_r;
logic glb_pio_l2h_pcfg_dma_ctrl_mode_r;
logic glb_pio_l2h_pcfg_dma_ctrl_relocation_is_msb_r;
logic [15:0] glb_pio_l2h_pcfg_dma_ctrl_relocation_value_r;
logic [15:0] glb_pio_l2h_pcfg_dma_header_num_cfg_num_cfg_r;
logic [18:0] glb_pio_l2h_pcfg_dma_header_start_addr_start_addr_r;
logic glb_pio_l2h_pcfg_network_ctrl_connected_r;
logic [5:0] glb_pio_l2h_pcfg_network_latency_value_r;
logic [1:0] glb_pio_l2h_st_dma_ctrl_data_mux_r;
logic [1:0] glb_pio_l2h_st_dma_ctrl_mode_r;
logic glb_pio_l2h_st_dma_ctrl_num_repeat_r;
logic glb_pio_l2h_st_dma_ctrl_use_valid_r;
logic [15:0] glb_pio_l2h_st_dma_header_0_cycle_start_addr_cycle_start_addr_r;
logic [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_0_cycle_stride_r;
logic [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_1_cycle_stride_r;
logic [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_2_cycle_stride_r;
logic [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_3_cycle_stride_r;
logic [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_4_cycle_stride_r;
logic [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_5_cycle_stride_r;
logic [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_6_cycle_stride_r;
logic [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_7_cycle_stride_r;
logic [3:0] glb_pio_l2h_st_dma_header_0_dim_dim_r;
logic [31:0] glb_pio_l2h_st_dma_header_0_range_0_range_r;
logic [31:0] glb_pio_l2h_st_dma_header_0_range_1_range_r;
logic [31:0] glb_pio_l2h_st_dma_header_0_range_2_range_r;
logic [31:0] glb_pio_l2h_st_dma_header_0_range_3_range_r;
logic [31:0] glb_pio_l2h_st_dma_header_0_range_4_range_r;
logic [31:0] glb_pio_l2h_st_dma_header_0_range_5_range_r;
logic [31:0] glb_pio_l2h_st_dma_header_0_range_6_range_r;
logic [31:0] glb_pio_l2h_st_dma_header_0_range_7_range_r;
logic [18:0] glb_pio_l2h_st_dma_header_0_start_addr_start_addr_r;
logic [19:0] glb_pio_l2h_st_dma_header_0_stride_0_stride_r;
logic [19:0] glb_pio_l2h_st_dma_header_0_stride_1_stride_r;
logic [19:0] glb_pio_l2h_st_dma_header_0_stride_2_stride_r;
logic [19:0] glb_pio_l2h_st_dma_header_0_stride_3_stride_r;
logic [19:0] glb_pio_l2h_st_dma_header_0_stride_4_stride_r;
logic [19:0] glb_pio_l2h_st_dma_header_0_stride_5_stride_r;
logic [19:0] glb_pio_l2h_st_dma_header_0_stride_6_stride_r;
logic [19:0] glb_pio_l2h_st_dma_header_0_stride_7_stride_r;
assign cfg_data_network.tile_connected = glb_pio_l2h_data_network_ctrl_connected_r;
assign cfg_data_network.latency = glb_pio_l2h_data_network_latency_value_r;
assign cfg_pcfg_network.tile_connected = glb_pio_l2h_pcfg_network_ctrl_connected_r;
assign cfg_pcfg_network.latency = glb_pio_l2h_pcfg_network_latency_value_r;
assign cfg_st_dma_ctrl.data_mux = glb_pio_l2h_st_dma_ctrl_data_mux_r;
assign cfg_st_dma_ctrl.mode = glb_pio_l2h_st_dma_ctrl_mode_r;
assign cfg_st_dma_ctrl.use_valid = glb_pio_l2h_st_dma_ctrl_use_valid_r;
assign cfg_st_dma_ctrl.num_repeat = glb_pio_l2h_st_dma_ctrl_num_repeat_r;
assign cfg_st_dma_header.start_addr = glb_pio_l2h_st_dma_header_0_start_addr_start_addr_r;
assign cfg_st_dma_header.cycle_start_addr = glb_pio_l2h_st_dma_header_0_cycle_start_addr_cycle_start_addr_r;
assign cfg_st_dma_header.dim = glb_pio_l2h_st_dma_header_0_dim_dim_r;
assign cfg_st_dma_header.cycle_stride_0 = glb_pio_l2h_st_dma_header_0_cycle_stride_0_cycle_stride_r;
assign cfg_st_dma_header.stride_0 = glb_pio_l2h_st_dma_header_0_stride_0_stride_r;
assign cfg_st_dma_header.range_0 = glb_pio_l2h_st_dma_header_0_range_0_range_r;
assign cfg_st_dma_header.cycle_stride_1 = glb_pio_l2h_st_dma_header_0_cycle_stride_1_cycle_stride_r;
assign cfg_st_dma_header.stride_1 = glb_pio_l2h_st_dma_header_0_stride_1_stride_r;
assign cfg_st_dma_header.range_1 = glb_pio_l2h_st_dma_header_0_range_1_range_r;
assign cfg_st_dma_header.cycle_stride_2 = glb_pio_l2h_st_dma_header_0_cycle_stride_2_cycle_stride_r;
assign cfg_st_dma_header.stride_2 = glb_pio_l2h_st_dma_header_0_stride_2_stride_r;
assign cfg_st_dma_header.range_2 = glb_pio_l2h_st_dma_header_0_range_2_range_r;
assign cfg_st_dma_header.cycle_stride_3 = glb_pio_l2h_st_dma_header_0_cycle_stride_3_cycle_stride_r;
assign cfg_st_dma_header.stride_3 = glb_pio_l2h_st_dma_header_0_stride_3_stride_r;
assign cfg_st_dma_header.range_3 = glb_pio_l2h_st_dma_header_0_range_3_range_r;
assign cfg_st_dma_header.cycle_stride_4 = glb_pio_l2h_st_dma_header_0_cycle_stride_4_cycle_stride_r;
assign cfg_st_dma_header.stride_4 = glb_pio_l2h_st_dma_header_0_stride_4_stride_r;
assign cfg_st_dma_header.range_4 = glb_pio_l2h_st_dma_header_0_range_4_range_r;
assign cfg_st_dma_header.cycle_stride_5 = glb_pio_l2h_st_dma_header_0_cycle_stride_5_cycle_stride_r;
assign cfg_st_dma_header.stride_5 = glb_pio_l2h_st_dma_header_0_stride_5_stride_r;
assign cfg_st_dma_header.range_5 = glb_pio_l2h_st_dma_header_0_range_5_range_r;
assign cfg_st_dma_header.cycle_stride_6 = glb_pio_l2h_st_dma_header_0_cycle_stride_6_cycle_stride_r;
assign cfg_st_dma_header.stride_6 = glb_pio_l2h_st_dma_header_0_stride_6_stride_r;
assign cfg_st_dma_header.range_6 = glb_pio_l2h_st_dma_header_0_range_6_range_r;
assign cfg_st_dma_header.cycle_stride_7 = glb_pio_l2h_st_dma_header_0_cycle_stride_7_cycle_stride_r;
assign cfg_st_dma_header.stride_7 = glb_pio_l2h_st_dma_header_0_stride_7_stride_r;
assign cfg_st_dma_header.range_7 = glb_pio_l2h_st_dma_header_0_range_7_range_r;
assign cfg_ld_dma_ctrl.data_mux = glb_pio_l2h_ld_dma_ctrl_data_mux_r;
assign cfg_ld_dma_ctrl.mode = glb_pio_l2h_ld_dma_ctrl_mode_r;
assign cfg_ld_dma_ctrl.use_valid = glb_pio_l2h_ld_dma_ctrl_use_valid_r;
assign cfg_ld_dma_ctrl.use_flush = glb_pio_l2h_ld_dma_ctrl_use_flush_r;
assign cfg_ld_dma_ctrl.num_repeat = glb_pio_l2h_ld_dma_ctrl_num_repeat_r;
assign cfg_ld_dma_header.start_addr = glb_pio_l2h_ld_dma_header_0_start_addr_start_addr_r;
assign cfg_ld_dma_header.cycle_start_addr = glb_pio_l2h_ld_dma_header_0_cycle_start_addr_cycle_start_addr_r;
assign cfg_ld_dma_header.dim = glb_pio_l2h_ld_dma_header_0_dim_dim_r;
assign cfg_ld_dma_header.cycle_stride_0 = glb_pio_l2h_ld_dma_header_0_cycle_stride_0_cycle_stride_r;
assign cfg_ld_dma_header.stride_0 = glb_pio_l2h_ld_dma_header_0_stride_0_stride_r;
assign cfg_ld_dma_header.range_0 = glb_pio_l2h_ld_dma_header_0_range_0_range_r;
assign cfg_ld_dma_header.cycle_stride_1 = glb_pio_l2h_ld_dma_header_0_cycle_stride_1_cycle_stride_r;
assign cfg_ld_dma_header.stride_1 = glb_pio_l2h_ld_dma_header_0_stride_1_stride_r;
assign cfg_ld_dma_header.range_1 = glb_pio_l2h_ld_dma_header_0_range_1_range_r;
assign cfg_ld_dma_header.cycle_stride_2 = glb_pio_l2h_ld_dma_header_0_cycle_stride_2_cycle_stride_r;
assign cfg_ld_dma_header.stride_2 = glb_pio_l2h_ld_dma_header_0_stride_2_stride_r;
assign cfg_ld_dma_header.range_2 = glb_pio_l2h_ld_dma_header_0_range_2_range_r;
assign cfg_ld_dma_header.cycle_stride_3 = glb_pio_l2h_ld_dma_header_0_cycle_stride_3_cycle_stride_r;
assign cfg_ld_dma_header.stride_3 = glb_pio_l2h_ld_dma_header_0_stride_3_stride_r;
assign cfg_ld_dma_header.range_3 = glb_pio_l2h_ld_dma_header_0_range_3_range_r;
assign cfg_ld_dma_header.cycle_stride_4 = glb_pio_l2h_ld_dma_header_0_cycle_stride_4_cycle_stride_r;
assign cfg_ld_dma_header.stride_4 = glb_pio_l2h_ld_dma_header_0_stride_4_stride_r;
assign cfg_ld_dma_header.range_4 = glb_pio_l2h_ld_dma_header_0_range_4_range_r;
assign cfg_ld_dma_header.cycle_stride_5 = glb_pio_l2h_ld_dma_header_0_cycle_stride_5_cycle_stride_r;
assign cfg_ld_dma_header.stride_5 = glb_pio_l2h_ld_dma_header_0_stride_5_stride_r;
assign cfg_ld_dma_header.range_5 = glb_pio_l2h_ld_dma_header_0_range_5_range_r;
assign cfg_ld_dma_header.cycle_stride_6 = glb_pio_l2h_ld_dma_header_0_cycle_stride_6_cycle_stride_r;
assign cfg_ld_dma_header.stride_6 = glb_pio_l2h_ld_dma_header_0_stride_6_stride_r;
assign cfg_ld_dma_header.range_6 = glb_pio_l2h_ld_dma_header_0_range_6_range_r;
assign cfg_ld_dma_header.cycle_stride_7 = glb_pio_l2h_ld_dma_header_0_cycle_stride_7_cycle_stride_r;
assign cfg_ld_dma_header.stride_7 = glb_pio_l2h_ld_dma_header_0_stride_7_stride_r;
assign cfg_ld_dma_header.range_7 = glb_pio_l2h_ld_dma_header_0_range_7_range_r;
assign cfg_pcfg_dma_ctrl.mode = glb_pio_l2h_pcfg_dma_ctrl_mode_r;
assign cfg_pcfg_dma_ctrl.relocation_value = glb_pio_l2h_pcfg_dma_ctrl_relocation_value_r;
assign cfg_pcfg_dma_ctrl.relocation_is_msb = glb_pio_l2h_pcfg_dma_ctrl_relocation_is_msb_r;
assign cfg_pcfg_dma_header.start_addr = glb_pio_l2h_pcfg_dma_header_start_addr_start_addr_r;
assign cfg_pcfg_dma_header.num_cfg = glb_pio_l2h_pcfg_dma_header_num_cfg_num_cfg_r;
assign cfg_pcfg_broadcast_mux.west = glb_pio_l2h_pcfg_broadcast_mux_west_r;
assign cfg_pcfg_broadcast_mux.east = glb_pio_l2h_pcfg_broadcast_mux_east_r;
assign cfg_pcfg_broadcast_mux.south = glb_pio_l2h_pcfg_broadcast_mux_south_r;
assign glb_pio_h2d_pio_dec_address = glb_cfg_ctrl_h2d_pio_dec_address[5:0];
glb_pio glb_pio (
  .clk(gclk),
  .h2d_pio_dec_address(glb_pio_h2d_pio_dec_address),
  .h2d_pio_dec_read(glb_pio_h2d_pio_dec_read),
  .h2d_pio_dec_write(glb_pio_h2d_pio_dec_write),
  .h2d_pio_dec_write_data(glb_pio_h2d_pio_dec_write_data),
  .reset(reset),
  .d2h_dec_pio_ack(glb_pio_d2h_dec_pio_ack),
  .d2h_dec_pio_nack(glb_pio_d2h_dec_pio_nack),
  .d2h_dec_pio_read_data(glb_pio_d2h_dec_pio_read_data),
  .l2h_data_network_ctrl_connected_r(glb_pio_l2h_data_network_ctrl_connected_r),
  .l2h_data_network_latency_value_r(glb_pio_l2h_data_network_latency_value_r),
  .l2h_ld_dma_ctrl_data_mux_r(glb_pio_l2h_ld_dma_ctrl_data_mux_r),
  .l2h_ld_dma_ctrl_mode_r(glb_pio_l2h_ld_dma_ctrl_mode_r),
  .l2h_ld_dma_ctrl_num_repeat_r(glb_pio_l2h_ld_dma_ctrl_num_repeat_r),
  .l2h_ld_dma_ctrl_use_flush_r(glb_pio_l2h_ld_dma_ctrl_use_flush_r),
  .l2h_ld_dma_ctrl_use_valid_r(glb_pio_l2h_ld_dma_ctrl_use_valid_r),
  .l2h_ld_dma_header_0_cycle_start_addr_cycle_start_addr_r(glb_pio_l2h_ld_dma_header_0_cycle_start_addr_cycle_start_addr_r),
  .l2h_ld_dma_header_0_cycle_stride_0_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_0_cycle_stride_r),
  .l2h_ld_dma_header_0_cycle_stride_1_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_1_cycle_stride_r),
  .l2h_ld_dma_header_0_cycle_stride_2_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_2_cycle_stride_r),
  .l2h_ld_dma_header_0_cycle_stride_3_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_3_cycle_stride_r),
  .l2h_ld_dma_header_0_cycle_stride_4_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_4_cycle_stride_r),
  .l2h_ld_dma_header_0_cycle_stride_5_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_5_cycle_stride_r),
  .l2h_ld_dma_header_0_cycle_stride_6_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_6_cycle_stride_r),
  .l2h_ld_dma_header_0_cycle_stride_7_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_7_cycle_stride_r),
  .l2h_ld_dma_header_0_dim_dim_r(glb_pio_l2h_ld_dma_header_0_dim_dim_r),
  .l2h_ld_dma_header_0_range_0_range_r(glb_pio_l2h_ld_dma_header_0_range_0_range_r),
  .l2h_ld_dma_header_0_range_1_range_r(glb_pio_l2h_ld_dma_header_0_range_1_range_r),
  .l2h_ld_dma_header_0_range_2_range_r(glb_pio_l2h_ld_dma_header_0_range_2_range_r),
  .l2h_ld_dma_header_0_range_3_range_r(glb_pio_l2h_ld_dma_header_0_range_3_range_r),
  .l2h_ld_dma_header_0_range_4_range_r(glb_pio_l2h_ld_dma_header_0_range_4_range_r),
  .l2h_ld_dma_header_0_range_5_range_r(glb_pio_l2h_ld_dma_header_0_range_5_range_r),
  .l2h_ld_dma_header_0_range_6_range_r(glb_pio_l2h_ld_dma_header_0_range_6_range_r),
  .l2h_ld_dma_header_0_range_7_range_r(glb_pio_l2h_ld_dma_header_0_range_7_range_r),
  .l2h_ld_dma_header_0_start_addr_start_addr_r(glb_pio_l2h_ld_dma_header_0_start_addr_start_addr_r),
  .l2h_ld_dma_header_0_stride_0_stride_r(glb_pio_l2h_ld_dma_header_0_stride_0_stride_r),
  .l2h_ld_dma_header_0_stride_1_stride_r(glb_pio_l2h_ld_dma_header_0_stride_1_stride_r),
  .l2h_ld_dma_header_0_stride_2_stride_r(glb_pio_l2h_ld_dma_header_0_stride_2_stride_r),
  .l2h_ld_dma_header_0_stride_3_stride_r(glb_pio_l2h_ld_dma_header_0_stride_3_stride_r),
  .l2h_ld_dma_header_0_stride_4_stride_r(glb_pio_l2h_ld_dma_header_0_stride_4_stride_r),
  .l2h_ld_dma_header_0_stride_5_stride_r(glb_pio_l2h_ld_dma_header_0_stride_5_stride_r),
  .l2h_ld_dma_header_0_stride_6_stride_r(glb_pio_l2h_ld_dma_header_0_stride_6_stride_r),
  .l2h_ld_dma_header_0_stride_7_stride_r(glb_pio_l2h_ld_dma_header_0_stride_7_stride_r),
  .l2h_pcfg_broadcast_mux_east_r(glb_pio_l2h_pcfg_broadcast_mux_east_r),
  .l2h_pcfg_broadcast_mux_south_r(glb_pio_l2h_pcfg_broadcast_mux_south_r),
  .l2h_pcfg_broadcast_mux_west_r(glb_pio_l2h_pcfg_broadcast_mux_west_r),
  .l2h_pcfg_dma_ctrl_mode_r(glb_pio_l2h_pcfg_dma_ctrl_mode_r),
  .l2h_pcfg_dma_ctrl_relocation_is_msb_r(glb_pio_l2h_pcfg_dma_ctrl_relocation_is_msb_r),
  .l2h_pcfg_dma_ctrl_relocation_value_r(glb_pio_l2h_pcfg_dma_ctrl_relocation_value_r),
  .l2h_pcfg_dma_header_num_cfg_num_cfg_r(glb_pio_l2h_pcfg_dma_header_num_cfg_num_cfg_r),
  .l2h_pcfg_dma_header_start_addr_start_addr_r(glb_pio_l2h_pcfg_dma_header_start_addr_start_addr_r),
  .l2h_pcfg_network_ctrl_connected_r(glb_pio_l2h_pcfg_network_ctrl_connected_r),
  .l2h_pcfg_network_latency_value_r(glb_pio_l2h_pcfg_network_latency_value_r),
  .l2h_st_dma_ctrl_data_mux_r(glb_pio_l2h_st_dma_ctrl_data_mux_r),
  .l2h_st_dma_ctrl_mode_r(glb_pio_l2h_st_dma_ctrl_mode_r),
  .l2h_st_dma_ctrl_num_repeat_r(glb_pio_l2h_st_dma_ctrl_num_repeat_r),
  .l2h_st_dma_ctrl_use_valid_r(glb_pio_l2h_st_dma_ctrl_use_valid_r),
  .l2h_st_dma_header_0_cycle_start_addr_cycle_start_addr_r(glb_pio_l2h_st_dma_header_0_cycle_start_addr_cycle_start_addr_r),
  .l2h_st_dma_header_0_cycle_stride_0_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_0_cycle_stride_r),
  .l2h_st_dma_header_0_cycle_stride_1_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_1_cycle_stride_r),
  .l2h_st_dma_header_0_cycle_stride_2_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_2_cycle_stride_r),
  .l2h_st_dma_header_0_cycle_stride_3_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_3_cycle_stride_r),
  .l2h_st_dma_header_0_cycle_stride_4_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_4_cycle_stride_r),
  .l2h_st_dma_header_0_cycle_stride_5_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_5_cycle_stride_r),
  .l2h_st_dma_header_0_cycle_stride_6_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_6_cycle_stride_r),
  .l2h_st_dma_header_0_cycle_stride_7_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_7_cycle_stride_r),
  .l2h_st_dma_header_0_dim_dim_r(glb_pio_l2h_st_dma_header_0_dim_dim_r),
  .l2h_st_dma_header_0_range_0_range_r(glb_pio_l2h_st_dma_header_0_range_0_range_r),
  .l2h_st_dma_header_0_range_1_range_r(glb_pio_l2h_st_dma_header_0_range_1_range_r),
  .l2h_st_dma_header_0_range_2_range_r(glb_pio_l2h_st_dma_header_0_range_2_range_r),
  .l2h_st_dma_header_0_range_3_range_r(glb_pio_l2h_st_dma_header_0_range_3_range_r),
  .l2h_st_dma_header_0_range_4_range_r(glb_pio_l2h_st_dma_header_0_range_4_range_r),
  .l2h_st_dma_header_0_range_5_range_r(glb_pio_l2h_st_dma_header_0_range_5_range_r),
  .l2h_st_dma_header_0_range_6_range_r(glb_pio_l2h_st_dma_header_0_range_6_range_r),
  .l2h_st_dma_header_0_range_7_range_r(glb_pio_l2h_st_dma_header_0_range_7_range_r),
  .l2h_st_dma_header_0_start_addr_start_addr_r(glb_pio_l2h_st_dma_header_0_start_addr_start_addr_r),
  .l2h_st_dma_header_0_stride_0_stride_r(glb_pio_l2h_st_dma_header_0_stride_0_stride_r),
  .l2h_st_dma_header_0_stride_1_stride_r(glb_pio_l2h_st_dma_header_0_stride_1_stride_r),
  .l2h_st_dma_header_0_stride_2_stride_r(glb_pio_l2h_st_dma_header_0_stride_2_stride_r),
  .l2h_st_dma_header_0_stride_3_stride_r(glb_pio_l2h_st_dma_header_0_stride_3_stride_r),
  .l2h_st_dma_header_0_stride_4_stride_r(glb_pio_l2h_st_dma_header_0_stride_4_stride_r),
  .l2h_st_dma_header_0_stride_5_stride_r(glb_pio_l2h_st_dma_header_0_stride_5_stride_r),
  .l2h_st_dma_header_0_stride_6_stride_r(glb_pio_l2h_st_dma_header_0_stride_6_stride_r),
  .l2h_st_dma_header_0_stride_7_stride_r(glb_pio_l2h_st_dma_header_0_stride_7_stride_r)
);

glb_cfg_ctrl glb_cfg_ctrl (
  .d2h_dec_pio_ack(glb_pio_d2h_dec_pio_ack),
  .d2h_dec_pio_nack(glb_pio_d2h_dec_pio_nack),
  .d2h_dec_pio_read_data(glb_pio_d2h_dec_pio_read_data),
  .gclk(gclk),
  .glb_tile_id(glb_tile_id),
  .mclk(mclk),
  .if_cfg_wst_s(if_cfg_wst_s),
  .if_cfg_est_m(if_cfg_est_m),
  .reset(reset),
  .h2d_pio_dec_address(glb_cfg_ctrl_h2d_pio_dec_address),
  .h2d_pio_dec_read(glb_pio_h2d_pio_dec_read),
  .h2d_pio_dec_write(glb_pio_h2d_pio_dec_write),
  .h2d_pio_dec_write_data(glb_pio_h2d_pio_dec_write_data)
);

endmodule   // glb_cfg

module glb_cfg_ctrl (
  glb_tile_ifc_A_12_D_32.master if_cfg_est_m,
  glb_tile_ifc_A_12_D_32.slave if_cfg_wst_s,
  input logic d2h_dec_pio_ack,
  input logic d2h_dec_pio_nack,
  input logic [31:0] d2h_dec_pio_read_data,
  input logic gclk,
  input logic glb_tile_id,
  input logic mclk,
  input logic reset,
  output logic [8:0] h2d_pio_dec_address,
  output logic h2d_pio_dec_read,
  output logic h2d_pio_dec_write,
  output logic [31:0] h2d_pio_dec_write_data
);

logic [8:0] addr_internal;
logic if_cfg_est_m_rd_clk_en_sel;
logic if_cfg_est_m_rd_clk_en_sel_first_cycle;
logic if_cfg_est_m_rd_clk_en_sel_latch;
logic if_cfg_est_m_wr_clk_en_sel;
logic if_cfg_est_m_wr_clk_en_sel_first_cycle;
logic if_cfg_est_m_wr_clk_en_sel_latch;
logic if_cfg_wst_s_rd_clk_en_d;
logic if_cfg_wst_s_wr_clk_en_d;
logic [31:0] rd_data_internal;
logic rd_data_valid_internal;
logic rd_en_d1;
logic rd_en_d2;
logic rd_tile_id_match;
logic read_internal;
logic [31:0] wr_data_internal;
logic wr_tile_id_match;
logic write_internal;
always_comb begin
  wr_tile_id_match = glb_tile_id == if_cfg_wst_s.wr_addr[11];
  rd_tile_id_match = glb_tile_id == if_cfg_wst_s.rd_addr[11];
end
always_comb begin
  wr_data_internal = 32'h0;
  addr_internal = 9'h0;
  read_internal = 1'h0;
  write_internal = 1'h0;
  if (if_cfg_wst_s.rd_en && rd_tile_id_match) begin
    addr_internal = if_cfg_wst_s.rd_addr[10:2];
    read_internal = 1'h1;
  end
  if (if_cfg_wst_s.wr_en && wr_tile_id_match) begin
    addr_internal = if_cfg_wst_s.wr_addr[10:2];
    wr_data_internal = if_cfg_wst_s.wr_data;
    write_internal = 1'h1;
  end
end

always_ff @(posedge gclk, posedge reset) begin
  if (reset) begin
    if_cfg_est_m.wr_en <= 1'h0;
    if_cfg_est_m.wr_addr <= 12'h0;
    if_cfg_est_m.wr_data <= 32'h0;
  end
  else if (~(wr_tile_id_match && (if_cfg_wst_s.wr_en == 1'h1))) begin
    if_cfg_est_m.wr_en <= if_cfg_wst_s.wr_en;
    if_cfg_est_m.wr_addr <= if_cfg_wst_s.wr_addr;
    if_cfg_est_m.wr_data <= if_cfg_wst_s.wr_data;
  end
  else begin
    if_cfg_est_m.wr_en <= 1'h0;
    if_cfg_est_m.wr_addr <= 12'h0;
    if_cfg_est_m.wr_data <= 32'h0;
  end
end

always_ff @(posedge gclk, posedge reset) begin
  if (reset) begin
    if_cfg_est_m.rd_en <= 1'h0;
    if_cfg_est_m.rd_addr <= 12'h0;
  end
  else if (~(rd_tile_id_match && (if_cfg_wst_s.rd_en == 1'h1))) begin
    if_cfg_est_m.rd_en <= if_cfg_wst_s.rd_en;
    if_cfg_est_m.rd_addr <= if_cfg_wst_s.rd_addr;
  end
  else begin
    if_cfg_est_m.rd_en <= 1'h0;
    if_cfg_est_m.rd_addr <= 12'h0;
  end
end

always_ff @(posedge gclk, posedge reset) begin
  if (reset) begin
    if_cfg_wst_s.rd_data <= 32'h0;
    if_cfg_wst_s.rd_data_valid <= 1'h0;
  end
  else if (rd_data_valid_internal) begin
    if_cfg_wst_s.rd_data <= rd_data_internal;
    if_cfg_wst_s.rd_data_valid <= rd_data_valid_internal;
  end
  else begin
    if_cfg_wst_s.rd_data <= if_cfg_est_m.rd_data;
    if_cfg_wst_s.rd_data_valid <= if_cfg_est_m.rd_data_valid;
  end
end

always_ff @(posedge gclk, posedge reset) begin
  if (reset) begin
    rd_en_d1 <= 1'h0;
    rd_en_d2 <= 1'h0;
  end
  else begin
    rd_en_d1 <= read_internal;
    rd_en_d2 <= rd_en_d1;
  end
end

always_ff @(posedge gclk, posedge reset) begin
  if (reset) begin
    rd_data_valid_internal <= 1'h0;
    rd_data_internal <= 32'h0;
  end
  else if ((rd_en_d2 == 1'h1) & (d2h_dec_pio_ack | d2h_dec_pio_nack)) begin
    rd_data_valid_internal <= 1'h1;
    rd_data_internal <= d2h_dec_pio_read_data;
  end
  else begin
    rd_data_valid_internal <= 1'h0;
    rd_data_internal <= 32'h0;
  end
end

always_ff @(posedge mclk, posedge reset) begin
  if (reset) begin
    if_cfg_wst_s_wr_clk_en_d <= 1'h0;
    if_cfg_wst_s_rd_clk_en_d <= 1'h0;
  end
  else begin
    if_cfg_wst_s_wr_clk_en_d <= if_cfg_wst_s.wr_clk_en;
    if_cfg_wst_s_rd_clk_en_d <= if_cfg_wst_s.rd_clk_en;
  end
end
always_comb begin
  if_cfg_est_m_wr_clk_en_sel_first_cycle = if_cfg_wst_s.wr_en & (~wr_tile_id_match);
  if_cfg_est_m_rd_clk_en_sel_first_cycle = if_cfg_wst_s.rd_en & (~rd_tile_id_match);
end

always_ff @(posedge mclk, posedge reset) begin
  if (reset) begin
    if_cfg_est_m_wr_clk_en_sel_latch <= 1'h0;
  end
  else if (if_cfg_wst_s.wr_en == 1'h1) begin
    if (wr_tile_id_match) begin
      if_cfg_est_m_wr_clk_en_sel_latch <= 1'h0;
    end
    else if_cfg_est_m_wr_clk_en_sel_latch <= 1'h1;
  end
  else if (if_cfg_wst_s.wr_clk_en == 1'h0) begin
    if_cfg_est_m_wr_clk_en_sel_latch <= 1'h0;
  end
end

always_ff @(posedge mclk, posedge reset) begin
  if (reset) begin
    if_cfg_est_m_rd_clk_en_sel_latch <= 1'h0;
  end
  else if (if_cfg_wst_s.rd_en == 1'h1) begin
    if (rd_tile_id_match) begin
      if_cfg_est_m_rd_clk_en_sel_latch <= 1'h0;
    end
    else if_cfg_est_m_rd_clk_en_sel_latch <= 1'h1;
  end
  else if (if_cfg_wst_s.rd_clk_en == 1'h0) begin
    if_cfg_est_m_rd_clk_en_sel_latch <= 1'h0;
  end
end
always_comb begin
  if_cfg_est_m_wr_clk_en_sel = if_cfg_est_m_wr_clk_en_sel_first_cycle | if_cfg_est_m_wr_clk_en_sel_latch;
  if_cfg_est_m_rd_clk_en_sel = if_cfg_est_m_rd_clk_en_sel_first_cycle | if_cfg_est_m_rd_clk_en_sel_latch;
end
always_comb begin
  if (if_cfg_est_m_wr_clk_en_sel) begin
    if_cfg_est_m.wr_clk_en = if_cfg_wst_s_wr_clk_en_d;
  end
  else if_cfg_est_m.wr_clk_en = 1'h0;
end
always_comb begin
  if (if_cfg_est_m_rd_clk_en_sel) begin
    if_cfg_est_m.rd_clk_en = if_cfg_wst_s_rd_clk_en_d;
  end
  else if_cfg_est_m.rd_clk_en = 1'h0;
end
assign h2d_pio_dec_write_data = wr_data_internal;
assign h2d_pio_dec_address = addr_internal;
assign h2d_pio_dec_read = read_internal;
assign h2d_pio_dec_write = write_internal;
endmodule   // glb_cfg_ctrl

module glb_clk_en_gen (
  input logic clk,
  input logic enable,
  input logic reset,
  output logic clk_en
);

logic [1:0] clk_en_cnt;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    clk_en_cnt <= 2'h0;
  end
  else if (enable) begin
    clk_en_cnt <= 2'h3;
  end
  else if (clk_en_cnt > 2'h0) begin
    clk_en_cnt <= clk_en_cnt - 2'h1;
  end
end
assign clk_en = enable | (clk_en_cnt > 2'h0);
endmodule   // glb_clk_en_gen

module glb_clk_en_gen_unq0 (
  input logic clk,
  input logic enable,
  input logic reset,
  output logic clk_en
);

logic [2:0] clk_en_cnt;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    clk_en_cnt <= 3'h0;
  end
  else if (enable) begin
    clk_en_cnt <= 3'h5;
  end
  else if (clk_en_cnt > 3'h0) begin
    clk_en_cnt <= clk_en_cnt - 3'h1;
  end
end
assign clk_en = enable | (clk_en_cnt > 3'h0);
endmodule   // glb_clk_en_gen_unq0

module glb_clk_en_gen_unq1 (
  input logic clk,
  input logic enable,
  input logic reset,
  output logic clk_en
);

logic [2:0] clk_en_cnt;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    clk_en_cnt <= 3'h0;
  end
  else if (enable) begin
    clk_en_cnt <= 3'h4;
  end
  else if (clk_en_cnt > 3'h0) begin
    clk_en_cnt <= clk_en_cnt - 3'h1;
  end
end
assign clk_en = enable | (clk_en_cnt > 3'h0);
endmodule   // glb_clk_en_gen_unq1

module glb_clk_en_gen_unq2 (
  input logic clk,
  input logic enable,
  input logic reset,
  output logic clk_en
);

logic [3:0] clk_en_cnt;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    clk_en_cnt <= 4'h0;
  end
  else if (enable) begin
    clk_en_cnt <= 4'hA;
  end
  else if (clk_en_cnt > 4'h0) begin
    clk_en_cnt <= clk_en_cnt - 4'h1;
  end
end
assign clk_en = enable | (clk_en_cnt > 4'h0);
endmodule   // glb_clk_en_gen_unq2

module glb_crossbar_I_2_O_1_W_1 (
  input logic [1:0] in_,
  input logic sel_,
  output logic out_
);

always_comb begin
  out_ = in_[sel_];
end
endmodule   // glb_crossbar_I_2_O_1_W_1

module glb_load_dma (
  input logic [1:0] cfg_data_network_g2f_mux,
  input logic [5:0] cfg_data_network_latency,
  input logic [1:0] cfg_ld_dma_ctrl_mode,
  input logic cfg_ld_dma_ctrl_use_flush,
  input logic cfg_ld_dma_ctrl_use_valid,
  input dma_header_t cfg_ld_dma_header,
  input logic cfg_ld_dma_num_repeat,
  input logic cfg_tile_connected_next,
  input logic cfg_tile_connected_prev,
  input logic clk,
  input logic glb_tile_id,
  input logic ld_dma_start_pulse,
  input rdrs_packet_t rdrs_packet_bank2dma,
  input rdrs_packet_t rdrs_packet_ring2dma,
  input logic reset,
  output logic clk_en_dma2bank,
  output logic data_flush,
  output logic [1:0] [15:0] data_g2f,
  output logic [1:0] data_valid_g2f,
  output logic ld_dma_done_interrupt,
  output rdrq_packet_t rdrq_packet_dma2bank,
  output rdrq_packet_t rdrq_packet_dma2ring
);

logic [18:0] bank_rdrq_rd_addr;
logic bank_rdrq_rd_en;
logic [63:0] bank_rdrs_data_cache_r;
dma_header_t current_dma_header;
logic [15:0] cycle_count;
logic [15:0] cycle_current_addr;
logic [7:0][15:0] cycle_stride_addr_gen_strides;
logic cycle_valid;
logic [19:0] data_current_addr;
logic data_flush_w;
logic [1:0][15:0] data_g2f_w;
logic [19:0] data_stride_addr_gen_start_addr;
logic [7:0][19:0] data_stride_addr_gen_strides;
logic [1:0] data_valid_g2f_w;
logic dma2bank_clk_en;
logic is_cached;
logic is_first;
logic [18:0] last_strm_rd_addr_r;
logic ld_dma_done_pulse;
logic ld_dma_done_pulse_d_arr [10:0];
logic ld_dma_done_pulse_last;
logic ld_dma_done_pulse_w;
logic ld_dma_start_pulse_next;
logic ld_dma_start_pulse_r;
logic loop_done;
logic [7:0][31:0] loop_iter_ranges;
logic [2:0] loop_mux_sel;
rdrq_packet_t rdrq_packet_dma2bank_w;
rdrq_packet_t rdrq_packet_dma2ring_w;
rdrs_packet_t rdrs_packet;
logic repeat_cnt;
logic [15:0] strm_data;
logic [15:0] strm_data_muxed;
logic [1:0] strm_data_sel_arr [9:0];
logic [1:0] strm_data_sel_w;
logic strm_data_start_pulse;
logic strm_data_start_pulse_d_arr [9:0];
logic strm_data_valid;
logic strm_data_valid_muxed;
logic [18:0] strm_rd_addr_w;
logic strm_rd_en_d_arr [9:0];
logic strm_rd_en_w;
logic strm_run;
assign current_dma_header = cfg_ld_dma_header;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    repeat_cnt <= 1'h0;
  end
  else if (cfg_ld_dma_ctrl_mode == 2'h2) begin
    if (ld_dma_done_pulse) begin
      if ((repeat_cnt + 1'h1) < cfg_ld_dma_num_repeat) begin
        repeat_cnt <= repeat_cnt + 1'h1;
      end
    end
  end
  else if (cfg_ld_dma_ctrl_mode == 2'h3) begin
    if (ld_dma_done_pulse) begin
      if (((repeat_cnt + 1'h1) < cfg_ld_dma_num_repeat) & ((repeat_cnt + 1'h1) < 1'h1)) begin
        repeat_cnt <= repeat_cnt + 1'h1;
      end
    end
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    cycle_count <= 16'h0;
  end
  else if (ld_dma_start_pulse_r) begin
    cycle_count <= 16'h0;
  end
  else if (loop_done) begin
    cycle_count <= 16'h0;
  end
  else if (strm_run) begin
    cycle_count <= cycle_count + 16'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    is_first <= 1'h0;
  end
  else if (ld_dma_start_pulse_r) begin
    is_first <= 1'h1;
  end
  else if (bank_rdrq_rd_en) begin
    is_first <= 1'h0;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    strm_run <= 1'h0;
  end
  else if (ld_dma_start_pulse_r) begin
    strm_run <= 1'h1;
  end
  else if (loop_done) begin
    strm_run <= 1'h0;
  end
end
always_comb begin
  if (cfg_ld_dma_ctrl_use_flush == 1'h1) begin
    strm_data_start_pulse = strm_data_start_pulse_d_arr[(4'(cfg_data_network_latency) + 4'h3) - 4'h1];
  end
  else strm_data_start_pulse = strm_data_start_pulse_d_arr[4'(cfg_data_network_latency) + 4'h3];
end
assign strm_data_valid = strm_rd_en_d_arr[4'(cfg_data_network_latency) + 4'h3];
assign strm_data_sel_w = strm_rd_addr_w[2:1];
always_comb begin
  if (cfg_ld_dma_ctrl_mode == 2'h0) begin
    ld_dma_start_pulse_next = 1'h0;
  end
  else if (cfg_ld_dma_ctrl_mode == 2'h1) begin
    ld_dma_start_pulse_next = (~strm_run) & ld_dma_start_pulse;
  end
  else if ((cfg_ld_dma_ctrl_mode == 2'h2) | (cfg_ld_dma_ctrl_mode == 2'h3)) begin
    ld_dma_start_pulse_next = ((~strm_run) & ld_dma_start_pulse) | (ld_dma_done_pulse & ((repeat_cnt + 1'h1) <
        cfg_ld_dma_num_repeat));
  end
  else ld_dma_start_pulse_next = 1'h0;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    ld_dma_start_pulse_r <= 1'h0;
  end
  else if (ld_dma_start_pulse_r) begin
    ld_dma_start_pulse_r <= 1'h0;
  end
  else ld_dma_start_pulse_r <= ld_dma_start_pulse_next;
end
always_comb begin
  strm_data_muxed = strm_data;
  if (cfg_ld_dma_ctrl_use_valid) begin
    strm_data_valid_muxed = strm_data_valid;
  end
  else if (~cfg_ld_dma_ctrl_use_flush) begin
    strm_data_valid_muxed = strm_data_start_pulse;
  end
  else strm_data_valid_muxed = 1'h0;
end
always_comb begin
  if (cfg_data_network_g2f_mux[0] == 1'h1) begin
    data_g2f_w[0] = strm_data_muxed;
    data_valid_g2f_w[0] = strm_data_valid_muxed;
  end
  else begin
    data_g2f_w[0] = 16'h0;
    data_valid_g2f_w[0] = 1'h0;
  end
  if (cfg_data_network_g2f_mux[1] == 1'h1) begin
    data_g2f_w[1] = strm_data_muxed;
    data_valid_g2f_w[1] = strm_data_valid_muxed;
  end
  else begin
    data_g2f_w[1] = 16'h0;
    data_valid_g2f_w[1] = 1'h0;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    data_g2f <= 32'h0;
    data_valid_g2f <= 2'h0;
  end
  else begin
    data_g2f[0] <= data_g2f_w[0];
    data_g2f[1] <= data_g2f_w[1];
    data_valid_g2f <= data_valid_g2f_w;
  end
end
always_comb begin
  ld_dma_done_pulse_w = strm_run & loop_done;
end
always_comb begin
  strm_rd_en_w = cycle_valid;
  strm_rd_addr_w = 19'(data_current_addr);
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    last_strm_rd_addr_r <= 19'h0;
  end
  else if (strm_rd_en_w) begin
    last_strm_rd_addr_r <= strm_rd_addr_w;
  end
end
always_comb begin
  if (cfg_tile_connected_next | cfg_tile_connected_prev) begin
    rdrq_packet_dma2bank_w = 20'h0;
    rdrq_packet_dma2ring_w.rd_en = bank_rdrq_rd_en;
    rdrq_packet_dma2ring_w.rd_addr = bank_rdrq_rd_addr;
  end
  else begin
    rdrq_packet_dma2bank_w.rd_en = bank_rdrq_rd_en;
    rdrq_packet_dma2bank_w.rd_addr = bank_rdrq_rd_addr;
    rdrq_packet_dma2ring_w = 20'h0;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    rdrq_packet_dma2bank <= 20'h0;
    rdrq_packet_dma2ring <= 20'h0;
  end
  else begin
    rdrq_packet_dma2bank <= rdrq_packet_dma2bank_w;
    rdrq_packet_dma2ring <= rdrq_packet_dma2ring_w;
  end
end
always_comb begin
  is_cached = strm_rd_addr_w[18:3] == last_strm_rd_addr_r[18:3];
  bank_rdrq_rd_en = strm_rd_en_w & (is_first | (~is_cached));
  bank_rdrq_rd_addr = strm_rd_addr_w;
end
always_comb begin
  if (cfg_tile_connected_next | cfg_tile_connected_prev) begin
    rdrs_packet = rdrs_packet_ring2dma;
  end
  else rdrs_packet = rdrs_packet_bank2dma;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    bank_rdrs_data_cache_r <= 64'h0;
  end
  else if (rdrs_packet.rd_data_valid) begin
    bank_rdrs_data_cache_r <= rdrs_packet.rd_data;
  end
end
always_comb begin
  unique case (strm_data_sel_arr[4'(cfg_data_network_latency) + 4'h3])
    2'h0: strm_data = bank_rdrs_data_cache_r[15:0];
    2'h1: strm_data = bank_rdrs_data_cache_r[31:16];
    2'h2: strm_data = bank_rdrs_data_cache_r[47:32];
    2'h3: strm_data = bank_rdrs_data_cache_r[63:48];
    default: strm_data = bank_rdrs_data_cache_r[15:0];
  endcase
end
assign ld_dma_done_pulse = ld_dma_done_pulse_d_arr[4'(cfg_data_network_latency) + 4'h3 + 4'h1];

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    ld_dma_done_interrupt <= 1'h0;
  end
  else if (ld_dma_done_pulse) begin
    ld_dma_done_interrupt <= 1'h1;
  end
  else if (ld_dma_done_pulse_last) begin
    ld_dma_done_interrupt <= 1'h0;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    data_flush <= 1'h0;
  end
  else data_flush <= data_flush_w;
end
always_comb begin
  if (cfg_ld_dma_ctrl_use_flush) begin
    data_flush_w = strm_data_start_pulse;
  end
  else data_flush_w = 1'h0;
end
assign clk_en_dma2bank = dma2bank_clk_en;
assign loop_iter_ranges[0] = current_dma_header.range_0;
assign loop_iter_ranges[1] = current_dma_header.range_1;
assign loop_iter_ranges[2] = current_dma_header.range_2;
assign loop_iter_ranges[3] = current_dma_header.range_3;
assign loop_iter_ranges[4] = current_dma_header.range_4;
assign loop_iter_ranges[5] = current_dma_header.range_5;
assign loop_iter_ranges[6] = current_dma_header.range_6;
assign loop_iter_ranges[7] = current_dma_header.range_7;
assign cycle_stride_addr_gen_strides[0] = current_dma_header.cycle_stride_0;
assign cycle_stride_addr_gen_strides[1] = current_dma_header.cycle_stride_1;
assign cycle_stride_addr_gen_strides[2] = current_dma_header.cycle_stride_2;
assign cycle_stride_addr_gen_strides[3] = current_dma_header.cycle_stride_3;
assign cycle_stride_addr_gen_strides[4] = current_dma_header.cycle_stride_4;
assign cycle_stride_addr_gen_strides[5] = current_dma_header.cycle_stride_5;
assign cycle_stride_addr_gen_strides[6] = current_dma_header.cycle_stride_6;
assign cycle_stride_addr_gen_strides[7] = current_dma_header.cycle_stride_7;
assign data_stride_addr_gen_start_addr = 20'(current_dma_header.start_addr);
assign data_stride_addr_gen_strides[0] = current_dma_header.stride_0;
assign data_stride_addr_gen_strides[1] = current_dma_header.stride_1;
assign data_stride_addr_gen_strides[2] = current_dma_header.stride_2;
assign data_stride_addr_gen_strides[3] = current_dma_header.stride_3;
assign data_stride_addr_gen_strides[4] = current_dma_header.stride_4;
assign data_stride_addr_gen_strides[5] = current_dma_header.stride_5;
assign data_stride_addr_gen_strides[6] = current_dma_header.stride_6;
assign data_stride_addr_gen_strides[7] = current_dma_header.stride_7;
pipeline_w_1_d_10_array strm_dma_start_pulse_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(ld_dma_start_pulse_r),
  .reset(reset),
  .out_(strm_data_start_pulse_d_arr)
);

pipeline_w_1_d_10_array strm_rd_en_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(strm_rd_en_w),
  .reset(reset),
  .out_(strm_rd_en_d_arr)
);

pipeline_w_2_d_10_array strm_data_sel_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(strm_data_sel_w),
  .reset(reset),
  .out_(strm_data_sel_arr)
);

pipeline_w_1_d_11_array ld_dma_done_pulse_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(ld_dma_done_pulse_w),
  .reset(reset),
  .out_(ld_dma_done_pulse_d_arr)
);

pipeline_w_1_d_5 ld_dma_interrupt_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(ld_dma_done_pulse),
  .reset(reset),
  .out_(ld_dma_done_pulse_last)
);

glb_clk_en_gen_unq0 dma2bank_clk_en_gen (
  .clk(clk),
  .enable(rdrq_packet_dma2bank_w.rd_en),
  .reset(reset),
  .clk_en(dma2bank_clk_en)
);

glb_loop_iter loop_iter (
  .clk(clk),
  .clk_en(1'h1),
  .dim(current_dma_header.dim),
  .ranges(loop_iter_ranges),
  .reset(reset),
  .step(cycle_valid),
  .mux_sel_out(loop_mux_sel),
  .restart(loop_done)
);

glb_sched_gen cycle_stride_sched_gen (
  .clk(clk),
  .clk_en(1'h1),
  .current_addr(cycle_current_addr),
  .cycle_count(cycle_count),
  .finished(loop_done),
  .reset(reset),
  .restart(ld_dma_start_pulse_r),
  .valid_output(cycle_valid)
);

glb_addr_gen #(
  .addr_width(32'h10))
cycle_stride_addr_gen (
  .clk(clk),
  .clk_en(1'h1),
  .mux_sel(loop_mux_sel),
  .reset(reset),
  .restart(ld_dma_start_pulse_r),
  .start_addr(current_dma_header.cycle_start_addr),
  .step(cycle_valid),
  .strides(cycle_stride_addr_gen_strides),
  .addr_out(cycle_current_addr)
);

glb_addr_gen #(
  .addr_width(32'h14))
data_stride_addr_gen (
  .clk(clk),
  .clk_en(1'h1),
  .mux_sel(loop_mux_sel),
  .reset(reset),
  .restart(ld_dma_start_pulse_r),
  .start_addr(data_stride_addr_gen_start_addr),
  .step(cycle_valid),
  .strides(data_stride_addr_gen_strides),
  .addr_out(data_current_addr)
);

endmodule   // glb_load_dma

module glb_loop_iter (
  input logic clk,
  input logic clk_en,
  input logic [3:0] dim,
  input logic [7:0] [31:0] ranges,
  input logic reset,
  input logic step,
  output logic [2:0] mux_sel_out,
  output logic restart
);

logic [7:0] clear;
logic [7:0][31:0] dim_counter;
logic [7:0] inc;
logic is_maxed;
logic [7:0] max_value;
logic [2:0] mux_sel;
logic not_done;
assign mux_sel_out = mux_sel;
assign is_maxed = (dim_counter[mux_sel] == ranges[mux_sel]) & inc[mux_sel];
always_comb begin
  mux_sel = 3'h0;
  not_done = 1'h0;
  for (int unsigned i = 0; i < 8; i += 1) begin
      if (~not_done) begin
        if ((~max_value[3'(i)]) & (4'(i) < dim)) begin
          mux_sel = 3'(i);
          not_done = 1'h1;
        end
      end
    end
end
always_comb begin
  clear[0] = 1'h0;
  if (((mux_sel > 3'h0) | (~not_done)) & step) begin
    clear[0] = 1'h1;
  end
end
always_comb begin
  inc[0] = 1'h0;
  if ((5'h0 == 5'h0) & step & (dim > 4'h0)) begin
    inc[0] = 1'h1;
  end
  else if ((mux_sel == 3'h0) & step & (dim > 4'h0)) begin
    inc[0] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[0] <= 32'h0;
  end
  else if (clear[0]) begin
    dim_counter[0] <= 32'h0;
  end
  else if (inc[0]) begin
    dim_counter[0] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[0] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[0]) begin
      max_value[0] <= 1'h0;
    end
    else if (inc[0]) begin
      max_value[0] <= is_maxed;
    end
  end
end
always_comb begin
  clear[1] = 1'h0;
  if (((mux_sel > 3'h1) | (~not_done)) & step) begin
    clear[1] = 1'h1;
  end
end
always_comb begin
  inc[1] = 1'h0;
  if ((5'h1 == 5'h0) & step & (dim > 4'h1)) begin
    inc[1] = 1'h1;
  end
  else if ((mux_sel == 3'h1) & step & (dim > 4'h1)) begin
    inc[1] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[1] <= 32'h0;
  end
  else if (clear[1]) begin
    dim_counter[1] <= 32'h0;
  end
  else if (inc[1]) begin
    dim_counter[1] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[1] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[1]) begin
      max_value[1] <= 1'h0;
    end
    else if (inc[1]) begin
      max_value[1] <= is_maxed;
    end
  end
end
always_comb begin
  clear[2] = 1'h0;
  if (((mux_sel > 3'h2) | (~not_done)) & step) begin
    clear[2] = 1'h1;
  end
end
always_comb begin
  inc[2] = 1'h0;
  if ((5'h2 == 5'h0) & step & (dim > 4'h2)) begin
    inc[2] = 1'h1;
  end
  else if ((mux_sel == 3'h2) & step & (dim > 4'h2)) begin
    inc[2] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[2] <= 32'h0;
  end
  else if (clear[2]) begin
    dim_counter[2] <= 32'h0;
  end
  else if (inc[2]) begin
    dim_counter[2] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[2] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[2]) begin
      max_value[2] <= 1'h0;
    end
    else if (inc[2]) begin
      max_value[2] <= is_maxed;
    end
  end
end
always_comb begin
  clear[3] = 1'h0;
  if (((mux_sel > 3'h3) | (~not_done)) & step) begin
    clear[3] = 1'h1;
  end
end
always_comb begin
  inc[3] = 1'h0;
  if ((5'h3 == 5'h0) & step & (dim > 4'h3)) begin
    inc[3] = 1'h1;
  end
  else if ((mux_sel == 3'h3) & step & (dim > 4'h3)) begin
    inc[3] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[3] <= 32'h0;
  end
  else if (clear[3]) begin
    dim_counter[3] <= 32'h0;
  end
  else if (inc[3]) begin
    dim_counter[3] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[3] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[3]) begin
      max_value[3] <= 1'h0;
    end
    else if (inc[3]) begin
      max_value[3] <= is_maxed;
    end
  end
end
always_comb begin
  clear[4] = 1'h0;
  if (((mux_sel > 3'h4) | (~not_done)) & step) begin
    clear[4] = 1'h1;
  end
end
always_comb begin
  inc[4] = 1'h0;
  if ((5'h4 == 5'h0) & step & (dim > 4'h4)) begin
    inc[4] = 1'h1;
  end
  else if ((mux_sel == 3'h4) & step & (dim > 4'h4)) begin
    inc[4] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[4] <= 32'h0;
  end
  else if (clear[4]) begin
    dim_counter[4] <= 32'h0;
  end
  else if (inc[4]) begin
    dim_counter[4] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[4] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[4]) begin
      max_value[4] <= 1'h0;
    end
    else if (inc[4]) begin
      max_value[4] <= is_maxed;
    end
  end
end
always_comb begin
  clear[5] = 1'h0;
  if (((mux_sel > 3'h5) | (~not_done)) & step) begin
    clear[5] = 1'h1;
  end
end
always_comb begin
  inc[5] = 1'h0;
  if ((5'h5 == 5'h0) & step & (dim > 4'h5)) begin
    inc[5] = 1'h1;
  end
  else if ((mux_sel == 3'h5) & step & (dim > 4'h5)) begin
    inc[5] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[5] <= 32'h0;
  end
  else if (clear[5]) begin
    dim_counter[5] <= 32'h0;
  end
  else if (inc[5]) begin
    dim_counter[5] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[5] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[5]) begin
      max_value[5] <= 1'h0;
    end
    else if (inc[5]) begin
      max_value[5] <= is_maxed;
    end
  end
end
always_comb begin
  clear[6] = 1'h0;
  if (((mux_sel > 3'h6) | (~not_done)) & step) begin
    clear[6] = 1'h1;
  end
end
always_comb begin
  inc[6] = 1'h0;
  if ((5'h6 == 5'h0) & step & (dim > 4'h6)) begin
    inc[6] = 1'h1;
  end
  else if ((mux_sel == 3'h6) & step & (dim > 4'h6)) begin
    inc[6] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[6] <= 32'h0;
  end
  else if (clear[6]) begin
    dim_counter[6] <= 32'h0;
  end
  else if (inc[6]) begin
    dim_counter[6] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[6] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[6]) begin
      max_value[6] <= 1'h0;
    end
    else if (inc[6]) begin
      max_value[6] <= is_maxed;
    end
  end
end
always_comb begin
  clear[7] = 1'h0;
  if (((mux_sel > 3'h7) | (~not_done)) & step) begin
    clear[7] = 1'h1;
  end
end
always_comb begin
  inc[7] = 1'h0;
  if ((5'h7 == 5'h0) & step & (dim > 4'h7)) begin
    inc[7] = 1'h1;
  end
  else if ((mux_sel == 3'h7) & step & (dim > 4'h7)) begin
    inc[7] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[7] <= 32'h0;
  end
  else if (clear[7]) begin
    dim_counter[7] <= 32'h0;
  end
  else if (inc[7]) begin
    dim_counter[7] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[7] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[7]) begin
      max_value[7] <= 1'h0;
    end
    else if (inc[7]) begin
      max_value[7] <= is_maxed;
    end
  end
end
assign restart = step & (~not_done);
endmodule   // glb_loop_iter

module glb_pcfg_broadcast (
  input pcfg_broadcast_mux_t cfg_pcfg_broadcast_mux,
  input cgra_cfg_t cgra_cfg_dma2mux,
  input logic [31:0] cgra_cfg_jtag_addr_bypass_wsti,
  input logic cgra_cfg_jtag_rd_en_bypass_wsti,
  input cgra_cfg_t cgra_cfg_jtag_wsti,
  input cgra_cfg_t cgra_cfg_pcfg_esti,
  input cgra_cfg_t cgra_cfg_pcfg_wsti,
  input logic clk,
  input logic reset,
  output cgra_cfg_t [1:0] cgra_cfg_g2f,
  output logic [31:0] cgra_cfg_jtag_addr_bypass_esto,
  output cgra_cfg_t cgra_cfg_jtag_esto,
  output logic cgra_cfg_jtag_rd_en_bypass_esto,
  output cgra_cfg_t cgra_cfg_pcfg_esto,
  output cgra_cfg_t cgra_cfg_pcfg_wsto
);

cgra_cfg_t [1:0] cgra_cfg_g2f_w;
cgra_cfg_t pcfg_east_muxed;
cgra_cfg_t pcfg_south_muxed;
cgra_cfg_t pcfg_west_muxed;
always_comb begin
  cgra_cfg_jtag_rd_en_bypass_esto = cgra_cfg_jtag_rd_en_bypass_wsti;
  cgra_cfg_jtag_addr_bypass_esto = cgra_cfg_jtag_addr_bypass_wsti;
end
always_comb begin
  if (cfg_pcfg_broadcast_mux.south == 2'h0) begin
    pcfg_south_muxed = 66'h0;
  end
  else if (cfg_pcfg_broadcast_mux.south == 2'h1) begin
    pcfg_south_muxed = cgra_cfg_dma2mux;
  end
  else if (cfg_pcfg_broadcast_mux.south == 2'h2) begin
    pcfg_south_muxed = cgra_cfg_pcfg_wsti;
  end
  else if (cfg_pcfg_broadcast_mux.south == 2'h3) begin
    pcfg_south_muxed = cgra_cfg_pcfg_esti;
  end
  else pcfg_south_muxed = 66'h0;
end
always_comb begin
  if (cfg_pcfg_broadcast_mux.west == 2'h0) begin
    pcfg_west_muxed = 66'h0;
  end
  else if (cfg_pcfg_broadcast_mux.west == 2'h1) begin
    pcfg_west_muxed = cgra_cfg_dma2mux;
  end
  else if (cfg_pcfg_broadcast_mux.west == 2'h2) begin
    pcfg_west_muxed = cgra_cfg_pcfg_esti;
  end
  else pcfg_west_muxed = 66'h0;
end
always_comb begin
  if (cfg_pcfg_broadcast_mux.east == 2'h0) begin
    pcfg_east_muxed = 66'h0;
  end
  else if (cfg_pcfg_broadcast_mux.east == 2'h1) begin
    pcfg_east_muxed = cgra_cfg_dma2mux;
  end
  else if (cfg_pcfg_broadcast_mux.east == 2'h2) begin
    pcfg_east_muxed = cgra_cfg_pcfg_wsti;
  end
  else pcfg_east_muxed = 66'h0;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    cgra_cfg_jtag_esto <= 66'h0;
  end
  else cgra_cfg_jtag_esto <= cgra_cfg_jtag_wsti;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    cgra_cfg_pcfg_esto <= 66'h0;
    cgra_cfg_pcfg_wsto <= 66'h0;
  end
  else begin
    cgra_cfg_pcfg_esto <= pcfg_east_muxed;
    cgra_cfg_pcfg_wsto <= pcfg_west_muxed;
  end
end
always_comb begin
  if (cgra_cfg_jtag_rd_en_bypass_esto) begin
    cgra_cfg_g2f_w[0].wr_en = 1'h0;
    cgra_cfg_g2f_w[0].rd_en = 1'h1;
    cgra_cfg_g2f_w[0].addr = cgra_cfg_jtag_addr_bypass_esto;
    cgra_cfg_g2f_w[0].data = 32'h0;
  end
  else cgra_cfg_g2f_w[0] = cgra_cfg_jtag_wsti | pcfg_south_muxed;
end
always_comb begin
  if (cgra_cfg_jtag_rd_en_bypass_esto) begin
    cgra_cfg_g2f_w[1].wr_en = 1'h0;
    cgra_cfg_g2f_w[1].rd_en = 1'h1;
    cgra_cfg_g2f_w[1].addr = cgra_cfg_jtag_addr_bypass_esto;
    cgra_cfg_g2f_w[1].data = 32'h0;
  end
  else cgra_cfg_g2f_w[1] = cgra_cfg_jtag_wsti | pcfg_south_muxed;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    for (int unsigned i = 0; i < 2; i += 1) begin
        cgra_cfg_g2f[1'(i)] <= 66'h0;
      end
  end
  else begin
    for (int unsigned i = 0; i < 2; i += 1) begin
        cgra_cfg_g2f[1'(i)] <= cgra_cfg_g2f_w[1'(i)];
      end
  end
end
endmodule   // glb_pcfg_broadcast

module glb_pcfg_dma (
  input logic cfg_pcfg_dma_ctrl_mode,
  input logic cfg_pcfg_dma_ctrl_relocation_is_msb,
  input logic [15:0] cfg_pcfg_dma_ctrl_relocation_value,
  input pcfg_dma_header_t cfg_pcfg_dma_header,
  input logic [5:0] cfg_pcfg_network_latency,
  input logic cfg_pcfg_tile_connected_next,
  input logic cfg_pcfg_tile_connected_prev,
  input logic clk,
  input logic glb_tile_id,
  input logic pcfg_dma_start_pulse,
  input rdrs_packet_t rdrs_packet_bank2dma,
  input rdrs_packet_t rdrs_packet_ring2dma,
  input logic reset,
  output cgra_cfg_t cgra_cfg_pcfg,
  output logic clk_en_dma2bank,
  output logic pcfg_dma_done_interrupt,
  output rdrq_packet_t rdrq_packet_dma2bank,
  output rdrq_packet_t rdrq_packet_dma2ring
);

logic [18:0] addr_next;
logic [18:0] addr_r;
logic dma2bank_clk_en;
logic done_pulse_d_arr [11:0];
logic done_pulse_r;
logic is_running_r;
logic [15:0] num_cfg_cnt_next;
logic [15:0] num_cfg_cnt_r;
logic pcfg_done_pulse;
logic pcfg_done_pulse_last;
rdrq_packet_t rdrq_packet_dma2bank_w;
rdrq_packet_t rdrq_packet_dma2ring_w;
logic [18:0] rdrq_packet_rd_addr_next;
logic rdrq_packet_rd_en_next;
rdrs_packet_t rdrs_packet;
logic [63:0] rdrs_packet_rd_data_r;
logic rdrs_packet_rd_data_valid_r;
logic start_pulse_r;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    start_pulse_r <= 1'h0;
  end
  else if ((cfg_pcfg_dma_ctrl_mode == 1'h1) & (~is_running_r) & pcfg_dma_start_pulse) begin
    start_pulse_r <= 1'h1;
  end
  else start_pulse_r <= 1'h0;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    done_pulse_r <= 1'h0;
  end
  else if (is_running_r & (num_cfg_cnt_r == 16'h0)) begin
    done_pulse_r <= 1'h1;
  end
  else done_pulse_r <= 1'h0;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    is_running_r <= 1'h0;
  end
  else if (start_pulse_r) begin
    is_running_r <= 1'h1;
  end
  else if ((is_running_r == 1'h1) & (num_cfg_cnt_r == 16'h0)) begin
    is_running_r <= 1'h0;
  end
end
always_comb begin
  if (start_pulse_r) begin
    num_cfg_cnt_next = cfg_pcfg_dma_header.num_cfg;
    addr_next = cfg_pcfg_dma_header.start_addr;
  end
  else if ((is_running_r == 1'h1) & (num_cfg_cnt_r > 16'h0)) begin
    num_cfg_cnt_next = num_cfg_cnt_r - 16'h1;
    addr_next = addr_r + 19'h8;
  end
  else begin
    num_cfg_cnt_next = 16'h0;
    addr_next = 19'h0;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    num_cfg_cnt_r <= 16'h0;
    addr_r <= 19'h0;
  end
  else begin
    num_cfg_cnt_r <= num_cfg_cnt_next;
    addr_r <= addr_next;
  end
end
always_comb begin
  if (is_running_r & (num_cfg_cnt_r > 16'h0)) begin
    rdrq_packet_rd_en_next = 1'h1;
    rdrq_packet_rd_addr_next = addr_r;
  end
  else begin
    rdrq_packet_rd_en_next = 1'h0;
    rdrq_packet_rd_addr_next = 19'h0;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    rdrq_packet_dma2ring <= 20'h0;
    rdrq_packet_dma2bank <= 20'h0;
  end
  else begin
    rdrq_packet_dma2ring <= rdrq_packet_dma2ring_w;
    rdrq_packet_dma2bank <= rdrq_packet_dma2bank_w;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    rdrs_packet_rd_data_r <= 64'h0;
    rdrs_packet_rd_data_valid_r <= 1'h0;
  end
  else if (rdrs_packet.rd_data_valid) begin
    rdrs_packet_rd_data_r <= rdrs_packet.rd_data;
    rdrs_packet_rd_data_valid_r <= 1'h1;
  end
  else begin
    rdrs_packet_rd_data_r <= 64'h0;
    rdrs_packet_rd_data_valid_r <= 1'h0;
  end
end
always_comb begin
  if (cfg_pcfg_tile_connected_next | cfg_pcfg_tile_connected_prev) begin
    rdrq_packet_dma2ring_w.rd_en = rdrq_packet_rd_en_next;
    rdrq_packet_dma2ring_w.rd_addr = rdrq_packet_rd_addr_next;
    rdrq_packet_dma2bank_w.rd_en = 1'h0;
    rdrq_packet_dma2bank_w.rd_addr = 19'h0;
  end
  else begin
    rdrq_packet_dma2ring_w.rd_en = 1'h0;
    rdrq_packet_dma2ring_w.rd_addr = 19'h0;
    rdrq_packet_dma2bank_w.rd_en = rdrq_packet_rd_en_next;
    rdrq_packet_dma2bank_w.rd_addr = rdrq_packet_rd_addr_next;
  end
end
always_comb begin
  if (cfg_pcfg_tile_connected_next | cfg_pcfg_tile_connected_prev) begin
    rdrs_packet = rdrs_packet_ring2dma;
  end
  else rdrs_packet = rdrs_packet_bank2dma;
end
always_comb begin
  cgra_cfg_pcfg.rd_en = 1'h0;
  cgra_cfg_pcfg.wr_en = rdrs_packet_rd_data_valid_r;
  cgra_cfg_pcfg.data = rdrs_packet_rd_data_r[31:0];
  if (cfg_pcfg_dma_ctrl_relocation_is_msb) begin
    cgra_cfg_pcfg.addr = rdrs_packet_rd_data_r[63:32] + 32'(cfg_pcfg_dma_ctrl_relocation_value << 16'h10);
  end
  else cgra_cfg_pcfg.addr = rdrs_packet_rd_data_r[63:32] + 32'(cfg_pcfg_dma_ctrl_relocation_value);
end
assign pcfg_done_pulse = done_pulse_d_arr[4'(cfg_pcfg_network_latency) + 4'h3 + 4'h2];

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    pcfg_dma_done_interrupt <= 1'h0;
  end
  else if (pcfg_done_pulse) begin
    pcfg_dma_done_interrupt <= 1'h1;
  end
  else if (pcfg_done_pulse_last) begin
    pcfg_dma_done_interrupt <= 1'h0;
  end
end
assign clk_en_dma2bank = dma2bank_clk_en;
pipeline_w_1_d_12_array done_pulse_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(done_pulse_r),
  .reset(reset),
  .out_(done_pulse_d_arr)
);

pipeline_w_1_d_5 pcfg_dma_interrupt_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(pcfg_done_pulse),
  .reset(reset),
  .out_(pcfg_done_pulse_last)
);

glb_clk_en_gen_unq0 dma2bank_clk_en_gen (
  .clk(clk),
  .enable(rdrq_packet_dma2bank_w.rd_en),
  .reset(reset),
  .clk_en(dma2bank_clk_en)
);

endmodule   // glb_pcfg_dma

module glb_ring_switch_RD (
  input logic cfg_ld_dma_on,
  input logic cfg_tile_connected_next,
  input logic cfg_tile_connected_prev,
  input logic clk,
  input logic glb_tile_id,
  input rdrq_packet_t rdrq_packet_dma2ring,
  input rdrq_packet_t rdrq_packet_e2w_esti,
  input rdrq_packet_t rdrq_packet_w2e_wsti,
  input rdrs_packet_t rdrs_packet_bank2ring,
  input rdrs_packet_t rdrs_packet_e2w_esti,
  input rdrs_packet_t rdrs_packet_w2e_wsti,
  input logic reset,
  output logic clk_en_ring2bank,
  output rdrq_packet_t rdrq_packet_e2w_wsto,
  output rdrq_packet_t rdrq_packet_ring2bank,
  output rdrq_packet_t rdrq_packet_w2e_esto,
  output rdrs_packet_t rdrs_packet_e2w_wsto,
  output rdrs_packet_t rdrs_packet_ring2dma,
  output rdrs_packet_t rdrs_packet_w2e_esto
);

rdrq_packet_t rdrq_packet_e2w_esti_muxed;
rdrq_packet_t rdrq_packet_e2w_wsto_w;
rdrq_packet_t rdrq_packet_ring2bank_w;
rdrq_packet_t rdrq_packet_w2e_esto_w;
rdrq_packet_t rdrq_packet_w2e_wsti_muxed;
rdrs_packet_t rdrs_packet_e2w_esti_muxed;
rdrs_packet_t rdrs_packet_e2w_wsto_w;
rdrs_packet_t rdrs_packet_ring2dma_w;
rdrs_packet_t rdrs_packet_w2e_esto_w;
rdrs_packet_t rdrs_packet_w2e_wsti_muxed;
logic ring2bank_rd_clk_en;
always_comb begin
  if (cfg_tile_connected_prev) begin
    rdrq_packet_w2e_wsti_muxed = rdrq_packet_w2e_wsti;
    rdrs_packet_w2e_wsti_muxed = rdrs_packet_w2e_wsti;
  end
  else begin
    rdrq_packet_w2e_wsti_muxed = rdrq_packet_e2w_wsto;
    rdrs_packet_w2e_wsti_muxed = rdrs_packet_e2w_wsto;
  end
end
always_comb begin
  if (cfg_tile_connected_next) begin
    rdrq_packet_e2w_esti_muxed = rdrq_packet_e2w_esti;
    rdrs_packet_e2w_esti_muxed = rdrs_packet_e2w_esti;
  end
  else begin
    rdrq_packet_e2w_esti_muxed = rdrq_packet_w2e_esto;
    rdrs_packet_e2w_esti_muxed = rdrs_packet_w2e_esto;
  end
end
always_comb begin
  if (rdrq_packet_dma2ring.rd_en == 1'h1) begin
    if (rdrq_packet_dma2ring.rd_addr[18] == glb_tile_id) begin
      rdrq_packet_ring2bank_w = rdrq_packet_dma2ring;
      rdrq_packet_w2e_esto_w = 20'h0;
    end
    else begin
      rdrq_packet_ring2bank_w = 20'h0;
      rdrq_packet_w2e_esto_w = rdrq_packet_dma2ring;
    end
  end
  else if (rdrq_packet_w2e_wsti_muxed.rd_en == 1'h1) begin
    if (rdrq_packet_w2e_wsti_muxed.rd_addr[18] == glb_tile_id) begin
      rdrq_packet_ring2bank_w = rdrq_packet_w2e_wsti_muxed;
      rdrq_packet_w2e_esto_w = 20'h0;
    end
    else begin
      rdrq_packet_ring2bank_w = 20'h0;
      rdrq_packet_w2e_esto_w = rdrq_packet_w2e_wsti_muxed;
    end
  end
  else begin
    rdrq_packet_ring2bank_w = 20'h0;
    rdrq_packet_w2e_esto_w = 20'h0;
  end
  rdrq_packet_e2w_wsto_w = rdrq_packet_e2w_esti_muxed;
end
always_comb begin
  if (rdrs_packet_bank2ring.rd_data_valid == 1'h1) begin
    rdrs_packet_w2e_esto_w = rdrs_packet_bank2ring;
  end
  else if (rdrs_packet_w2e_wsti_muxed.rd_data_valid & cfg_ld_dma_on) begin
    rdrs_packet_w2e_esto_w = 65'h0;
  end
  else rdrs_packet_w2e_esto_w = rdrs_packet_w2e_wsti_muxed;
  if (rdrs_packet_w2e_wsti_muxed.rd_data_valid & cfg_ld_dma_on) begin
    rdrs_packet_ring2dma_w = rdrs_packet_w2e_wsti_muxed;
  end
  else rdrs_packet_ring2dma_w = 65'h0;
  rdrs_packet_e2w_wsto_w = rdrs_packet_e2w_esti_muxed;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    rdrq_packet_w2e_esto <= 20'h0;
    rdrq_packet_e2w_wsto <= 20'h0;
    rdrq_packet_ring2bank <= 20'h0;
    rdrs_packet_w2e_esto <= 65'h0;
    rdrs_packet_e2w_wsto <= 65'h0;
  end
  else begin
    rdrq_packet_w2e_esto <= rdrq_packet_w2e_esto_w;
    rdrq_packet_e2w_wsto <= rdrq_packet_e2w_wsto_w;
    rdrq_packet_ring2bank <= rdrq_packet_ring2bank_w;
    rdrs_packet_w2e_esto <= rdrs_packet_w2e_esto_w;
    rdrs_packet_e2w_wsto <= rdrs_packet_e2w_wsto_w;
  end
end
always_comb begin
  rdrs_packet_ring2dma = rdrs_packet_ring2dma_w;
end
assign clk_en_ring2bank = ring2bank_rd_clk_en;
glb_clk_en_gen_unq0 ring2bank_rd_clk_en_gen (
  .clk(clk),
  .enable(rdrq_packet_ring2bank_w.rd_en),
  .reset(reset),
  .clk_en(ring2bank_rd_clk_en)
);

endmodule   // glb_ring_switch_RD

module glb_ring_switch_WR_RD (
  input logic cfg_ld_dma_on,
  input logic cfg_tile_connected_next,
  input logic cfg_tile_connected_prev,
  input logic clk,
  input logic glb_tile_id,
  input rdrq_packet_t rdrq_packet_dma2ring,
  input rdrq_packet_t rdrq_packet_e2w_esti,
  input rdrq_packet_t rdrq_packet_w2e_wsti,
  input rdrs_packet_t rdrs_packet_bank2ring,
  input rdrs_packet_t rdrs_packet_e2w_esti,
  input rdrs_packet_t rdrs_packet_w2e_wsti,
  input logic reset,
  input wr_packet_t wr_packet_dma2ring,
  input wr_packet_t wr_packet_e2w_esti,
  input wr_packet_t wr_packet_w2e_wsti,
  output logic clk_en_ring2bank,
  output rdrq_packet_t rdrq_packet_e2w_wsto,
  output rdrq_packet_t rdrq_packet_ring2bank,
  output rdrq_packet_t rdrq_packet_w2e_esto,
  output rdrs_packet_t rdrs_packet_e2w_wsto,
  output rdrs_packet_t rdrs_packet_ring2dma,
  output rdrs_packet_t rdrs_packet_w2e_esto,
  output wr_packet_t wr_packet_e2w_wsto,
  output wr_packet_t wr_packet_ring2bank,
  output wr_packet_t wr_packet_w2e_esto
);

rdrq_packet_t rdrq_packet_e2w_esti_muxed;
rdrq_packet_t rdrq_packet_e2w_wsto_w;
rdrq_packet_t rdrq_packet_ring2bank_w;
rdrq_packet_t rdrq_packet_w2e_esto_w;
rdrq_packet_t rdrq_packet_w2e_wsti_muxed;
rdrs_packet_t rdrs_packet_e2w_esti_muxed;
rdrs_packet_t rdrs_packet_e2w_wsto_w;
rdrs_packet_t rdrs_packet_ring2dma_w;
rdrs_packet_t rdrs_packet_w2e_esto_w;
rdrs_packet_t rdrs_packet_w2e_wsti_muxed;
logic ring2bank_rd_clk_en;
logic ring2bank_wr_clk_en;
wr_packet_t wr_packet_e2w_esti_muxed;
wr_packet_t wr_packet_e2w_wsto_w;
wr_packet_t wr_packet_ring2bank_w;
wr_packet_t wr_packet_w2e_esto_w;
wr_packet_t wr_packet_w2e_wsti_muxed;
always_comb begin
  if (cfg_tile_connected_prev) begin
    wr_packet_w2e_wsti_muxed = wr_packet_w2e_wsti;
    rdrq_packet_w2e_wsti_muxed = rdrq_packet_w2e_wsti;
    rdrs_packet_w2e_wsti_muxed = rdrs_packet_w2e_wsti;
  end
  else begin
    wr_packet_w2e_wsti_muxed = wr_packet_e2w_wsto;
    rdrq_packet_w2e_wsti_muxed = rdrq_packet_e2w_wsto;
    rdrs_packet_w2e_wsti_muxed = rdrs_packet_e2w_wsto;
  end
end
always_comb begin
  if (cfg_tile_connected_next) begin
    wr_packet_e2w_esti_muxed = wr_packet_e2w_esti;
    rdrq_packet_e2w_esti_muxed = rdrq_packet_e2w_esti;
    rdrs_packet_e2w_esti_muxed = rdrs_packet_e2w_esti;
  end
  else begin
    wr_packet_e2w_esti_muxed = wr_packet_w2e_esto;
    rdrq_packet_e2w_esti_muxed = rdrq_packet_w2e_esto;
    rdrs_packet_e2w_esti_muxed = rdrs_packet_w2e_esto;
  end
end
always_comb begin
  if (wr_packet_dma2ring.wr_en == 1'h1) begin
    if (wr_packet_dma2ring.wr_addr[18] == glb_tile_id) begin
      wr_packet_ring2bank_w = wr_packet_dma2ring;
      wr_packet_w2e_esto_w = 92'h0;
    end
    else begin
      wr_packet_ring2bank_w = 92'h0;
      wr_packet_w2e_esto_w = wr_packet_dma2ring;
    end
  end
  else if (wr_packet_w2e_wsti_muxed.wr_en == 1'h1) begin
    if (wr_packet_w2e_wsti_muxed.wr_addr[18] == glb_tile_id) begin
      wr_packet_ring2bank_w = wr_packet_w2e_wsti_muxed;
      wr_packet_w2e_esto_w = 92'h0;
    end
    else begin
      wr_packet_ring2bank_w = 92'h0;
      wr_packet_w2e_esto_w = wr_packet_w2e_wsti_muxed;
    end
  end
  else begin
    wr_packet_ring2bank_w = 92'h0;
    wr_packet_w2e_esto_w = 92'h0;
  end
  wr_packet_e2w_wsto_w = wr_packet_e2w_esti_muxed;
end
always_comb begin
  if (rdrq_packet_dma2ring.rd_en == 1'h1) begin
    if (rdrq_packet_dma2ring.rd_addr[18] == glb_tile_id) begin
      rdrq_packet_ring2bank_w = rdrq_packet_dma2ring;
      rdrq_packet_w2e_esto_w = 20'h0;
    end
    else begin
      rdrq_packet_ring2bank_w = 20'h0;
      rdrq_packet_w2e_esto_w = rdrq_packet_dma2ring;
    end
  end
  else if (rdrq_packet_w2e_wsti_muxed.rd_en == 1'h1) begin
    if (rdrq_packet_w2e_wsti_muxed.rd_addr[18] == glb_tile_id) begin
      rdrq_packet_ring2bank_w = rdrq_packet_w2e_wsti_muxed;
      rdrq_packet_w2e_esto_w = 20'h0;
    end
    else begin
      rdrq_packet_ring2bank_w = 20'h0;
      rdrq_packet_w2e_esto_w = rdrq_packet_w2e_wsti_muxed;
    end
  end
  else begin
    rdrq_packet_ring2bank_w = 20'h0;
    rdrq_packet_w2e_esto_w = 20'h0;
  end
  rdrq_packet_e2w_wsto_w = rdrq_packet_e2w_esti_muxed;
end
always_comb begin
  if (rdrs_packet_bank2ring.rd_data_valid == 1'h1) begin
    rdrs_packet_w2e_esto_w = rdrs_packet_bank2ring;
  end
  else if (rdrs_packet_w2e_wsti_muxed.rd_data_valid & cfg_ld_dma_on) begin
    rdrs_packet_w2e_esto_w = 65'h0;
  end
  else rdrs_packet_w2e_esto_w = rdrs_packet_w2e_wsti_muxed;
  if (rdrs_packet_w2e_wsti_muxed.rd_data_valid & cfg_ld_dma_on) begin
    rdrs_packet_ring2dma_w = rdrs_packet_w2e_wsti_muxed;
  end
  else rdrs_packet_ring2dma_w = 65'h0;
  rdrs_packet_e2w_wsto_w = rdrs_packet_e2w_esti_muxed;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    wr_packet_w2e_esto <= 92'h0;
    wr_packet_e2w_wsto <= 92'h0;
    wr_packet_ring2bank <= 92'h0;
    rdrq_packet_w2e_esto <= 20'h0;
    rdrq_packet_e2w_wsto <= 20'h0;
    rdrq_packet_ring2bank <= 20'h0;
    rdrs_packet_w2e_esto <= 65'h0;
    rdrs_packet_e2w_wsto <= 65'h0;
  end
  else begin
    wr_packet_w2e_esto <= wr_packet_w2e_esto_w;
    wr_packet_e2w_wsto <= wr_packet_e2w_wsto_w;
    wr_packet_ring2bank <= wr_packet_ring2bank_w;
    rdrq_packet_w2e_esto <= rdrq_packet_w2e_esto_w;
    rdrq_packet_e2w_wsto <= rdrq_packet_e2w_wsto_w;
    rdrq_packet_ring2bank <= rdrq_packet_ring2bank_w;
    rdrs_packet_w2e_esto <= rdrs_packet_w2e_esto_w;
    rdrs_packet_e2w_wsto <= rdrs_packet_e2w_wsto_w;
  end
end
always_comb begin
  rdrs_packet_ring2dma = rdrs_packet_ring2dma_w;
end
assign clk_en_ring2bank = ring2bank_wr_clk_en | ring2bank_rd_clk_en;
glb_clk_en_gen ring2bank_wr_clk_en_gen (
  .clk(clk),
  .enable(wr_packet_ring2bank_w.wr_en),
  .reset(reset),
  .clk_en(ring2bank_wr_clk_en)
);

glb_clk_en_gen_unq0 ring2bank_rd_clk_en_gen (
  .clk(clk),
  .enable(rdrq_packet_ring2bank_w.rd_en),
  .reset(reset),
  .clk_en(ring2bank_rd_clk_en)
);

endmodule   // glb_ring_switch_WR_RD

module glb_sched_gen (
  input logic clk,
  input logic clk_en,
  input logic [15:0] current_addr,
  input logic [15:0] cycle_count,
  input logic finished,
  input logic reset,
  input logic restart,
  output logic valid_output
);

logic valid_gate;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    valid_gate <= 1'h1;
  end
  else if (clk_en) begin
    if (restart) begin
      valid_gate <= 1'h0;
    end
    else if (finished) begin
      valid_gate <= 1'h1;
    end
  end
end
always_comb begin
  valid_output = (cycle_count == current_addr) & (~valid_gate);
end
endmodule   // glb_sched_gen

module glb_store_dma (
  input logic [1:0] cfg_data_network_f2g_mux,
  input logic [5:0] cfg_data_network_latency,
  input logic [1:0] cfg_st_dma_ctrl_mode,
  input logic cfg_st_dma_ctrl_use_valid,
  input dma_header_t cfg_st_dma_header,
  input logic cfg_st_dma_num_repeat,
  input logic cfg_tile_connected_next,
  input logic cfg_tile_connected_prev,
  input logic clk,
  input logic [1:0] [15:0] data_f2g,
  input logic [1:0] data_valid_f2g,
  input logic reset,
  input logic st_dma_start_pulse,
  output logic clk_en_dma2bank,
  output logic st_dma_done_interrupt,
  output wr_packet_t wr_packet_dma2bank,
  output wr_packet_t wr_packet_dma2ring
);

logic bank_addr_match;
logic [18:0] bank_wr_addr;
logic [63:0] bank_wr_data_cache_r;
logic [63:0] bank_wr_data_cache_w;
logic bank_wr_en;
logic [7:0] bank_wr_strb_cache_r;
logic [7:0] bank_wr_strb_cache_w;
dma_header_t current_dma_header;
logic [15:0] cycle_count;
logic [15:0] cycle_current_addr;
logic [7:0][15:0] cycle_stride_addr_gen_strides;
logic cycle_valid;
logic cycle_valid_muxed;
logic [19:0] data_current_addr;
logic [1:0][15:0] data_f2g_r;
logic [19:0] data_stride_addr_gen_start_addr;
logic [7:0][19:0] data_stride_addr_gen_strides;
logic [1:0] data_valid_f2g_r;
logic dma2bank_clk_en;
logic done_pulse_d_arr [7:0];
logic done_pulse_w;
logic is_first;
logic is_last;
logic [18:0] last_strm_wr_addr_r;
logic loop_done;
logic [7:0][31:0] loop_iter_ranges;
logic [2:0] loop_mux_sel;
logic repeat_cnt;
logic st_dma_done_pulse;
logic st_dma_done_pulse_last;
logic st_dma_start_pulse_next;
logic st_dma_start_pulse_r;
logic [15:0] strm_data;
logic [1:0] strm_data_sel;
logic strm_data_valid;
logic strm_run;
logic [18:0] strm_wr_addr_w;
logic [15:0] strm_wr_data_w;
logic strm_wr_en_w;
wr_packet_t wr_packet_dma2bank_w;
wr_packet_t wr_packet_dma2ring_w;
assign current_dma_header = cfg_st_dma_header;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    repeat_cnt <= 1'h0;
  end
  else if (cfg_st_dma_ctrl_mode == 2'h2) begin
    if (st_dma_done_pulse) begin
      if ((repeat_cnt + 1'h1) < cfg_st_dma_num_repeat) begin
        repeat_cnt <= repeat_cnt + 1'h1;
      end
    end
  end
  else if (cfg_st_dma_ctrl_mode == 2'h3) begin
    if (st_dma_done_pulse) begin
      if (((repeat_cnt + 1'h1) < cfg_st_dma_num_repeat) & ((repeat_cnt + 1'h1) < 1'h1)) begin
        repeat_cnt <= repeat_cnt + 1'h1;
      end
    end
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    is_first <= 1'h0;
  end
  else if (st_dma_start_pulse_r) begin
    is_first <= 1'h1;
  end
  else if (strm_wr_en_w) begin
    is_first <= 1'h0;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    is_last <= 1'h0;
  end
  else if (loop_done) begin
    is_last <= 1'h1;
  end
  else if (bank_wr_en) begin
    is_last <= 1'h0;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    strm_run <= 1'h0;
  end
  else if (st_dma_start_pulse_r) begin
    strm_run <= 1'h1;
  end
  else if (loop_done) begin
    strm_run <= 1'h0;
  end
end
always_comb begin
  if (cfg_st_dma_ctrl_mode == 2'h0) begin
    st_dma_start_pulse_next = 1'h0;
  end
  else if (cfg_st_dma_ctrl_mode == 2'h1) begin
    st_dma_start_pulse_next = (~strm_run) & st_dma_start_pulse;
  end
  else if ((cfg_st_dma_ctrl_mode == 2'h2) | (cfg_st_dma_ctrl_mode == 2'h3)) begin
    st_dma_start_pulse_next = ((~strm_run) & st_dma_start_pulse) | (st_dma_done_pulse & ((repeat_cnt + 1'h1) <
        cfg_st_dma_num_repeat));
  end
  else st_dma_start_pulse_next = 1'h0;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    st_dma_start_pulse_r <= 1'h0;
  end
  else if (st_dma_start_pulse_r) begin
    st_dma_start_pulse_r <= 1'h0;
  end
  else st_dma_start_pulse_r <= st_dma_start_pulse_next;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    cycle_count <= 16'h0;
  end
  else if (st_dma_start_pulse_r) begin
    cycle_count <= 16'h0;
  end
  else if (loop_done) begin
    cycle_count <= 16'h0;
  end
  else if (strm_run) begin
    cycle_count <= cycle_count + 16'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    data_f2g_r <= 32'h0;
    data_valid_f2g_r <= 2'h0;
  end
  else begin
    data_f2g_r[0] <= data_f2g[0];
    data_f2g_r[1] <= data_f2g[1];
    data_valid_f2g_r <= data_valid_f2g;
  end
end
always_comb begin
  strm_data = 16'h0;
  strm_data_valid = 1'h0;
  if (cfg_data_network_f2g_mux[0] == 1'h1) begin
    strm_data = data_f2g_r[0];
    strm_data_valid = data_valid_f2g_r[0];
  end
  else begin
    strm_data = strm_data;
    strm_data_valid = strm_data_valid;
  end
  if (cfg_data_network_f2g_mux[1] == 1'h1) begin
    strm_data = data_f2g_r[1];
    strm_data_valid = data_valid_f2g_r[1];
  end
  else begin
    strm_data = strm_data;
    strm_data_valid = strm_data_valid;
  end
end
always_comb begin
  if (cfg_st_dma_ctrl_use_valid) begin
    cycle_valid_muxed = strm_data_valid;
  end
  else cycle_valid_muxed = cycle_valid;
end
always_comb begin
  strm_wr_en_w = cycle_valid_muxed;
  strm_wr_addr_w = 19'(data_current_addr);
  strm_wr_data_w = strm_data;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    last_strm_wr_addr_r <= 19'h0;
  end
  else if (strm_wr_en_w) begin
    last_strm_wr_addr_r <= strm_wr_addr_w;
  end
end
always_comb begin
  strm_data_sel = strm_wr_addr_w[2:1];
end
always_comb begin
  bank_wr_strb_cache_w = bank_wr_strb_cache_r;
  bank_wr_data_cache_w = bank_wr_data_cache_r;
  if (bank_wr_en) begin
    bank_wr_strb_cache_w = 8'h0;
    bank_wr_data_cache_w = 64'h0;
  end
  if (strm_wr_en_w) begin
    if (strm_data_sel == 2'h0) begin
      bank_wr_strb_cache_w[1:0] = 2'h3;
      bank_wr_data_cache_w[15:0] = strm_wr_data_w;
    end
    else if (strm_data_sel == 2'h1) begin
      bank_wr_strb_cache_w[3:2] = 2'h3;
      bank_wr_data_cache_w[31:16] = strm_wr_data_w;
    end
    else if (strm_data_sel == 2'h2) begin
      bank_wr_strb_cache_w[5:4] = 2'h3;
      bank_wr_data_cache_w[47:32] = strm_wr_data_w;
    end
    else if (strm_data_sel == 2'h3) begin
      bank_wr_strb_cache_w[7:6] = 2'h3;
      bank_wr_data_cache_w[63:48] = strm_wr_data_w;
    end
    else begin
      bank_wr_strb_cache_w = bank_wr_strb_cache_r;
      bank_wr_data_cache_w = bank_wr_data_cache_r;
    end
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    bank_wr_strb_cache_r <= 8'h0;
    bank_wr_data_cache_r <= 64'h0;
  end
  else begin
    bank_wr_strb_cache_r <= bank_wr_strb_cache_w;
    bank_wr_data_cache_r <= bank_wr_data_cache_w;
  end
end
always_comb begin
  bank_addr_match = strm_wr_addr_w[18:3] == last_strm_wr_addr_r[18:3];
  bank_wr_en = (strm_wr_en_w & (~bank_addr_match) & (~is_first)) | is_last;
  bank_wr_addr = last_strm_wr_addr_r;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    wr_packet_dma2bank <= 92'h0;
    wr_packet_dma2ring <= 92'h0;
  end
  else begin
    wr_packet_dma2bank <= wr_packet_dma2bank_w;
    wr_packet_dma2ring <= wr_packet_dma2ring_w;
  end
end
always_comb begin
  if (cfg_tile_connected_next | cfg_tile_connected_prev) begin
    wr_packet_dma2bank_w = 92'h0;
    wr_packet_dma2ring_w.wr_en = bank_wr_en;
    wr_packet_dma2ring_w.wr_strb = bank_wr_strb_cache_r;
    wr_packet_dma2ring_w.wr_data = bank_wr_data_cache_r;
    wr_packet_dma2ring_w.wr_addr = bank_wr_addr;
  end
  else begin
    wr_packet_dma2bank_w.wr_en = bank_wr_en;
    wr_packet_dma2bank_w.wr_strb = bank_wr_strb_cache_r;
    wr_packet_dma2bank_w.wr_data = bank_wr_data_cache_r;
    wr_packet_dma2bank_w.wr_addr = bank_wr_addr;
    wr_packet_dma2ring_w = 92'h0;
  end
end
assign clk_en_dma2bank = dma2bank_clk_en;
always_comb begin
  done_pulse_w = loop_done & strm_run;
end
assign st_dma_done_pulse = done_pulse_d_arr[3'(cfg_data_network_latency) + 3'h1];

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    st_dma_done_interrupt <= 1'h0;
  end
  else if (st_dma_done_pulse) begin
    st_dma_done_interrupt <= 1'h1;
  end
  else if (st_dma_done_pulse_last) begin
    st_dma_done_interrupt <= 1'h0;
  end
end
assign loop_iter_ranges[0] = current_dma_header.range_0;
assign loop_iter_ranges[1] = current_dma_header.range_1;
assign loop_iter_ranges[2] = current_dma_header.range_2;
assign loop_iter_ranges[3] = current_dma_header.range_3;
assign loop_iter_ranges[4] = current_dma_header.range_4;
assign loop_iter_ranges[5] = current_dma_header.range_5;
assign loop_iter_ranges[6] = current_dma_header.range_6;
assign loop_iter_ranges[7] = current_dma_header.range_7;
assign cycle_stride_addr_gen_strides[0] = current_dma_header.cycle_stride_0;
assign cycle_stride_addr_gen_strides[1] = current_dma_header.cycle_stride_1;
assign cycle_stride_addr_gen_strides[2] = current_dma_header.cycle_stride_2;
assign cycle_stride_addr_gen_strides[3] = current_dma_header.cycle_stride_3;
assign cycle_stride_addr_gen_strides[4] = current_dma_header.cycle_stride_4;
assign cycle_stride_addr_gen_strides[5] = current_dma_header.cycle_stride_5;
assign cycle_stride_addr_gen_strides[6] = current_dma_header.cycle_stride_6;
assign cycle_stride_addr_gen_strides[7] = current_dma_header.cycle_stride_7;
assign data_stride_addr_gen_start_addr = 20'(current_dma_header.start_addr);
assign data_stride_addr_gen_strides[0] = current_dma_header.stride_0;
assign data_stride_addr_gen_strides[1] = current_dma_header.stride_1;
assign data_stride_addr_gen_strides[2] = current_dma_header.stride_2;
assign data_stride_addr_gen_strides[3] = current_dma_header.stride_3;
assign data_stride_addr_gen_strides[4] = current_dma_header.stride_4;
assign data_stride_addr_gen_strides[5] = current_dma_header.stride_5;
assign data_stride_addr_gen_strides[6] = current_dma_header.stride_6;
assign data_stride_addr_gen_strides[7] = current_dma_header.stride_7;
glb_clk_en_gen dma2bank_clk_en_gen (
  .clk(clk),
  .enable(wr_packet_dma2bank_w.wr_en),
  .reset(reset),
  .clk_en(dma2bank_clk_en)
);

pipeline_w_1_d_8_array done_pulse_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(done_pulse_w),
  .reset(reset),
  .out_(done_pulse_d_arr)
);

pipeline_w_1_d_5 st_dma_interrupt_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(st_dma_done_pulse),
  .reset(reset),
  .out_(st_dma_done_pulse_last)
);

glb_loop_iter loop_iter (
  .clk(clk),
  .clk_en(1'h1),
  .dim(current_dma_header.dim),
  .ranges(loop_iter_ranges),
  .reset(reset),
  .step(cycle_valid_muxed),
  .mux_sel_out(loop_mux_sel),
  .restart(loop_done)
);

glb_sched_gen cycle_stride_sched_gen (
  .clk(clk),
  .clk_en(1'h1),
  .current_addr(cycle_current_addr),
  .cycle_count(cycle_count),
  .finished(loop_done),
  .reset(reset),
  .restart(st_dma_start_pulse_r),
  .valid_output(cycle_valid)
);

glb_addr_gen #(
  .addr_width(32'h10))
cycle_stride_addr_gen (
  .clk(clk),
  .clk_en(1'h1),
  .mux_sel(loop_mux_sel),
  .reset(reset),
  .restart(st_dma_start_pulse_r),
  .start_addr(current_dma_header.cycle_start_addr),
  .step(cycle_valid_muxed),
  .strides(cycle_stride_addr_gen_strides),
  .addr_out(cycle_current_addr)
);

glb_addr_gen #(
  .addr_width(32'h14))
data_stride_addr_gen (
  .clk(clk),
  .clk_en(1'h1),
  .mux_sel(loop_mux_sel),
  .reset(reset),
  .restart(st_dma_start_pulse_r),
  .start_addr(data_stride_addr_gen_start_addr),
  .step(cycle_valid_muxed),
  .strides(data_stride_addr_gen_strides),
  .addr_out(data_current_addr)
);

endmodule   // glb_store_dma

module glb_switch (
  glb_tile_ifc_A_19_D_64.master if_est_m,
  glb_tile_ifc_A_19_D_64.slave if_wst_s,
  input logic gclk,
  input logic glb_tile_id,
  input logic mclk,
  input rdrs_packet_t rdrs_packet,
  input logic reset,
  output logic clk_en_sw2bank,
  output rdrq_packet_t rdrq_packet,
  output wr_packet_t wr_packet
);

logic [18:0] bank_rd_addr;
logic bank_rd_en;
logic [18:0] bank_wr_addr;
logic [63:0] bank_wr_data;
logic bank_wr_en;
logic [7:0] bank_wr_strb;
logic [18:0] if_est_m_rd_addr_w;
logic if_est_m_rd_clk_en_sel;
logic if_est_m_rd_clk_en_sel_first_cycle;
logic if_est_m_rd_clk_en_sel_latch;
logic if_est_m_rd_en_w;
logic [18:0] if_est_m_wr_addr_w;
logic if_est_m_wr_clk_en_sel;
logic if_est_m_wr_clk_en_sel_first_cycle;
logic if_est_m_wr_clk_en_sel_latch;
logic [63:0] if_est_m_wr_data_w;
logic if_est_m_wr_en_w;
logic [7:0] if_est_m_wr_strb_w;
logic if_wst_s_rd_clk_en_d;
logic if_wst_s_wr_clk_en_d;
logic rd_data_valid_w;
logic [63:0] rd_data_w;
logic rd_tile_id_match;
logic sw2bank_rd_clk_en;
logic sw2bank_rd_clk_en_gen_enable;
logic sw2bank_wr_clk_en;
logic sw2bank_wr_clk_en_gen_enable;
logic wr_tile_id_match;
always_comb begin
  wr_tile_id_match = glb_tile_id == if_wst_s.wr_addr[18];
  rd_tile_id_match = glb_tile_id == if_wst_s.rd_addr[18];
end
always_comb begin
  if (if_wst_s.wr_en) begin
    if (wr_tile_id_match) begin
      if_est_m_wr_en_w = 1'h0;
      if_est_m_wr_addr_w = 19'h0;
      if_est_m_wr_data_w = 64'h0;
      if_est_m_wr_strb_w = 8'h0;
      bank_wr_en = 1'h1;
      bank_wr_addr = if_wst_s.wr_addr;
      bank_wr_data = if_wst_s.wr_data;
      bank_wr_strb = if_wst_s.wr_strb;
    end
    else begin
      if_est_m_wr_en_w = if_wst_s.wr_en;
      if_est_m_wr_addr_w = if_wst_s.wr_addr;
      if_est_m_wr_data_w = if_wst_s.wr_data;
      if_est_m_wr_strb_w = if_wst_s.wr_strb;
      bank_wr_en = 1'h0;
      bank_wr_addr = 19'h0;
      bank_wr_data = 64'h0;
      bank_wr_strb = 8'h0;
    end
  end
  else begin
    if_est_m_wr_en_w = 1'h0;
    if_est_m_wr_addr_w = 19'h0;
    if_est_m_wr_data_w = 64'h0;
    if_est_m_wr_strb_w = 8'h0;
    bank_wr_en = 1'h0;
    bank_wr_addr = 19'h0;
    bank_wr_data = 64'h0;
    bank_wr_strb = 8'h0;
  end
end
always_comb begin
  if (if_wst_s.rd_en) begin
    if (rd_tile_id_match) begin
      if_est_m_rd_en_w = 1'h0;
      if_est_m_rd_addr_w = 19'h0;
      bank_rd_en = 1'h1;
      bank_rd_addr = if_wst_s.rd_addr;
    end
    else begin
      if_est_m_rd_en_w = if_wst_s.rd_en;
      if_est_m_rd_addr_w = if_wst_s.rd_addr;
      bank_rd_en = 1'h0;
      bank_rd_addr = 19'h0;
    end
  end
  else begin
    if_est_m_rd_en_w = 1'h0;
    if_est_m_rd_addr_w = 19'h0;
    bank_rd_en = 1'h0;
    bank_rd_addr = 19'h0;
  end
end
always_comb begin
  rd_data_w = 64'h0;
  rd_data_valid_w = 1'h0;
  if (rdrs_packet.rd_data_valid == 1'h1) begin
    rd_data_w = rdrs_packet.rd_data;
    rd_data_valid_w = 1'h1;
  end
  else if (if_est_m.rd_data_valid == 1'h1) begin
    rd_data_w = if_est_m.rd_data;
    rd_data_valid_w = 1'h1;
  end
end

always_ff @(posedge gclk, posedge reset) begin
  if (reset) begin
    if_est_m.wr_en <= 1'h0;
    if_est_m.wr_strb <= 8'h0;
    if_est_m.wr_addr <= 19'h0;
    if_est_m.wr_data <= 64'h0;
    if_est_m.rd_en <= 1'h0;
    if_est_m.rd_addr <= 19'h0;
    if_wst_s.rd_data <= 64'h0;
    if_wst_s.rd_data_valid <= 1'h0;
    wr_packet.wr_en <= 1'h0;
    wr_packet.wr_strb <= 8'h0;
    wr_packet.wr_addr <= 19'h0;
    wr_packet.wr_data <= 64'h0;
    rdrq_packet.rd_en <= 1'h0;
    rdrq_packet.rd_addr <= 19'h0;
  end
  else begin
    if_est_m.wr_en <= if_est_m_wr_en_w;
    if_est_m.wr_strb <= if_est_m_wr_strb_w;
    if_est_m.wr_addr <= if_est_m_wr_addr_w;
    if_est_m.wr_data <= if_est_m_wr_data_w;
    if_est_m.rd_en <= if_est_m_rd_en_w;
    if_est_m.rd_addr <= if_est_m_rd_addr_w;
    if_wst_s.rd_data <= rd_data_w;
    if_wst_s.rd_data_valid <= rd_data_valid_w;
    wr_packet.wr_en <= bank_wr_en;
    wr_packet.wr_strb <= bank_wr_strb;
    wr_packet.wr_addr <= bank_wr_addr;
    wr_packet.wr_data <= bank_wr_data;
    rdrq_packet.rd_en <= bank_rd_en;
    rdrq_packet.rd_addr <= bank_rd_addr;
  end
end

always_ff @(posedge mclk, posedge reset) begin
  if (reset) begin
    if_wst_s_wr_clk_en_d <= 1'h0;
    if_wst_s_rd_clk_en_d <= 1'h0;
  end
  else begin
    if_wst_s_wr_clk_en_d <= if_wst_s.wr_clk_en;
    if_wst_s_rd_clk_en_d <= if_wst_s.rd_clk_en;
  end
end
always_comb begin
  if_est_m_wr_clk_en_sel_first_cycle = if_wst_s.wr_en & (~wr_tile_id_match);
  if_est_m_rd_clk_en_sel_first_cycle = if_wst_s.rd_en & (~rd_tile_id_match);
end

always_ff @(posedge mclk, posedge reset) begin
  if (reset) begin
    if_est_m_wr_clk_en_sel_latch <= 1'h0;
  end
  else if (if_wst_s.wr_en == 1'h1) begin
    if (wr_tile_id_match) begin
      if_est_m_wr_clk_en_sel_latch <= 1'h0;
    end
    else if_est_m_wr_clk_en_sel_latch <= 1'h1;
  end
  else if (if_wst_s.wr_clk_en == 1'h0) begin
    if_est_m_wr_clk_en_sel_latch <= 1'h0;
  end
end

always_ff @(posedge mclk, posedge reset) begin
  if (reset) begin
    if_est_m_rd_clk_en_sel_latch <= 1'h0;
  end
  else if (if_wst_s.rd_en == 1'h1) begin
    if (rd_tile_id_match) begin
      if_est_m_rd_clk_en_sel_latch <= 1'h0;
    end
    else if_est_m_rd_clk_en_sel_latch <= 1'h1;
  end
  else if (if_wst_s.rd_clk_en == 1'h0) begin
    if_est_m_rd_clk_en_sel_latch <= 1'h0;
  end
end
always_comb begin
  if_est_m_wr_clk_en_sel = if_est_m_wr_clk_en_sel_first_cycle | if_est_m_wr_clk_en_sel_latch;
  if_est_m_rd_clk_en_sel = if_est_m_rd_clk_en_sel_first_cycle | if_est_m_rd_clk_en_sel_latch;
end
always_comb begin
  if (if_est_m_wr_clk_en_sel) begin
    if_est_m.wr_clk_en = if_wst_s_wr_clk_en_d;
  end
  else if_est_m.wr_clk_en = 1'h0;
end
always_comb begin
  if (if_est_m_rd_clk_en_sel) begin
    if_est_m.rd_clk_en = if_wst_s_rd_clk_en_d;
  end
  else if_est_m.rd_clk_en = 1'h0;
end
assign sw2bank_wr_clk_en_gen_enable = if_wst_s.wr_en & wr_tile_id_match;
assign sw2bank_rd_clk_en_gen_enable = if_wst_s.rd_en & rd_tile_id_match;
assign clk_en_sw2bank = sw2bank_wr_clk_en | sw2bank_rd_clk_en;
glb_clk_en_gen sw2bank_wr_clk_en_gen (
  .clk(mclk),
  .enable(sw2bank_wr_clk_en_gen_enable),
  .reset(reset),
  .clk_en(sw2bank_wr_clk_en)
);

glb_clk_en_gen_unq0 sw2bank_rd_clk_en_gen (
  .clk(mclk),
  .enable(sw2bank_rd_clk_en_gen_enable),
  .reset(reset),
  .clk_en(sw2bank_rd_clk_en)
);

endmodule   // glb_switch

module glb_tile (
  input logic cfg_pcfg_tile_connected_wsti,
  input logic cfg_tile_connected_wsti,
  input logic [31:0] cgra_cfg_jtag_addr_bypass_wsti,
  input logic [31:0] cgra_cfg_jtag_addr_wsti,
  input logic [31:0] cgra_cfg_jtag_data_wsti,
  input logic cgra_cfg_jtag_rd_en_bypass_wsti,
  input logic cgra_cfg_jtag_rd_en_wsti,
  input logic cgra_cfg_jtag_wr_en_wsti,
  input logic [31:0] cgra_cfg_pcfg_addr_e2w_esti,
  input logic [31:0] cgra_cfg_pcfg_addr_w2e_wsti,
  input logic [31:0] cgra_cfg_pcfg_data_e2w_esti,
  input logic [31:0] cgra_cfg_pcfg_data_w2e_wsti,
  input logic cgra_cfg_pcfg_rd_en_e2w_esti,
  input logic cgra_cfg_pcfg_rd_en_w2e_wsti,
  input logic cgra_cfg_pcfg_wr_en_e2w_esti,
  input logic cgra_cfg_pcfg_wr_en_w2e_wsti,
  input logic clk,
  input logic clk_en_bank_master,
  input logic clk_en_master,
  input logic clk_en_pcfg_broadcast,
  input logic glb_tile_id,
  input logic [31:0] if_cfg_est_m_rd_data,
  input logic if_cfg_est_m_rd_data_valid,
  input logic [11:0] if_cfg_wst_s_rd_addr,
  input logic if_cfg_wst_s_rd_clk_en,
  input logic if_cfg_wst_s_rd_en,
  input logic [11:0] if_cfg_wst_s_wr_addr,
  input logic if_cfg_wst_s_wr_clk_en,
  input logic [31:0] if_cfg_wst_s_wr_data,
  input logic if_cfg_wst_s_wr_en,
  input logic [63:0] if_proc_est_m_rd_data,
  input logic if_proc_est_m_rd_data_valid,
  input logic [18:0] if_proc_wst_s_rd_addr,
  input logic if_proc_wst_s_rd_clk_en,
  input logic if_proc_wst_s_rd_en,
  input logic [18:0] if_proc_wst_s_wr_addr,
  input logic if_proc_wst_s_wr_clk_en,
  input logic [63:0] if_proc_wst_s_wr_data,
  input logic if_proc_wst_s_wr_en,
  input logic [7:0] if_proc_wst_s_wr_strb,
  input logic [18:0] pcfg_rd_addr_e2w_esti,
  input logic [18:0] pcfg_rd_addr_w2e_wsti,
  input logic [63:0] pcfg_rd_data_e2w_esti,
  input logic pcfg_rd_data_valid_e2w_esti,
  input logic pcfg_rd_data_valid_w2e_wsti,
  input logic [63:0] pcfg_rd_data_w2e_wsti,
  input logic pcfg_rd_en_e2w_esti,
  input logic pcfg_rd_en_w2e_wsti,
  input logic pcfg_start_pulse,
  input logic reset,
  input logic [1:0] [15:0] strm_data_f2g,
  input logic [1:0] strm_data_valid_f2g,
  input logic strm_f2g_start_pulse,
  input logic strm_g2f_start_pulse,
  input logic [18:0] strm_rd_addr_e2w_esti,
  input logic [18:0] strm_rd_addr_w2e_wsti,
  input logic [63:0] strm_rd_data_e2w_esti,
  input logic strm_rd_data_valid_e2w_esti,
  input logic strm_rd_data_valid_w2e_wsti,
  input logic [63:0] strm_rd_data_w2e_wsti,
  input logic strm_rd_en_e2w_esti,
  input logic strm_rd_en_w2e_wsti,
  input logic [18:0] strm_wr_addr_e2w_esti,
  input logic [18:0] strm_wr_addr_w2e_wsti,
  input logic [63:0] strm_wr_data_e2w_esti,
  input logic [63:0] strm_wr_data_w2e_wsti,
  input logic strm_wr_en_e2w_esti,
  input logic strm_wr_en_w2e_wsti,
  input logic [7:0] strm_wr_strb_e2w_esti,
  input logic [7:0] strm_wr_strb_w2e_wsti,
  output logic cfg_pcfg_tile_connected_esto,
  output logic cfg_tile_connected_esto,
  output logic [1:0] [31:0] cgra_cfg_g2f_cfg_addr,
  output logic [1:0] [31:0] cgra_cfg_g2f_cfg_data,
  output logic [1:0] cgra_cfg_g2f_cfg_rd_en,
  output logic [1:0] cgra_cfg_g2f_cfg_wr_en,
  output logic [31:0] cgra_cfg_jtag_addr_bypass_esto,
  output logic [31:0] cgra_cfg_jtag_addr_esto,
  output logic [31:0] cgra_cfg_jtag_data_esto,
  output logic cgra_cfg_jtag_rd_en_bypass_esto,
  output logic cgra_cfg_jtag_rd_en_esto,
  output logic cgra_cfg_jtag_wr_en_esto,
  output logic [31:0] cgra_cfg_pcfg_addr_e2w_wsto,
  output logic [31:0] cgra_cfg_pcfg_addr_w2e_esto,
  output logic [31:0] cgra_cfg_pcfg_data_e2w_wsto,
  output logic [31:0] cgra_cfg_pcfg_data_w2e_esto,
  output logic cgra_cfg_pcfg_rd_en_e2w_wsto,
  output logic cgra_cfg_pcfg_rd_en_w2e_esto,
  output logic cgra_cfg_pcfg_wr_en_e2w_wsto,
  output logic cgra_cfg_pcfg_wr_en_w2e_esto,
  output logic data_flush,
  output logic [11:0] if_cfg_est_m_rd_addr,
  output logic if_cfg_est_m_rd_clk_en,
  output logic if_cfg_est_m_rd_en,
  output logic [11:0] if_cfg_est_m_wr_addr,
  output logic if_cfg_est_m_wr_clk_en,
  output logic [31:0] if_cfg_est_m_wr_data,
  output logic if_cfg_est_m_wr_en,
  output logic [31:0] if_cfg_wst_s_rd_data,
  output logic if_cfg_wst_s_rd_data_valid,
  output logic [18:0] if_proc_est_m_rd_addr,
  output logic if_proc_est_m_rd_clk_en,
  output logic if_proc_est_m_rd_en,
  output logic [18:0] if_proc_est_m_wr_addr,
  output logic if_proc_est_m_wr_clk_en,
  output logic [63:0] if_proc_est_m_wr_data,
  output logic if_proc_est_m_wr_en,
  output logic [7:0] if_proc_est_m_wr_strb,
  output logic [63:0] if_proc_wst_s_rd_data,
  output logic if_proc_wst_s_rd_data_valid,
  output logic pcfg_g2f_interrupt_pulse,
  output logic [18:0] pcfg_rd_addr_e2w_wsto,
  output logic [18:0] pcfg_rd_addr_w2e_esto,
  output logic [63:0] pcfg_rd_data_e2w_wsto,
  output logic pcfg_rd_data_valid_e2w_wsto,
  output logic pcfg_rd_data_valid_w2e_esto,
  output logic [63:0] pcfg_rd_data_w2e_esto,
  output logic pcfg_rd_en_e2w_wsto,
  output logic pcfg_rd_en_w2e_esto,
  output logic [1:0] [15:0] strm_data_g2f,
  output logic [1:0] strm_data_valid_g2f,
  output logic strm_f2g_interrupt_pulse,
  output logic strm_g2f_interrupt_pulse,
  output logic [18:0] strm_rd_addr_e2w_wsto,
  output logic [18:0] strm_rd_addr_w2e_esto,
  output logic [63:0] strm_rd_data_e2w_wsto,
  output logic strm_rd_data_valid_e2w_wsto,
  output logic strm_rd_data_valid_w2e_esto,
  output logic [63:0] strm_rd_data_w2e_esto,
  output logic strm_rd_en_e2w_wsto,
  output logic strm_rd_en_w2e_esto,
  output logic [18:0] strm_wr_addr_e2w_wsto,
  output logic [18:0] strm_wr_addr_w2e_esto,
  output logic [63:0] strm_wr_data_e2w_wsto,
  output logic [63:0] strm_wr_data_w2e_esto,
  output logic strm_wr_en_e2w_wsto,
  output logic strm_wr_en_w2e_esto,
  output logic [7:0] strm_wr_strb_e2w_wsto,
  output logic [7:0] strm_wr_strb_w2e_esto
);

load_dma_ctrl_t cfg_ld_dma_ctrl;
dma_header_t cfg_ld_dma_header;
pcfg_broadcast_mux_t cfg_pcfg_broadcast_mux;
pcfg_dma_ctrl_t cfg_pcfg_dma_ctrl;
pcfg_dma_header_t cfg_pcfg_dma_header;
logic cfg_pcfg_tile_connected_next;
logic cfg_pcfg_tile_connected_prev;
store_dma_ctrl_t cfg_st_dma_ctrl;
dma_header_t cfg_st_dma_header;
logic cfg_tile_connected_next;
logic cfg_tile_connected_prev;
cgra_cfg_t [1:0] cgra_cfg_g2f_cfg_w;
cgra_cfg_t cgra_cfg_pcfgdma2mux;
logic clk_en_bank;
logic clk_en_cfg;
logic clk_en_ld_dma;
logic clk_en_lddma2bank;
logic clk_en_pcfg_dma;
logic clk_en_pcfg_switch;
logic clk_en_pcfgdma2bank;
logic clk_en_pcfgring2bank;
logic clk_en_proc_switch;
logic clk_en_procsw2bank;
logic clk_en_ring2bank;
logic clk_en_st_dma;
logic clk_en_stdma2bank;
logic clk_en_strm_switch;
logic gclk_bank;
logic gclk_cfg;
logic gclk_ld_dma;
logic gclk_pcfg_broadcast;
logic gclk_pcfg_dma;
logic gclk_pcfg_switch;
logic gclk_proc_switch;
logic gclk_st_dma;
logic gclk_strm_switch;
logic glb_bank_0_clk;
rdrs_packet_t glb_bank_0_rdrs_packet;
logic glb_bank_1_clk;
rdrs_packet_t glb_bank_1_rdrs_packet;
logic glb_bank_mux_clk;
cfg_data_network_t glb_cfg_cfg_data_network;
cfg_pcfg_network_t glb_cfg_cfg_pcfg_network;
logic glb_cfg_gclk;
logic glb_clk_gate_bank_enable;
logic glb_clk_gate_cfg_enable;
logic glb_clk_gate_ld_dma_enable;
logic glb_clk_gate_pcfg_broadcast_enable;
logic glb_clk_gate_pcfg_dma_enable;
logic glb_clk_gate_pcfg_switch_enable;
logic glb_clk_gate_proc_switch_enable;
logic glb_clk_gate_st_dma_enable;
logic glb_clk_gate_strm_switch_enable;
logic glb_load_dma_clk;
cgra_cfg_t glb_pcfg_broadcast_cgra_cfg_jtag_esto;
cgra_cfg_t glb_pcfg_broadcast_cgra_cfg_jtag_wsti;
cgra_cfg_t glb_pcfg_broadcast_cgra_cfg_pcfg_esti;
cgra_cfg_t glb_pcfg_broadcast_cgra_cfg_pcfg_esto;
cgra_cfg_t glb_pcfg_broadcast_cgra_cfg_pcfg_wsti;
cgra_cfg_t glb_pcfg_broadcast_cgra_cfg_pcfg_wsto;
logic glb_pcfg_broadcast_clk;
logic glb_pcfg_dma_clk;
logic glb_pcfg_ring_switch_cfg_ld_dma_on;
logic glb_pcfg_ring_switch_clk;
logic glb_proc_switch_gclk;
logic glb_store_dma_clk;
logic glb_strm_ring_switch_cfg_ld_dma_on;
logic glb_strm_ring_switch_clk;
rdrq_packet_t pcfg_rdrq_packet_e2w_esti;
rdrq_packet_t pcfg_rdrq_packet_e2w_wsto;
rdrq_packet_t pcfg_rdrq_packet_w2e_esto;
rdrq_packet_t pcfg_rdrq_packet_w2e_wsti;
rdrs_packet_t pcfg_rdrs_packet_e2w_esti;
rdrs_packet_t pcfg_rdrs_packet_e2w_wsto;
rdrs_packet_t pcfg_rdrs_packet_w2e_esto;
rdrs_packet_t pcfg_rdrs_packet_w2e_wsti;
rdrq_packet_t rdrq_packet_dma2bank;
rdrq_packet_t rdrq_packet_dma2ring;
rdrq_packet_t rdrq_packet_pcfgdma2bank;
rdrq_packet_t rdrq_packet_pcfgdma2ring;
rdrq_packet_t rdrq_packet_pcfgring2bank;
rdrq_packet_t rdrq_packet_procsw2bank;
rdrq_packet_t rdrq_packet_ring2bank;
rdrq_bank_packet_t [1:0] rdrq_packet_sw2bankarr;
rdrs_packet_t rdrs_packet_bank2dma;
rdrs_packet_t rdrs_packet_bank2pcfgdma;
rdrs_packet_t rdrs_packet_bank2pcfgring;
rdrs_packet_t rdrs_packet_bank2procsw;
rdrs_packet_t rdrs_packet_bank2ring;
rdrs_packet_t [1:0] rdrs_packet_bankarr2sw;
rdrs_packet_t rdrs_packet_pcfgring2dma;
rdrs_packet_t rdrs_packet_ring2dma;
rdrq_packet_t strm_rdrq_packet_e2w_esti;
rdrq_packet_t strm_rdrq_packet_e2w_wsto;
rdrq_packet_t strm_rdrq_packet_w2e_esto;
rdrq_packet_t strm_rdrq_packet_w2e_wsti;
rdrs_packet_t strm_rdrs_packet_e2w_esti;
rdrs_packet_t strm_rdrs_packet_e2w_wsto;
rdrs_packet_t strm_rdrs_packet_w2e_esto;
rdrs_packet_t strm_rdrs_packet_w2e_wsti;
wr_packet_t strm_wr_packet_e2w_esti;
wr_packet_t strm_wr_packet_e2w_wsto;
wr_packet_t strm_wr_packet_w2e_esto;
wr_packet_t strm_wr_packet_w2e_wsti;
wr_packet_t wr_packet_dma2bank;
wr_packet_t wr_packet_dma2ring;
wr_packet_t wr_packet_procsw2bank;
wr_packet_t wr_packet_ring2bank;
wr_bank_packet_t [1:0] wr_packet_sw2bankarr;
glb_tile_ifc_A_12_D_32 if_cfg_est_m();
glb_tile_ifc_A_12_D_32 if_cfg_wst_s();
glb_tile_ifc_A_19_D_64 if_proc_est_m();
glb_tile_ifc_A_19_D_64 if_proc_wst_s();
assign if_proc_est_m_wr_en = if_proc_est_m.wr_en;
assign if_proc_wst_s.wr_en = if_proc_wst_s_wr_en;
assign if_proc_est_m_wr_addr = if_proc_est_m.wr_addr;
assign if_proc_wst_s.wr_addr = if_proc_wst_s_wr_addr;
assign if_proc_est_m_wr_data = if_proc_est_m.wr_data;
assign if_proc_wst_s.wr_data = if_proc_wst_s_wr_data;
assign if_proc_est_m_rd_en = if_proc_est_m.rd_en;
assign if_proc_wst_s.rd_en = if_proc_wst_s_rd_en;
assign if_proc_est_m_rd_addr = if_proc_est_m.rd_addr;
assign if_proc_wst_s.rd_addr = if_proc_wst_s_rd_addr;
assign if_proc_est_m_wr_strb = if_proc_est_m.wr_strb;
assign if_proc_wst_s.wr_strb = if_proc_wst_s_wr_strb;
assign if_proc_est_m_wr_clk_en = if_proc_est_m.wr_clk_en;
assign if_proc_wst_s.wr_clk_en = if_proc_wst_s_wr_clk_en;
assign if_proc_est_m_rd_clk_en = if_proc_est_m.rd_clk_en;
assign if_proc_wst_s.rd_clk_en = if_proc_wst_s_rd_clk_en;
assign if_proc_est_m.rd_data = if_proc_est_m_rd_data;
assign if_proc_wst_s_rd_data = if_proc_wst_s.rd_data;
assign if_proc_est_m.rd_data_valid = if_proc_est_m_rd_data_valid;
assign if_proc_wst_s_rd_data_valid = if_proc_wst_s.rd_data_valid;
assign if_cfg_est_m_wr_en = if_cfg_est_m.wr_en;
assign if_cfg_wst_s.wr_en = if_cfg_wst_s_wr_en;
assign if_cfg_est_m_wr_addr = if_cfg_est_m.wr_addr;
assign if_cfg_wst_s.wr_addr = if_cfg_wst_s_wr_addr;
assign if_cfg_est_m_wr_data = if_cfg_est_m.wr_data;
assign if_cfg_wst_s.wr_data = if_cfg_wst_s_wr_data;
assign if_cfg_est_m_rd_en = if_cfg_est_m.rd_en;
assign if_cfg_wst_s.rd_en = if_cfg_wst_s_rd_en;
assign if_cfg_est_m_rd_addr = if_cfg_est_m.rd_addr;
assign if_cfg_wst_s.rd_addr = if_cfg_wst_s_rd_addr;
assign if_cfg_est_m_wr_clk_en = if_cfg_est_m.wr_clk_en;
assign if_cfg_wst_s.wr_clk_en = if_cfg_wst_s_wr_clk_en;
assign if_cfg_est_m_rd_clk_en = if_cfg_est_m.rd_clk_en;
assign if_cfg_wst_s.rd_clk_en = if_cfg_wst_s_rd_clk_en;
assign if_cfg_est_m.rd_data = if_cfg_est_m_rd_data;
assign if_cfg_wst_s_rd_data = if_cfg_wst_s.rd_data;
assign if_cfg_est_m.rd_data_valid = if_cfg_est_m_rd_data_valid;
assign if_cfg_wst_s_rd_data_valid = if_cfg_wst_s.rd_data_valid;
assign strm_wr_packet_w2e_wsti.wr_en = strm_wr_en_w2e_wsti;
assign strm_wr_packet_w2e_wsti.wr_strb = strm_wr_strb_w2e_wsti;
assign strm_wr_packet_w2e_wsti.wr_addr = strm_wr_addr_w2e_wsti;
assign strm_wr_packet_w2e_wsti.wr_data = strm_wr_data_w2e_wsti;
assign strm_wr_en_w2e_esto = strm_wr_packet_w2e_esto.wr_en;
assign strm_wr_strb_w2e_esto = strm_wr_packet_w2e_esto.wr_strb;
assign strm_wr_addr_w2e_esto = strm_wr_packet_w2e_esto.wr_addr;
assign strm_wr_data_w2e_esto = strm_wr_packet_w2e_esto.wr_data;
assign strm_wr_packet_e2w_esti.wr_en = strm_wr_en_e2w_esti;
assign strm_wr_packet_e2w_esti.wr_strb = strm_wr_strb_e2w_esti;
assign strm_wr_packet_e2w_esti.wr_addr = strm_wr_addr_e2w_esti;
assign strm_wr_packet_e2w_esti.wr_data = strm_wr_data_e2w_esti;
assign strm_wr_en_e2w_wsto = strm_wr_packet_e2w_wsto.wr_en;
assign strm_wr_strb_e2w_wsto = strm_wr_packet_e2w_wsto.wr_strb;
assign strm_wr_addr_e2w_wsto = strm_wr_packet_e2w_wsto.wr_addr;
assign strm_wr_data_e2w_wsto = strm_wr_packet_e2w_wsto.wr_data;
assign strm_rdrq_packet_w2e_wsti.rd_en = strm_rd_en_w2e_wsti;
assign strm_rdrq_packet_w2e_wsti.rd_addr = strm_rd_addr_w2e_wsti;
assign strm_rd_en_w2e_esto = strm_rdrq_packet_w2e_esto.rd_en;
assign strm_rd_addr_w2e_esto = strm_rdrq_packet_w2e_esto.rd_addr;
assign strm_rdrq_packet_e2w_esti.rd_en = strm_rd_en_e2w_esti;
assign strm_rdrq_packet_e2w_esti.rd_addr = strm_rd_addr_e2w_esti;
assign strm_rd_en_e2w_wsto = strm_rdrq_packet_e2w_wsto.rd_en;
assign strm_rd_addr_e2w_wsto = strm_rdrq_packet_e2w_wsto.rd_addr;
assign strm_rd_data_e2w_wsto = strm_rdrs_packet_e2w_wsto.rd_data;
assign strm_rd_data_valid_e2w_wsto = strm_rdrs_packet_e2w_wsto.rd_data_valid;
assign strm_rdrs_packet_e2w_esti.rd_data = strm_rd_data_e2w_esti;
assign strm_rdrs_packet_e2w_esti.rd_data_valid = strm_rd_data_valid_e2w_esti;
assign strm_rdrs_packet_w2e_wsti.rd_data = strm_rd_data_w2e_wsti;
assign strm_rdrs_packet_w2e_wsti.rd_data_valid = strm_rd_data_valid_w2e_wsti;
assign strm_rd_data_w2e_esto = strm_rdrs_packet_w2e_esto.rd_data;
assign strm_rd_data_valid_w2e_esto = strm_rdrs_packet_w2e_esto.rd_data_valid;
assign pcfg_rdrq_packet_w2e_wsti.rd_en = pcfg_rd_en_w2e_wsti;
assign pcfg_rdrq_packet_w2e_wsti.rd_addr = pcfg_rd_addr_w2e_wsti;
assign pcfg_rd_en_w2e_esto = pcfg_rdrq_packet_w2e_esto.rd_en;
assign pcfg_rd_addr_w2e_esto = pcfg_rdrq_packet_w2e_esto.rd_addr;
assign pcfg_rdrq_packet_e2w_esti.rd_en = pcfg_rd_en_e2w_esti;
assign pcfg_rdrq_packet_e2w_esti.rd_addr = pcfg_rd_addr_e2w_esti;
assign pcfg_rd_en_e2w_wsto = pcfg_rdrq_packet_e2w_wsto.rd_en;
assign pcfg_rd_addr_e2w_wsto = pcfg_rdrq_packet_e2w_wsto.rd_addr;
assign pcfg_rd_data_e2w_wsto = pcfg_rdrs_packet_e2w_wsto.rd_data;
assign pcfg_rd_data_valid_e2w_wsto = pcfg_rdrs_packet_e2w_wsto.rd_data_valid;
assign pcfg_rdrs_packet_e2w_esti.rd_data = pcfg_rd_data_e2w_esti;
assign pcfg_rdrs_packet_e2w_esti.rd_data_valid = pcfg_rd_data_valid_e2w_esti;
assign pcfg_rdrs_packet_w2e_wsti.rd_data = pcfg_rd_data_w2e_wsti;
assign pcfg_rdrs_packet_w2e_wsti.rd_data_valid = pcfg_rd_data_valid_w2e_wsti;
assign pcfg_rd_data_w2e_esto = pcfg_rdrs_packet_w2e_esto.rd_data;
assign pcfg_rd_data_valid_w2e_esto = pcfg_rdrs_packet_w2e_esto.rd_data_valid;
assign clk_en_cfg = if_cfg_wst_s.wr_clk_en | if_cfg_wst_s.rd_clk_en;
assign glb_clk_gate_cfg_enable = clk_en_cfg | clk_en_master;
assign glb_clk_gate_pcfg_broadcast_enable = clk_en_pcfg_broadcast | clk_en_master;
assign clk_en_ld_dma = cfg_ld_dma_ctrl.mode != 2'h0;
assign glb_clk_gate_ld_dma_enable = clk_en_ld_dma | clk_en_master;
assign clk_en_st_dma = cfg_st_dma_ctrl.mode != 2'h0;
assign glb_clk_gate_st_dma_enable = clk_en_st_dma | clk_en_master;
assign clk_en_proc_switch = if_proc_wst_s.wr_clk_en | if_proc_wst_s.rd_clk_en;
assign glb_clk_gate_proc_switch_enable = clk_en_proc_switch | clk_en_master;
assign clk_en_pcfg_dma = cfg_pcfg_dma_ctrl.mode != 1'h0;
assign glb_clk_gate_pcfg_dma_enable = clk_en_pcfg_dma | clk_en_master;
assign clk_en_strm_switch = cfg_tile_connected_next | cfg_tile_connected_prev;
assign glb_clk_gate_strm_switch_enable = clk_en_strm_switch | clk_en_master;
assign clk_en_pcfg_switch = cfg_pcfg_tile_connected_next | cfg_pcfg_tile_connected_prev;
assign glb_clk_gate_pcfg_switch_enable = clk_en_pcfg_switch | clk_en_master;
assign clk_en_bank = clk_en_lddma2bank | clk_en_stdma2bank | clk_en_pcfgdma2bank | clk_en_ring2bank |
    clk_en_pcfgring2bank | clk_en_procsw2bank;
assign glb_clk_gate_bank_enable = clk_en_bank | clk_en_master | clk_en_bank_master;
assign glb_cfg_gclk = gclk_cfg;
assign cfg_tile_connected_next = glb_cfg_cfg_data_network.tile_connected;
assign cfg_tile_connected_prev = cfg_tile_connected_wsti;
assign cfg_tile_connected_esto = cfg_tile_connected_next;
assign cfg_pcfg_tile_connected_next = glb_cfg_cfg_pcfg_network.tile_connected;
assign cfg_pcfg_tile_connected_prev = cfg_pcfg_tile_connected_wsti;
assign cfg_pcfg_tile_connected_esto = cfg_pcfg_tile_connected_next;
assign glb_pcfg_broadcast_clk = gclk_pcfg_broadcast;
assign glb_store_dma_clk = gclk_st_dma;
assign glb_load_dma_clk = gclk_ld_dma;
assign glb_pcfg_dma_clk = gclk_pcfg_dma;
assign glb_bank_mux_clk = gclk_bank;
assign glb_proc_switch_gclk = gclk_proc_switch;
assign glb_strm_ring_switch_clk = gclk_strm_switch;
assign glb_strm_ring_switch_cfg_ld_dma_on = cfg_ld_dma_ctrl.mode != 2'h0;
assign glb_pcfg_ring_switch_clk = gclk_pcfg_switch;
assign glb_pcfg_ring_switch_cfg_ld_dma_on = cfg_pcfg_dma_ctrl.mode != 1'h0;
assign glb_bank_0_clk = gclk_bank;
assign rdrs_packet_bankarr2sw[0] = glb_bank_0_rdrs_packet;
assign glb_bank_1_clk = gclk_bank;
assign rdrs_packet_bankarr2sw[1] = glb_bank_1_rdrs_packet;
assign cgra_cfg_g2f_cfg_wr_en[0] = cgra_cfg_g2f_cfg_w[0].wr_en;
assign cgra_cfg_g2f_cfg_rd_en[0] = cgra_cfg_g2f_cfg_w[0].rd_en;
assign cgra_cfg_g2f_cfg_addr[0] = cgra_cfg_g2f_cfg_w[0].addr;
assign cgra_cfg_g2f_cfg_data[0] = cgra_cfg_g2f_cfg_w[0].data;
assign cgra_cfg_g2f_cfg_wr_en[1] = cgra_cfg_g2f_cfg_w[1].wr_en;
assign cgra_cfg_g2f_cfg_rd_en[1] = cgra_cfg_g2f_cfg_w[1].rd_en;
assign cgra_cfg_g2f_cfg_addr[1] = cgra_cfg_g2f_cfg_w[1].addr;
assign cgra_cfg_g2f_cfg_data[1] = cgra_cfg_g2f_cfg_w[1].data;
assign glb_pcfg_broadcast_cgra_cfg_jtag_wsti.wr_en = cgra_cfg_jtag_wr_en_wsti;
assign glb_pcfg_broadcast_cgra_cfg_jtag_wsti.rd_en = cgra_cfg_jtag_rd_en_wsti;
assign glb_pcfg_broadcast_cgra_cfg_jtag_wsti.addr = cgra_cfg_jtag_addr_wsti;
assign glb_pcfg_broadcast_cgra_cfg_jtag_wsti.data = cgra_cfg_jtag_data_wsti;
assign cgra_cfg_jtag_wr_en_esto = glb_pcfg_broadcast_cgra_cfg_jtag_esto.wr_en;
assign cgra_cfg_jtag_rd_en_esto = glb_pcfg_broadcast_cgra_cfg_jtag_esto.rd_en;
assign cgra_cfg_jtag_addr_esto = glb_pcfg_broadcast_cgra_cfg_jtag_esto.addr;
assign cgra_cfg_jtag_data_esto = glb_pcfg_broadcast_cgra_cfg_jtag_esto.data;
assign glb_pcfg_broadcast_cgra_cfg_pcfg_wsti.wr_en = cgra_cfg_pcfg_wr_en_w2e_wsti;
assign glb_pcfg_broadcast_cgra_cfg_pcfg_wsti.rd_en = cgra_cfg_pcfg_rd_en_w2e_wsti;
assign glb_pcfg_broadcast_cgra_cfg_pcfg_wsti.addr = cgra_cfg_pcfg_addr_w2e_wsti;
assign glb_pcfg_broadcast_cgra_cfg_pcfg_wsti.data = cgra_cfg_pcfg_data_w2e_wsti;
assign cgra_cfg_pcfg_wr_en_w2e_esto = glb_pcfg_broadcast_cgra_cfg_pcfg_esto.wr_en;
assign cgra_cfg_pcfg_rd_en_w2e_esto = glb_pcfg_broadcast_cgra_cfg_pcfg_esto.rd_en;
assign cgra_cfg_pcfg_addr_w2e_esto = glb_pcfg_broadcast_cgra_cfg_pcfg_esto.addr;
assign cgra_cfg_pcfg_data_w2e_esto = glb_pcfg_broadcast_cgra_cfg_pcfg_esto.data;
assign glb_pcfg_broadcast_cgra_cfg_pcfg_esti.wr_en = cgra_cfg_pcfg_wr_en_e2w_esti;
assign glb_pcfg_broadcast_cgra_cfg_pcfg_esti.rd_en = cgra_cfg_pcfg_rd_en_e2w_esti;
assign glb_pcfg_broadcast_cgra_cfg_pcfg_esti.addr = cgra_cfg_pcfg_addr_e2w_esti;
assign glb_pcfg_broadcast_cgra_cfg_pcfg_esti.data = cgra_cfg_pcfg_data_e2w_esti;
assign cgra_cfg_pcfg_wr_en_e2w_wsto = glb_pcfg_broadcast_cgra_cfg_pcfg_wsto.wr_en;
assign cgra_cfg_pcfg_rd_en_e2w_wsto = glb_pcfg_broadcast_cgra_cfg_pcfg_wsto.rd_en;
assign cgra_cfg_pcfg_addr_e2w_wsto = glb_pcfg_broadcast_cgra_cfg_pcfg_wsto.addr;
assign cgra_cfg_pcfg_data_e2w_wsto = glb_pcfg_broadcast_cgra_cfg_pcfg_wsto.data;
clk_gate glb_clk_gate_cfg (
  .clk(clk),
  .enable(glb_clk_gate_cfg_enable),
  .gclk(gclk_cfg)
);

clk_gate glb_clk_gate_pcfg_broadcast (
  .clk(clk),
  .enable(glb_clk_gate_pcfg_broadcast_enable),
  .gclk(gclk_pcfg_broadcast)
);

clk_gate glb_clk_gate_ld_dma (
  .clk(clk),
  .enable(glb_clk_gate_ld_dma_enable),
  .gclk(gclk_ld_dma)
);

clk_gate glb_clk_gate_st_dma (
  .clk(clk),
  .enable(glb_clk_gate_st_dma_enable),
  .gclk(gclk_st_dma)
);

clk_gate glb_clk_gate_proc_switch (
  .clk(clk),
  .enable(glb_clk_gate_proc_switch_enable),
  .gclk(gclk_proc_switch)
);

clk_gate glb_clk_gate_pcfg_dma (
  .clk(clk),
  .enable(glb_clk_gate_pcfg_dma_enable),
  .gclk(gclk_pcfg_dma)
);

clk_gate glb_clk_gate_strm_switch (
  .clk(clk),
  .enable(glb_clk_gate_strm_switch_enable),
  .gclk(gclk_strm_switch)
);

clk_gate glb_clk_gate_pcfg_switch (
  .clk(clk),
  .enable(glb_clk_gate_pcfg_switch_enable),
  .gclk(gclk_pcfg_switch)
);

clk_gate glb_clk_gate_bank (
  .clk(clk),
  .enable(glb_clk_gate_bank_enable),
  .gclk(gclk_bank)
);

glb_cfg glb_cfg (
  .gclk(glb_cfg_gclk),
  .glb_tile_id(glb_tile_id),
  .mclk(clk),
  .if_cfg_wst_s(if_cfg_wst_s.slave),
  .if_cfg_est_m(if_cfg_est_m.master),
  .reset(reset),
  .cfg_data_network(glb_cfg_cfg_data_network),
  .cfg_ld_dma_ctrl(cfg_ld_dma_ctrl),
  .cfg_ld_dma_header(cfg_ld_dma_header),
  .cfg_pcfg_broadcast_mux(cfg_pcfg_broadcast_mux),
  .cfg_pcfg_dma_ctrl(cfg_pcfg_dma_ctrl),
  .cfg_pcfg_dma_header(cfg_pcfg_dma_header),
  .cfg_pcfg_network(glb_cfg_cfg_pcfg_network),
  .cfg_st_dma_ctrl(cfg_st_dma_ctrl),
  .cfg_st_dma_header(cfg_st_dma_header)
);

glb_pcfg_broadcast glb_pcfg_broadcast (
  .cfg_pcfg_broadcast_mux(cfg_pcfg_broadcast_mux),
  .cgra_cfg_dma2mux(cgra_cfg_pcfgdma2mux),
  .cgra_cfg_jtag_addr_bypass_wsti(cgra_cfg_jtag_addr_bypass_wsti),
  .cgra_cfg_jtag_rd_en_bypass_wsti(cgra_cfg_jtag_rd_en_bypass_wsti),
  .cgra_cfg_jtag_wsti(glb_pcfg_broadcast_cgra_cfg_jtag_wsti),
  .cgra_cfg_pcfg_esti(glb_pcfg_broadcast_cgra_cfg_pcfg_esti),
  .cgra_cfg_pcfg_wsti(glb_pcfg_broadcast_cgra_cfg_pcfg_wsti),
  .clk(glb_pcfg_broadcast_clk),
  .reset(reset),
  .cgra_cfg_g2f(cgra_cfg_g2f_cfg_w),
  .cgra_cfg_jtag_addr_bypass_esto(cgra_cfg_jtag_addr_bypass_esto),
  .cgra_cfg_jtag_esto(glb_pcfg_broadcast_cgra_cfg_jtag_esto),
  .cgra_cfg_jtag_rd_en_bypass_esto(cgra_cfg_jtag_rd_en_bypass_esto),
  .cgra_cfg_pcfg_esto(glb_pcfg_broadcast_cgra_cfg_pcfg_esto),
  .cgra_cfg_pcfg_wsto(glb_pcfg_broadcast_cgra_cfg_pcfg_wsto)
);

glb_store_dma glb_store_dma (
  .cfg_data_network_f2g_mux(cfg_st_dma_ctrl.data_mux),
  .cfg_data_network_latency(glb_cfg_cfg_data_network.latency),
  .cfg_st_dma_ctrl_mode(cfg_st_dma_ctrl.mode),
  .cfg_st_dma_ctrl_use_valid(cfg_st_dma_ctrl.use_valid),
  .cfg_st_dma_header(cfg_st_dma_header),
  .cfg_st_dma_num_repeat(cfg_st_dma_ctrl.num_repeat),
  .cfg_tile_connected_next(cfg_tile_connected_next),
  .cfg_tile_connected_prev(cfg_tile_connected_prev),
  .clk(glb_store_dma_clk),
  .data_f2g(strm_data_f2g),
  .data_valid_f2g(strm_data_valid_f2g),
  .reset(reset),
  .st_dma_start_pulse(strm_f2g_start_pulse),
  .clk_en_dma2bank(clk_en_stdma2bank),
  .st_dma_done_interrupt(strm_f2g_interrupt_pulse),
  .wr_packet_dma2bank(wr_packet_dma2bank),
  .wr_packet_dma2ring(wr_packet_dma2ring)
);

glb_load_dma glb_load_dma (
  .cfg_data_network_g2f_mux(cfg_ld_dma_ctrl.data_mux),
  .cfg_data_network_latency(glb_cfg_cfg_data_network.latency),
  .cfg_ld_dma_ctrl_mode(cfg_ld_dma_ctrl.mode),
  .cfg_ld_dma_ctrl_use_flush(cfg_ld_dma_ctrl.use_flush),
  .cfg_ld_dma_ctrl_use_valid(cfg_ld_dma_ctrl.use_valid),
  .cfg_ld_dma_header(cfg_ld_dma_header),
  .cfg_ld_dma_num_repeat(cfg_ld_dma_ctrl.num_repeat),
  .cfg_tile_connected_next(cfg_tile_connected_next),
  .cfg_tile_connected_prev(cfg_tile_connected_prev),
  .clk(glb_load_dma_clk),
  .glb_tile_id(glb_tile_id),
  .ld_dma_start_pulse(strm_g2f_start_pulse),
  .rdrs_packet_bank2dma(rdrs_packet_bank2dma),
  .rdrs_packet_ring2dma(rdrs_packet_ring2dma),
  .reset(reset),
  .clk_en_dma2bank(clk_en_lddma2bank),
  .data_flush(data_flush),
  .data_g2f(strm_data_g2f),
  .data_valid_g2f(strm_data_valid_g2f),
  .ld_dma_done_interrupt(strm_g2f_interrupt_pulse),
  .rdrq_packet_dma2bank(rdrq_packet_dma2bank),
  .rdrq_packet_dma2ring(rdrq_packet_dma2ring)
);

glb_pcfg_dma glb_pcfg_dma (
  .cfg_pcfg_dma_ctrl_mode(cfg_pcfg_dma_ctrl.mode),
  .cfg_pcfg_dma_ctrl_relocation_is_msb(cfg_pcfg_dma_ctrl.relocation_is_msb),
  .cfg_pcfg_dma_ctrl_relocation_value(cfg_pcfg_dma_ctrl.relocation_value),
  .cfg_pcfg_dma_header(cfg_pcfg_dma_header),
  .cfg_pcfg_network_latency(glb_cfg_cfg_pcfg_network.latency),
  .cfg_pcfg_tile_connected_next(cfg_pcfg_tile_connected_next),
  .cfg_pcfg_tile_connected_prev(cfg_pcfg_tile_connected_prev),
  .clk(glb_pcfg_dma_clk),
  .glb_tile_id(glb_tile_id),
  .pcfg_dma_start_pulse(pcfg_start_pulse),
  .rdrs_packet_bank2dma(rdrs_packet_bank2pcfgdma),
  .rdrs_packet_ring2dma(rdrs_packet_pcfgring2dma),
  .reset(reset),
  .cgra_cfg_pcfg(cgra_cfg_pcfgdma2mux),
  .clk_en_dma2bank(clk_en_pcfgdma2bank),
  .pcfg_dma_done_interrupt(pcfg_g2f_interrupt_pulse),
  .rdrq_packet_dma2bank(rdrq_packet_pcfgdma2bank),
  .rdrq_packet_dma2ring(rdrq_packet_pcfgdma2ring)
);

glb_bank_mux glb_bank_mux (
  .cfg_pcfg_tile_connected_next(cfg_pcfg_tile_connected_next),
  .cfg_pcfg_tile_connected_prev(cfg_pcfg_tile_connected_prev),
  .cfg_tile_connected_next(cfg_tile_connected_next),
  .cfg_tile_connected_prev(cfg_tile_connected_prev),
  .clk(glb_bank_mux_clk),
  .glb_tile_id(glb_tile_id),
  .rdrq_packet_dma2bank(rdrq_packet_dma2bank),
  .rdrq_packet_pcfgdma2bank(rdrq_packet_pcfgdma2bank),
  .rdrq_packet_pcfgring2bank(rdrq_packet_pcfgring2bank),
  .rdrq_packet_procsw2bank(rdrq_packet_procsw2bank),
  .rdrq_packet_ring2bank(rdrq_packet_ring2bank),
  .rdrs_packet_bankarr2sw(rdrs_packet_bankarr2sw),
  .reset(reset),
  .wr_packet_dma2bank(wr_packet_dma2bank),
  .wr_packet_procsw2bank(wr_packet_procsw2bank),
  .wr_packet_ring2bank(wr_packet_ring2bank),
  .rdrq_packet_sw2bankarr(rdrq_packet_sw2bankarr),
  .rdrs_packet_bank2dma(rdrs_packet_bank2dma),
  .rdrs_packet_bank2pcfgdma(rdrs_packet_bank2pcfgdma),
  .rdrs_packet_bank2pcfgring(rdrs_packet_bank2pcfgring),
  .rdrs_packet_bank2procsw(rdrs_packet_bank2procsw),
  .rdrs_packet_bank2ring(rdrs_packet_bank2ring),
  .wr_packet_sw2bankarr(wr_packet_sw2bankarr)
);

glb_switch glb_proc_switch (
  .gclk(glb_proc_switch_gclk),
  .glb_tile_id(glb_tile_id),
  .mclk(clk),
  .if_wst_s(if_proc_wst_s.slave),
  .if_est_m(if_proc_est_m.master),
  .rdrs_packet(rdrs_packet_bank2procsw),
  .reset(reset),
  .clk_en_sw2bank(clk_en_procsw2bank),
  .rdrq_packet(rdrq_packet_procsw2bank),
  .wr_packet(wr_packet_procsw2bank)
);

glb_ring_switch_WR_RD glb_strm_ring_switch (
  .cfg_ld_dma_on(glb_strm_ring_switch_cfg_ld_dma_on),
  .cfg_tile_connected_next(cfg_tile_connected_next),
  .cfg_tile_connected_prev(cfg_tile_connected_prev),
  .clk(glb_strm_ring_switch_clk),
  .glb_tile_id(glb_tile_id),
  .rdrq_packet_dma2ring(rdrq_packet_dma2ring),
  .rdrq_packet_e2w_esti(strm_rdrq_packet_e2w_esti),
  .rdrq_packet_w2e_wsti(strm_rdrq_packet_w2e_wsti),
  .rdrs_packet_bank2ring(rdrs_packet_bank2ring),
  .rdrs_packet_e2w_esti(strm_rdrs_packet_e2w_esti),
  .rdrs_packet_w2e_wsti(strm_rdrs_packet_w2e_wsti),
  .reset(reset),
  .wr_packet_dma2ring(wr_packet_dma2ring),
  .wr_packet_e2w_esti(strm_wr_packet_e2w_esti),
  .wr_packet_w2e_wsti(strm_wr_packet_w2e_wsti),
  .clk_en_ring2bank(clk_en_ring2bank),
  .rdrq_packet_e2w_wsto(strm_rdrq_packet_e2w_wsto),
  .rdrq_packet_ring2bank(rdrq_packet_ring2bank),
  .rdrq_packet_w2e_esto(strm_rdrq_packet_w2e_esto),
  .rdrs_packet_e2w_wsto(strm_rdrs_packet_e2w_wsto),
  .rdrs_packet_ring2dma(rdrs_packet_ring2dma),
  .rdrs_packet_w2e_esto(strm_rdrs_packet_w2e_esto),
  .wr_packet_e2w_wsto(strm_wr_packet_e2w_wsto),
  .wr_packet_ring2bank(wr_packet_ring2bank),
  .wr_packet_w2e_esto(strm_wr_packet_w2e_esto)
);

glb_ring_switch_RD glb_pcfg_ring_switch (
  .cfg_ld_dma_on(glb_pcfg_ring_switch_cfg_ld_dma_on),
  .cfg_tile_connected_next(cfg_pcfg_tile_connected_next),
  .cfg_tile_connected_prev(cfg_pcfg_tile_connected_prev),
  .clk(glb_pcfg_ring_switch_clk),
  .glb_tile_id(glb_tile_id),
  .rdrq_packet_dma2ring(rdrq_packet_pcfgdma2ring),
  .rdrq_packet_e2w_esti(pcfg_rdrq_packet_e2w_esti),
  .rdrq_packet_w2e_wsti(pcfg_rdrq_packet_w2e_wsti),
  .rdrs_packet_bank2ring(rdrs_packet_bank2pcfgring),
  .rdrs_packet_e2w_esti(pcfg_rdrs_packet_e2w_esti),
  .rdrs_packet_w2e_wsti(pcfg_rdrs_packet_w2e_wsti),
  .reset(reset),
  .clk_en_ring2bank(clk_en_pcfgring2bank),
  .rdrq_packet_e2w_wsto(pcfg_rdrq_packet_e2w_wsto),
  .rdrq_packet_ring2bank(rdrq_packet_pcfgring2bank),
  .rdrq_packet_w2e_esto(pcfg_rdrq_packet_w2e_esto),
  .rdrs_packet_e2w_wsto(pcfg_rdrs_packet_e2w_wsto),
  .rdrs_packet_ring2dma(rdrs_packet_pcfgring2dma),
  .rdrs_packet_w2e_esto(pcfg_rdrs_packet_w2e_esto)
);

glb_bank glb_bank_0 (
  .clk(glb_bank_0_clk),
  .rdrq_packet(rdrq_packet_sw2bankarr[0]),
  .reset(reset),
  .wr_packet(wr_packet_sw2bankarr[0]),
  .rdrs_packet(glb_bank_0_rdrs_packet)
);

glb_bank glb_bank_1 (
  .clk(glb_bank_1_clk),
  .rdrq_packet(rdrq_packet_sw2bankarr[1]),
  .reset(reset),
  .wr_packet(wr_packet_sw2bankarr[1]),
  .rdrs_packet(glb_bank_1_rdrs_packet)
);

endmodule   // glb_tile

module global_buffer (
  input logic [31:0] cgra_cfg_jtag_gc2glb_addr,
  input logic [31:0] cgra_cfg_jtag_gc2glb_data,
  input logic cgra_cfg_jtag_gc2glb_rd_en,
  input logic cgra_cfg_jtag_gc2glb_wr_en,
  input logic [3:0] cgra_stall_in,
  input logic clk,
  input logic flush_crossbar_sel,
  input logic [1:0] glb_clk_en_bank_master,
  input logic [1:0] glb_clk_en_master,
  input logic [11:0] if_cfg_rd_addr,
  input logic if_cfg_rd_clk_en,
  input logic if_cfg_rd_en,
  input logic [11:0] if_cfg_wr_addr,
  input logic if_cfg_wr_clk_en,
  input logic [31:0] if_cfg_wr_data,
  input logic if_cfg_wr_en,
  input logic [18:0] if_sram_cfg_rd_addr,
  input logic if_sram_cfg_rd_en,
  input logic [18:0] if_sram_cfg_wr_addr,
  input logic [31:0] if_sram_cfg_wr_data,
  input logic if_sram_cfg_wr_en,
  input logic [1:0] pcfg_broadcast_stall,
  input logic [1:0] pcfg_start_pulse,
  input logic [18:0] proc_rd_addr,
  input logic proc_rd_en,
  input logic [18:0] proc_wr_addr,
  input logic [63:0] proc_wr_data,
  input logic proc_wr_en,
  input logic [7:0] proc_wr_strb,
  input logic reset,
  input logic [1:0][1:0] [15:0] strm_data_f2g,
  input logic [1:0][1:0] strm_data_valid_f2g,
  input logic [1:0] strm_f2g_start_pulse,
  input logic [1:0] strm_g2f_start_pulse,
  output logic [1:0][1:0] [31:0] cgra_cfg_g2f_cfg_addr,
  output logic [1:0][1:0] [31:0] cgra_cfg_g2f_cfg_data,
  output logic [1:0][1:0] cgra_cfg_g2f_cfg_rd_en,
  output logic [1:0][1:0] cgra_cfg_g2f_cfg_wr_en,
  output logic [3:0] cgra_stall,
  output logic [31:0] if_cfg_rd_data,
  output logic if_cfg_rd_data_valid,
  output logic [31:0] if_sram_cfg_rd_data,
  output logic if_sram_cfg_rd_data_valid,
  output logic [1:0] pcfg_g2f_interrupt_pulse,
  output logic [63:0] proc_rd_data,
  output logic proc_rd_data_valid,
  output logic strm_data_flush_g2f,
  output logic [1:0][1:0] [15:0] strm_data_g2f,
  output logic [1:0][1:0] strm_data_valid_g2f,
  output logic [1:0] strm_f2g_interrupt_pulse,
  output logic [1:0] strm_g2f_interrupt_pulse
);

typedef enum logic {
  axi = 1'h0,
  jtag = 1'h1
} proc_rd_type_e;
logic [2:0] cfg_pcfg_tile_connected;
logic [2:0] cfg_tile_connected;
logic [1:0][31:0] cgra_cfg_jtag_addr_bypass_esto;
logic [1:0][31:0] cgra_cfg_jtag_addr_bypass_wsti;
logic [1:0][31:0] cgra_cfg_jtag_addr_esto;
logic [1:0][31:0] cgra_cfg_jtag_addr_wsti;
logic [1:0][31:0] cgra_cfg_jtag_data_esto;
logic [1:0][31:0] cgra_cfg_jtag_data_wsti;
logic [31:0] cgra_cfg_jtag_gc2glb_addr_d;
logic [31:0] cgra_cfg_jtag_gc2glb_data_d;
logic cgra_cfg_jtag_gc2glb_rd_en_d;
logic cgra_cfg_jtag_gc2glb_wr_en_d;
logic [1:0] cgra_cfg_jtag_rd_en_bypass_esto;
logic [1:0] cgra_cfg_jtag_rd_en_bypass_wsti;
logic [1:0] cgra_cfg_jtag_rd_en_esto;
logic [1:0] cgra_cfg_jtag_rd_en_wsti;
logic [1:0] cgra_cfg_jtag_wr_en_esto;
logic [1:0] cgra_cfg_jtag_wr_en_wsti;
logic [1:0][31:0] cgra_cfg_pcfg_addr_esti;
logic [1:0][31:0] cgra_cfg_pcfg_addr_esto;
logic [1:0][31:0] cgra_cfg_pcfg_addr_wsti;
logic [1:0][31:0] cgra_cfg_pcfg_addr_wsto;
logic [1:0][31:0] cgra_cfg_pcfg_data_esti;
logic [1:0][31:0] cgra_cfg_pcfg_data_esto;
logic [1:0][31:0] cgra_cfg_pcfg_data_wsti;
logic [1:0][31:0] cgra_cfg_pcfg_data_wsto;
logic [1:0] cgra_cfg_pcfg_rd_en_esti;
logic [1:0] cgra_cfg_pcfg_rd_en_esto;
logic [1:0] cgra_cfg_pcfg_rd_en_wsti;
logic [1:0] cgra_cfg_pcfg_rd_en_wsto;
logic [1:0] cgra_cfg_pcfg_wr_en_esti;
logic [1:0] cgra_cfg_pcfg_wr_en_esto;
logic [1:0] cgra_cfg_pcfg_wr_en_wsti;
logic [1:0] cgra_cfg_pcfg_wr_en_wsto;
logic [1:0] data_flush;
logic [1:0] data_flush_d;
logic [1:0] flush_crossbar_in;
logic flush_crossbar_sel_w;
logic glb_tile_gen_0_cfg_pcfg_tile_connected_esto;
logic glb_tile_gen_0_cfg_tile_connected_esto;
logic [1:0][31:0] glb_tile_gen_0_cgra_cfg_g2f_cfg_addr;
logic [1:0][31:0] glb_tile_gen_0_cgra_cfg_g2f_cfg_data;
logic [1:0] glb_tile_gen_0_cgra_cfg_g2f_cfg_rd_en;
logic [1:0] glb_tile_gen_0_cgra_cfg_g2f_cfg_wr_en;
logic [31:0] glb_tile_gen_0_cgra_cfg_jtag_addr_bypass_esto;
logic [31:0] glb_tile_gen_0_cgra_cfg_jtag_addr_esto;
logic [31:0] glb_tile_gen_0_cgra_cfg_jtag_data_esto;
logic glb_tile_gen_0_cgra_cfg_jtag_rd_en_bypass_esto;
logic glb_tile_gen_0_cgra_cfg_jtag_rd_en_esto;
logic glb_tile_gen_0_cgra_cfg_jtag_wr_en_esto;
logic [31:0] glb_tile_gen_0_cgra_cfg_pcfg_addr_e2w_wsto;
logic [31:0] glb_tile_gen_0_cgra_cfg_pcfg_addr_w2e_esto;
logic [31:0] glb_tile_gen_0_cgra_cfg_pcfg_data_e2w_wsto;
logic [31:0] glb_tile_gen_0_cgra_cfg_pcfg_data_w2e_esto;
logic glb_tile_gen_0_cgra_cfg_pcfg_rd_en_e2w_wsto;
logic glb_tile_gen_0_cgra_cfg_pcfg_rd_en_w2e_esto;
logic glb_tile_gen_0_cgra_cfg_pcfg_wr_en_e2w_wsto;
logic glb_tile_gen_0_cgra_cfg_pcfg_wr_en_w2e_esto;
logic glb_tile_gen_0_clk_en_bank_master;
logic glb_tile_gen_0_clk_en_master;
logic glb_tile_gen_0_clk_en_pcfg_broadcast;
logic glb_tile_gen_0_data_flush;
logic glb_tile_gen_0_pcfg_g2f_interrupt_pulse;
logic [18:0] glb_tile_gen_0_pcfg_rd_addr_e2w_wsto;
logic [18:0] glb_tile_gen_0_pcfg_rd_addr_w2e_esto;
logic [63:0] glb_tile_gen_0_pcfg_rd_data_e2w_wsto;
logic glb_tile_gen_0_pcfg_rd_data_valid_e2w_wsto;
logic glb_tile_gen_0_pcfg_rd_data_valid_w2e_esto;
logic [63:0] glb_tile_gen_0_pcfg_rd_data_w2e_esto;
logic glb_tile_gen_0_pcfg_rd_en_e2w_wsto;
logic glb_tile_gen_0_pcfg_rd_en_w2e_esto;
logic [1:0][15:0] glb_tile_gen_0_strm_data_g2f;
logic [1:0] glb_tile_gen_0_strm_data_valid_g2f;
logic glb_tile_gen_0_strm_f2g_interrupt_pulse;
logic glb_tile_gen_0_strm_g2f_interrupt_pulse;
logic [18:0] glb_tile_gen_0_strm_rd_addr_e2w_wsto;
logic [18:0] glb_tile_gen_0_strm_rd_addr_w2e_esto;
logic [63:0] glb_tile_gen_0_strm_rd_data_e2w_wsto;
logic glb_tile_gen_0_strm_rd_data_valid_e2w_wsto;
logic glb_tile_gen_0_strm_rd_data_valid_w2e_esto;
logic [63:0] glb_tile_gen_0_strm_rd_data_w2e_esto;
logic glb_tile_gen_0_strm_rd_en_e2w_wsto;
logic glb_tile_gen_0_strm_rd_en_w2e_esto;
logic [18:0] glb_tile_gen_0_strm_wr_addr_e2w_wsto;
logic [18:0] glb_tile_gen_0_strm_wr_addr_w2e_esto;
logic [63:0] glb_tile_gen_0_strm_wr_data_e2w_wsto;
logic [63:0] glb_tile_gen_0_strm_wr_data_w2e_esto;
logic glb_tile_gen_0_strm_wr_en_e2w_wsto;
logic glb_tile_gen_0_strm_wr_en_w2e_esto;
logic [7:0] glb_tile_gen_0_strm_wr_strb_e2w_wsto;
logic [7:0] glb_tile_gen_0_strm_wr_strb_w2e_esto;
logic glb_tile_gen_1_cfg_pcfg_tile_connected_esto;
logic glb_tile_gen_1_cfg_tile_connected_esto;
logic [1:0][31:0] glb_tile_gen_1_cgra_cfg_g2f_cfg_addr;
logic [1:0][31:0] glb_tile_gen_1_cgra_cfg_g2f_cfg_data;
logic [1:0] glb_tile_gen_1_cgra_cfg_g2f_cfg_rd_en;
logic [1:0] glb_tile_gen_1_cgra_cfg_g2f_cfg_wr_en;
logic [31:0] glb_tile_gen_1_cgra_cfg_jtag_addr_bypass_esto;
logic [31:0] glb_tile_gen_1_cgra_cfg_jtag_addr_esto;
logic [31:0] glb_tile_gen_1_cgra_cfg_jtag_data_esto;
logic glb_tile_gen_1_cgra_cfg_jtag_rd_en_bypass_esto;
logic glb_tile_gen_1_cgra_cfg_jtag_rd_en_esto;
logic glb_tile_gen_1_cgra_cfg_jtag_wr_en_esto;
logic [31:0] glb_tile_gen_1_cgra_cfg_pcfg_addr_e2w_wsto;
logic [31:0] glb_tile_gen_1_cgra_cfg_pcfg_addr_w2e_esto;
logic [31:0] glb_tile_gen_1_cgra_cfg_pcfg_data_e2w_wsto;
logic [31:0] glb_tile_gen_1_cgra_cfg_pcfg_data_w2e_esto;
logic glb_tile_gen_1_cgra_cfg_pcfg_rd_en_e2w_wsto;
logic glb_tile_gen_1_cgra_cfg_pcfg_rd_en_w2e_esto;
logic glb_tile_gen_1_cgra_cfg_pcfg_wr_en_e2w_wsto;
logic glb_tile_gen_1_cgra_cfg_pcfg_wr_en_w2e_esto;
logic glb_tile_gen_1_clk_en_bank_master;
logic glb_tile_gen_1_clk_en_master;
logic glb_tile_gen_1_clk_en_pcfg_broadcast;
logic glb_tile_gen_1_data_flush;
logic glb_tile_gen_1_pcfg_g2f_interrupt_pulse;
logic [18:0] glb_tile_gen_1_pcfg_rd_addr_e2w_wsto;
logic [18:0] glb_tile_gen_1_pcfg_rd_addr_w2e_esto;
logic [63:0] glb_tile_gen_1_pcfg_rd_data_e2w_wsto;
logic glb_tile_gen_1_pcfg_rd_data_valid_e2w_wsto;
logic glb_tile_gen_1_pcfg_rd_data_valid_w2e_esto;
logic [63:0] glb_tile_gen_1_pcfg_rd_data_w2e_esto;
logic glb_tile_gen_1_pcfg_rd_en_e2w_wsto;
logic glb_tile_gen_1_pcfg_rd_en_w2e_esto;
logic [1:0][15:0] glb_tile_gen_1_strm_data_g2f;
logic [1:0] glb_tile_gen_1_strm_data_valid_g2f;
logic glb_tile_gen_1_strm_f2g_interrupt_pulse;
logic glb_tile_gen_1_strm_g2f_interrupt_pulse;
logic [18:0] glb_tile_gen_1_strm_rd_addr_e2w_wsto;
logic [18:0] glb_tile_gen_1_strm_rd_addr_w2e_esto;
logic [63:0] glb_tile_gen_1_strm_rd_data_e2w_wsto;
logic glb_tile_gen_1_strm_rd_data_valid_e2w_wsto;
logic glb_tile_gen_1_strm_rd_data_valid_w2e_esto;
logic [63:0] glb_tile_gen_1_strm_rd_data_w2e_esto;
logic glb_tile_gen_1_strm_rd_en_e2w_wsto;
logic glb_tile_gen_1_strm_rd_en_w2e_esto;
logic [18:0] glb_tile_gen_1_strm_wr_addr_e2w_wsto;
logic [18:0] glb_tile_gen_1_strm_wr_addr_w2e_esto;
logic [63:0] glb_tile_gen_1_strm_wr_data_e2w_wsto;
logic [63:0] glb_tile_gen_1_strm_wr_data_w2e_esto;
logic glb_tile_gen_1_strm_wr_en_e2w_wsto;
logic glb_tile_gen_1_strm_wr_en_w2e_esto;
logic [7:0] glb_tile_gen_1_strm_wr_strb_e2w_wsto;
logic [7:0] glb_tile_gen_1_strm_wr_strb_w2e_esto;
logic if_sram_cfg_rd_data_valid_w;
logic [31:0] if_sram_cfg_rd_data_w;
logic [1:0] pcfg_g2f_interrupt_pulse_d;
logic [1:0] pcfg_g2f_interrupt_pulse_w;
rd_packet_t [1:0] pcfg_packet_e2w_esti;
rd_packet_t [1:0] pcfg_packet_e2w_wsto;
rd_packet_t [1:0] pcfg_packet_w2e_esto;
rd_packet_t [1:0] pcfg_packet_w2e_wsti;
logic [18:0] proc_rd_addr_d;
logic proc_rd_addr_sel;
logic proc_rd_clk_en;
logic proc_rd_clk_en_gen_enable;
logic proc_rd_data_valid_w;
logic [63:0] proc_rd_data_w;
logic proc_rd_en_d;
proc_rd_type_e proc_rd_type;
logic [18:0] proc_wr_addr_d;
logic proc_wr_clk_en;
logic proc_wr_clk_en_gen_enable;
logic [63:0] proc_wr_data_d;
logic proc_wr_en_d;
logic [7:0] proc_wr_strb_d;
logic [18:0] sram_cfg_rd_addr_d;
logic sram_cfg_rd_en_d;
logic [18:0] sram_cfg_wr_addr_d;
logic [63:0] sram_cfg_wr_data_d;
logic sram_cfg_wr_en_d;
logic [7:0] sram_cfg_wr_strb_d;
logic [1:0] strm_f2g_interrupt_pulse_d;
logic [1:0] strm_f2g_interrupt_pulse_w;
logic [1:0] strm_g2f_interrupt_pulse_d;
logic [1:0] strm_g2f_interrupt_pulse_w;
packet_t [1:0] strm_packet_e2w_esti;
packet_t [1:0] strm_packet_e2w_wsto;
packet_t [1:0] strm_packet_w2e_esto;
packet_t [1:0] strm_packet_w2e_wsti;
glb_tile_ifc_A_12_D_32 if_cfg_tile2tile_0();
glb_tile_ifc_A_12_D_32 if_cfg_tile2tile_1();
glb_tile_ifc_A_12_D_32 if_cfg_tile2tile_2();
glb_tile_ifc_A_19_D_64 if_proc_tile2tile_0();
glb_tile_ifc_A_19_D_64 if_proc_tile2tile_1();
glb_tile_ifc_A_19_D_64 if_proc_tile2tile_2();
glb_tile_ifc_A_19_D_32 if_sram_cfg_tile2tile_0();
glb_tile_ifc_A_19_D_32 if_sram_cfg_tile2tile_1();
glb_tile_ifc_A_19_D_32 if_sram_cfg_tile2tile_2();
assign cfg_tile_connected[0] = 1'h0;
assign cfg_pcfg_tile_connected[0] = 1'h0;
assign strm_f2g_interrupt_pulse = strm_f2g_interrupt_pulse_d;
assign strm_g2f_interrupt_pulse = strm_g2f_interrupt_pulse_d;
assign pcfg_g2f_interrupt_pulse = pcfg_g2f_interrupt_pulse_d;
assign cgra_stall = cgra_stall_in;
assign if_sram_cfg_tile2tile_2.rd_data = 32'h0;
assign if_sram_cfg_tile2tile_2.rd_data_valid = 1'h0;
assign glb_tile_gen_0_clk_en_pcfg_broadcast = ~pcfg_broadcast_stall[0];
assign glb_tile_gen_0_clk_en_master = glb_clk_en_master[0];
assign glb_tile_gen_0_clk_en_bank_master = glb_clk_en_bank_master[0];
assign strm_packet_w2e_esto[0].wr.wr_en = glb_tile_gen_0_strm_wr_en_w2e_esto;
assign strm_packet_w2e_esto[0].wr.wr_strb = glb_tile_gen_0_strm_wr_strb_w2e_esto;
assign strm_packet_w2e_esto[0].wr.wr_addr = glb_tile_gen_0_strm_wr_addr_w2e_esto;
assign strm_packet_w2e_esto[0].wr.wr_data = glb_tile_gen_0_strm_wr_data_w2e_esto;
assign strm_packet_w2e_esto[0].rdrq.rd_en = glb_tile_gen_0_strm_rd_en_w2e_esto;
assign strm_packet_w2e_esto[0].rdrq.rd_addr = glb_tile_gen_0_strm_rd_addr_w2e_esto;
assign strm_packet_w2e_esto[0].rdrs.rd_data = glb_tile_gen_0_strm_rd_data_w2e_esto;
assign strm_packet_w2e_esto[0].rdrs.rd_data_valid = glb_tile_gen_0_strm_rd_data_valid_w2e_esto;
assign strm_packet_e2w_wsto[0].wr.wr_en = glb_tile_gen_0_strm_wr_en_e2w_wsto;
assign strm_packet_e2w_wsto[0].wr.wr_strb = glb_tile_gen_0_strm_wr_strb_e2w_wsto;
assign strm_packet_e2w_wsto[0].wr.wr_addr = glb_tile_gen_0_strm_wr_addr_e2w_wsto;
assign strm_packet_e2w_wsto[0].wr.wr_data = glb_tile_gen_0_strm_wr_data_e2w_wsto;
assign strm_packet_e2w_wsto[0].rdrq.rd_en = glb_tile_gen_0_strm_rd_en_e2w_wsto;
assign strm_packet_e2w_wsto[0].rdrq.rd_addr = glb_tile_gen_0_strm_rd_addr_e2w_wsto;
assign strm_packet_e2w_wsto[0].rdrs.rd_data = glb_tile_gen_0_strm_rd_data_e2w_wsto;
assign strm_packet_e2w_wsto[0].rdrs.rd_data_valid = glb_tile_gen_0_strm_rd_data_valid_e2w_wsto;
assign pcfg_packet_w2e_esto[0].rdrq.rd_en = glb_tile_gen_0_pcfg_rd_en_w2e_esto;
assign pcfg_packet_w2e_esto[0].rdrq.rd_addr = glb_tile_gen_0_pcfg_rd_addr_w2e_esto;
assign pcfg_packet_w2e_esto[0].rdrs.rd_data = glb_tile_gen_0_pcfg_rd_data_w2e_esto;
assign pcfg_packet_w2e_esto[0].rdrs.rd_data_valid = glb_tile_gen_0_pcfg_rd_data_valid_w2e_esto;
assign pcfg_packet_e2w_wsto[0].rdrq.rd_en = glb_tile_gen_0_pcfg_rd_en_e2w_wsto;
assign pcfg_packet_e2w_wsto[0].rdrq.rd_addr = glb_tile_gen_0_pcfg_rd_addr_e2w_wsto;
assign pcfg_packet_e2w_wsto[0].rdrs.rd_data = glb_tile_gen_0_pcfg_rd_data_e2w_wsto;
assign pcfg_packet_e2w_wsto[0].rdrs.rd_data_valid = glb_tile_gen_0_pcfg_rd_data_valid_e2w_wsto;
assign cfg_tile_connected[1] = glb_tile_gen_0_cfg_tile_connected_esto;
assign cfg_pcfg_tile_connected[1] = glb_tile_gen_0_cfg_pcfg_tile_connected_esto;
assign strm_data_g2f[0] = glb_tile_gen_0_strm_data_g2f;
assign strm_data_valid_g2f[0] = glb_tile_gen_0_strm_data_valid_g2f;
assign data_flush[0] = glb_tile_gen_0_data_flush;
assign cgra_cfg_g2f_cfg_wr_en[0] = glb_tile_gen_0_cgra_cfg_g2f_cfg_wr_en;
assign cgra_cfg_g2f_cfg_rd_en[0] = glb_tile_gen_0_cgra_cfg_g2f_cfg_rd_en;
assign cgra_cfg_g2f_cfg_addr[0] = glb_tile_gen_0_cgra_cfg_g2f_cfg_addr;
assign cgra_cfg_g2f_cfg_data[0] = glb_tile_gen_0_cgra_cfg_g2f_cfg_data;
assign cgra_cfg_pcfg_wr_en_esto[0] = glb_tile_gen_0_cgra_cfg_pcfg_wr_en_w2e_esto;
assign cgra_cfg_pcfg_rd_en_esto[0] = glb_tile_gen_0_cgra_cfg_pcfg_rd_en_w2e_esto;
assign cgra_cfg_pcfg_addr_esto[0] = glb_tile_gen_0_cgra_cfg_pcfg_addr_w2e_esto;
assign cgra_cfg_pcfg_data_esto[0] = glb_tile_gen_0_cgra_cfg_pcfg_data_w2e_esto;
assign cgra_cfg_pcfg_wr_en_wsto[0] = glb_tile_gen_0_cgra_cfg_pcfg_wr_en_e2w_wsto;
assign cgra_cfg_pcfg_rd_en_wsto[0] = glb_tile_gen_0_cgra_cfg_pcfg_rd_en_e2w_wsto;
assign cgra_cfg_pcfg_addr_wsto[0] = glb_tile_gen_0_cgra_cfg_pcfg_addr_e2w_wsto;
assign cgra_cfg_pcfg_data_wsto[0] = glb_tile_gen_0_cgra_cfg_pcfg_data_e2w_wsto;
assign cgra_cfg_jtag_wr_en_esto[0] = glb_tile_gen_0_cgra_cfg_jtag_wr_en_esto;
assign cgra_cfg_jtag_rd_en_esto[0] = glb_tile_gen_0_cgra_cfg_jtag_rd_en_esto;
assign cgra_cfg_jtag_addr_esto[0] = glb_tile_gen_0_cgra_cfg_jtag_addr_esto;
assign cgra_cfg_jtag_data_esto[0] = glb_tile_gen_0_cgra_cfg_jtag_data_esto;
assign cgra_cfg_jtag_rd_en_bypass_esto[0] = glb_tile_gen_0_cgra_cfg_jtag_rd_en_bypass_esto;
assign cgra_cfg_jtag_addr_bypass_esto[0] = glb_tile_gen_0_cgra_cfg_jtag_addr_bypass_esto;
assign strm_f2g_interrupt_pulse_w[0] = glb_tile_gen_0_strm_f2g_interrupt_pulse;
assign strm_g2f_interrupt_pulse_w[0] = glb_tile_gen_0_strm_g2f_interrupt_pulse;
assign pcfg_g2f_interrupt_pulse_w[0] = glb_tile_gen_0_pcfg_g2f_interrupt_pulse;
assign glb_tile_gen_1_clk_en_pcfg_broadcast = ~pcfg_broadcast_stall[1];
assign glb_tile_gen_1_clk_en_master = glb_clk_en_master[1];
assign glb_tile_gen_1_clk_en_bank_master = glb_clk_en_bank_master[1];
assign strm_packet_w2e_esto[1].wr.wr_en = glb_tile_gen_1_strm_wr_en_w2e_esto;
assign strm_packet_w2e_esto[1].wr.wr_strb = glb_tile_gen_1_strm_wr_strb_w2e_esto;
assign strm_packet_w2e_esto[1].wr.wr_addr = glb_tile_gen_1_strm_wr_addr_w2e_esto;
assign strm_packet_w2e_esto[1].wr.wr_data = glb_tile_gen_1_strm_wr_data_w2e_esto;
assign strm_packet_w2e_esto[1].rdrq.rd_en = glb_tile_gen_1_strm_rd_en_w2e_esto;
assign strm_packet_w2e_esto[1].rdrq.rd_addr = glb_tile_gen_1_strm_rd_addr_w2e_esto;
assign strm_packet_w2e_esto[1].rdrs.rd_data = glb_tile_gen_1_strm_rd_data_w2e_esto;
assign strm_packet_w2e_esto[1].rdrs.rd_data_valid = glb_tile_gen_1_strm_rd_data_valid_w2e_esto;
assign strm_packet_e2w_wsto[1].wr.wr_en = glb_tile_gen_1_strm_wr_en_e2w_wsto;
assign strm_packet_e2w_wsto[1].wr.wr_strb = glb_tile_gen_1_strm_wr_strb_e2w_wsto;
assign strm_packet_e2w_wsto[1].wr.wr_addr = glb_tile_gen_1_strm_wr_addr_e2w_wsto;
assign strm_packet_e2w_wsto[1].wr.wr_data = glb_tile_gen_1_strm_wr_data_e2w_wsto;
assign strm_packet_e2w_wsto[1].rdrq.rd_en = glb_tile_gen_1_strm_rd_en_e2w_wsto;
assign strm_packet_e2w_wsto[1].rdrq.rd_addr = glb_tile_gen_1_strm_rd_addr_e2w_wsto;
assign strm_packet_e2w_wsto[1].rdrs.rd_data = glb_tile_gen_1_strm_rd_data_e2w_wsto;
assign strm_packet_e2w_wsto[1].rdrs.rd_data_valid = glb_tile_gen_1_strm_rd_data_valid_e2w_wsto;
assign pcfg_packet_w2e_esto[1].rdrq.rd_en = glb_tile_gen_1_pcfg_rd_en_w2e_esto;
assign pcfg_packet_w2e_esto[1].rdrq.rd_addr = glb_tile_gen_1_pcfg_rd_addr_w2e_esto;
assign pcfg_packet_w2e_esto[1].rdrs.rd_data = glb_tile_gen_1_pcfg_rd_data_w2e_esto;
assign pcfg_packet_w2e_esto[1].rdrs.rd_data_valid = glb_tile_gen_1_pcfg_rd_data_valid_w2e_esto;
assign pcfg_packet_e2w_wsto[1].rdrq.rd_en = glb_tile_gen_1_pcfg_rd_en_e2w_wsto;
assign pcfg_packet_e2w_wsto[1].rdrq.rd_addr = glb_tile_gen_1_pcfg_rd_addr_e2w_wsto;
assign pcfg_packet_e2w_wsto[1].rdrs.rd_data = glb_tile_gen_1_pcfg_rd_data_e2w_wsto;
assign pcfg_packet_e2w_wsto[1].rdrs.rd_data_valid = glb_tile_gen_1_pcfg_rd_data_valid_e2w_wsto;
assign cfg_tile_connected[2] = glb_tile_gen_1_cfg_tile_connected_esto;
assign cfg_pcfg_tile_connected[2] = glb_tile_gen_1_cfg_pcfg_tile_connected_esto;
assign strm_data_g2f[1] = glb_tile_gen_1_strm_data_g2f;
assign strm_data_valid_g2f[1] = glb_tile_gen_1_strm_data_valid_g2f;
assign data_flush[1] = glb_tile_gen_1_data_flush;
assign cgra_cfg_g2f_cfg_wr_en[1] = glb_tile_gen_1_cgra_cfg_g2f_cfg_wr_en;
assign cgra_cfg_g2f_cfg_rd_en[1] = glb_tile_gen_1_cgra_cfg_g2f_cfg_rd_en;
assign cgra_cfg_g2f_cfg_addr[1] = glb_tile_gen_1_cgra_cfg_g2f_cfg_addr;
assign cgra_cfg_g2f_cfg_data[1] = glb_tile_gen_1_cgra_cfg_g2f_cfg_data;
assign cgra_cfg_pcfg_wr_en_esto[1] = glb_tile_gen_1_cgra_cfg_pcfg_wr_en_w2e_esto;
assign cgra_cfg_pcfg_rd_en_esto[1] = glb_tile_gen_1_cgra_cfg_pcfg_rd_en_w2e_esto;
assign cgra_cfg_pcfg_addr_esto[1] = glb_tile_gen_1_cgra_cfg_pcfg_addr_w2e_esto;
assign cgra_cfg_pcfg_data_esto[1] = glb_tile_gen_1_cgra_cfg_pcfg_data_w2e_esto;
assign cgra_cfg_pcfg_wr_en_wsto[1] = glb_tile_gen_1_cgra_cfg_pcfg_wr_en_e2w_wsto;
assign cgra_cfg_pcfg_rd_en_wsto[1] = glb_tile_gen_1_cgra_cfg_pcfg_rd_en_e2w_wsto;
assign cgra_cfg_pcfg_addr_wsto[1] = glb_tile_gen_1_cgra_cfg_pcfg_addr_e2w_wsto;
assign cgra_cfg_pcfg_data_wsto[1] = glb_tile_gen_1_cgra_cfg_pcfg_data_e2w_wsto;
assign cgra_cfg_jtag_wr_en_esto[1] = glb_tile_gen_1_cgra_cfg_jtag_wr_en_esto;
assign cgra_cfg_jtag_rd_en_esto[1] = glb_tile_gen_1_cgra_cfg_jtag_rd_en_esto;
assign cgra_cfg_jtag_addr_esto[1] = glb_tile_gen_1_cgra_cfg_jtag_addr_esto;
assign cgra_cfg_jtag_data_esto[1] = glb_tile_gen_1_cgra_cfg_jtag_data_esto;
assign cgra_cfg_jtag_rd_en_bypass_esto[1] = glb_tile_gen_1_cgra_cfg_jtag_rd_en_bypass_esto;
assign cgra_cfg_jtag_addr_bypass_esto[1] = glb_tile_gen_1_cgra_cfg_jtag_addr_bypass_esto;
assign strm_f2g_interrupt_pulse_w[1] = glb_tile_gen_1_strm_f2g_interrupt_pulse;
assign strm_g2f_interrupt_pulse_w[1] = glb_tile_gen_1_strm_g2f_interrupt_pulse;
assign pcfg_g2f_interrupt_pulse_w[1] = glb_tile_gen_1_pcfg_g2f_interrupt_pulse;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    proc_wr_en_d <= 1'h0;
    proc_wr_strb_d <= 8'h0;
    proc_wr_addr_d <= 19'h0;
    proc_wr_data_d <= 64'h0;
    proc_rd_en_d <= 1'h0;
    proc_rd_addr_d <= 19'h0;
  end
  else begin
    proc_wr_en_d <= proc_wr_en;
    proc_wr_strb_d <= proc_wr_strb;
    proc_wr_addr_d <= proc_wr_addr;
    proc_wr_data_d <= proc_wr_data;
    proc_rd_en_d <= proc_rd_en;
    proc_rd_addr_d <= proc_rd_addr;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    sram_cfg_wr_en_d <= 1'h0;
    sram_cfg_wr_strb_d <= 8'h0;
    sram_cfg_wr_addr_d <= 19'h0;
    sram_cfg_wr_data_d <= 64'h0;
    sram_cfg_rd_en_d <= 1'h0;
    sram_cfg_rd_addr_d <= 19'h0;
  end
  else begin
    sram_cfg_wr_en_d <= if_sram_cfg_wr_en;
    sram_cfg_wr_addr_d <= if_sram_cfg_wr_addr;
    if (if_sram_cfg_wr_addr[2] == 1'h0) begin
      sram_cfg_wr_data_d <= {32'h0, if_sram_cfg_wr_data};
      sram_cfg_wr_strb_d <= {4'h0, 4'hF};
    end
    else begin
      sram_cfg_wr_data_d <= {if_sram_cfg_wr_data[31:0], 32'h0};
      sram_cfg_wr_strb_d <= {4'hF, 4'h0};
    end
    sram_cfg_rd_en_d <= if_sram_cfg_rd_en;
    sram_cfg_rd_addr_d <= if_sram_cfg_rd_addr;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    if_proc_tile2tile_0.wr_en <= 1'h0;
    if_proc_tile2tile_0.wr_strb <= 8'h0;
    if_proc_tile2tile_0.wr_addr <= 19'h0;
    if_proc_tile2tile_0.wr_data <= 64'h0;
  end
  else if (proc_wr_en_d) begin
    if_proc_tile2tile_0.wr_en <= proc_wr_en_d;
    if_proc_tile2tile_0.wr_strb <= proc_wr_strb_d;
    if_proc_tile2tile_0.wr_addr <= proc_wr_addr_d;
    if_proc_tile2tile_0.wr_data <= proc_wr_data_d;
  end
  else if (sram_cfg_wr_en_d) begin
    if_proc_tile2tile_0.wr_en <= sram_cfg_wr_en_d;
    if_proc_tile2tile_0.wr_strb <= sram_cfg_wr_strb_d;
    if_proc_tile2tile_0.wr_addr <= sram_cfg_wr_addr_d;
    if_proc_tile2tile_0.wr_data <= sram_cfg_wr_data_d;
  end
  else begin
    if_proc_tile2tile_0.wr_en <= proc_wr_en_d;
    if_proc_tile2tile_0.wr_strb <= proc_wr_strb_d;
    if_proc_tile2tile_0.wr_addr <= proc_wr_addr_d;
    if_proc_tile2tile_0.wr_data <= proc_wr_data_d;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    if_proc_tile2tile_0.rd_en <= 1'h0;
    if_proc_tile2tile_0.rd_addr <= 19'h0;
    proc_rd_type <= axi;
    proc_rd_addr_sel <= 1'h0;
  end
  else if (proc_rd_en_d) begin
    if_proc_tile2tile_0.rd_en <= proc_rd_en_d;
    if_proc_tile2tile_0.rd_addr <= proc_rd_addr_d;
    proc_rd_type <= axi;
    proc_rd_addr_sel <= 1'h0;
  end
  else if (sram_cfg_rd_en_d) begin
    if_proc_tile2tile_0.rd_en <= sram_cfg_rd_en_d;
    if_proc_tile2tile_0.rd_addr <= sram_cfg_rd_addr_d;
    proc_rd_addr_sel <= sram_cfg_rd_addr_d[2];
    proc_rd_type <= jtag;
  end
  else begin
    if_proc_tile2tile_0.rd_en <= proc_rd_en_d;
    if_proc_tile2tile_0.rd_addr <= proc_rd_addr_d;
    proc_rd_type <= proc_rd_type;
    proc_rd_addr_sel <= proc_rd_addr_sel;
  end
end
always_comb begin
  if (proc_rd_type == axi) begin
    proc_rd_data_w = if_proc_tile2tile_0.rd_data;
    proc_rd_data_valid_w = if_proc_tile2tile_0.rd_data_valid;
    if_sram_cfg_rd_data_w = 32'h0;
    if_sram_cfg_rd_data_valid_w = 1'h0;
  end
  else if (proc_rd_type == jtag) begin
    proc_rd_data_w = 64'h0;
    proc_rd_data_valid_w = 1'h0;
    if (proc_rd_addr_sel == 1'h0) begin
      if_sram_cfg_rd_data_w = if_proc_tile2tile_0.rd_data[31:0];
    end
    else if_sram_cfg_rd_data_w = if_proc_tile2tile_0.rd_data[63:32];
    if_sram_cfg_rd_data_valid_w = if_proc_tile2tile_0.rd_data_valid;
  end
  else begin
    proc_rd_data_w = if_proc_tile2tile_0.rd_data;
    proc_rd_data_valid_w = if_proc_tile2tile_0.rd_data_valid;
    if_sram_cfg_rd_data_w = 32'h0;
    if_sram_cfg_rd_data_valid_w = 1'h0;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    proc_rd_data <= 64'h0;
    proc_rd_data_valid <= 1'h0;
    if_sram_cfg_rd_data <= 32'h0;
    if_sram_cfg_rd_data_valid <= 1'h0;
  end
  else begin
    proc_rd_data <= proc_rd_data_w;
    proc_rd_data_valid <= proc_rd_data_valid_w;
    if_sram_cfg_rd_data <= if_sram_cfg_rd_data_w;
    if_sram_cfg_rd_data_valid <= if_sram_cfg_rd_data_valid_w;
  end
end
assign proc_wr_clk_en_gen_enable = proc_wr_en_d | sram_cfg_wr_en_d;
assign if_proc_tile2tile_0.wr_clk_en = proc_wr_clk_en;
assign proc_rd_clk_en_gen_enable = proc_rd_en_d | sram_cfg_rd_en_d;
assign if_proc_tile2tile_0.rd_clk_en = proc_rd_clk_en;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    if_cfg_tile2tile_0.wr_en <= 1'h0;
    if_cfg_tile2tile_0.wr_clk_en <= 1'h0;
    if_cfg_tile2tile_0.wr_addr <= 12'h0;
    if_cfg_tile2tile_0.wr_data <= 32'h0;
    if_cfg_tile2tile_0.rd_en <= 1'h0;
    if_cfg_tile2tile_0.rd_clk_en <= 1'h0;
    if_cfg_tile2tile_0.rd_addr <= 12'h0;
  end
  else begin
    if_cfg_tile2tile_0.wr_en <= if_cfg_wr_en;
    if_cfg_tile2tile_0.wr_clk_en <= if_cfg_wr_clk_en;
    if_cfg_tile2tile_0.wr_addr <= if_cfg_wr_addr;
    if_cfg_tile2tile_0.wr_data <= if_cfg_wr_data;
    if_cfg_tile2tile_0.rd_en <= if_cfg_rd_en;
    if_cfg_tile2tile_0.rd_clk_en <= if_cfg_rd_clk_en;
    if_cfg_tile2tile_0.rd_addr <= if_cfg_rd_addr;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    cgra_cfg_jtag_gc2glb_wr_en_d <= 1'h0;
    cgra_cfg_jtag_gc2glb_rd_en_d <= 1'h0;
    cgra_cfg_jtag_gc2glb_addr_d <= 32'h0;
    cgra_cfg_jtag_gc2glb_data_d <= 32'h0;
  end
  else begin
    cgra_cfg_jtag_gc2glb_wr_en_d <= cgra_cfg_jtag_gc2glb_wr_en;
    cgra_cfg_jtag_gc2glb_rd_en_d <= cgra_cfg_jtag_gc2glb_rd_en;
    cgra_cfg_jtag_gc2glb_addr_d <= cgra_cfg_jtag_gc2glb_addr;
    cgra_cfg_jtag_gc2glb_data_d <= cgra_cfg_jtag_gc2glb_data;
  end
end
assign strm_packet_e2w_esti[1] = 177'h0;
assign pcfg_packet_e2w_esti[1] = 85'h0;
assign strm_packet_e2w_esti[0] = strm_packet_e2w_wsto[1];
assign pcfg_packet_e2w_esti[0] = pcfg_packet_e2w_wsto[1];
assign strm_packet_w2e_wsti[0] = 177'h0;
assign pcfg_packet_w2e_wsti[0] = 85'h0;
assign strm_packet_w2e_wsti[1] = strm_packet_w2e_esto[0];
assign pcfg_packet_w2e_wsti[1] = pcfg_packet_w2e_esto[0];
always_comb begin
  cgra_cfg_jtag_rd_en_wsti[0] = 1'h0;
  cgra_cfg_jtag_wr_en_wsti[0] = cgra_cfg_jtag_gc2glb_wr_en_d;
  cgra_cfg_jtag_addr_wsti[0] = cgra_cfg_jtag_gc2glb_addr_d;
  cgra_cfg_jtag_data_wsti[0] = cgra_cfg_jtag_gc2glb_data_d;
  cgra_cfg_jtag_rd_en_bypass_wsti[0] = cgra_cfg_jtag_gc2glb_rd_en_d;
  cgra_cfg_jtag_addr_bypass_wsti[0] = cgra_cfg_jtag_gc2glb_addr_d;
  cgra_cfg_pcfg_rd_en_wsti[0] = 1'h0;
  cgra_cfg_pcfg_wr_en_wsti[0] = 1'h0;
  cgra_cfg_pcfg_addr_wsti[0] = 32'h0;
  cgra_cfg_pcfg_data_wsti[0] = 32'h0;
  cgra_cfg_jtag_rd_en_wsti[1] = cgra_cfg_jtag_rd_en_esto[0];
  cgra_cfg_jtag_wr_en_wsti[1] = cgra_cfg_jtag_wr_en_esto[0];
  cgra_cfg_jtag_addr_wsti[1] = cgra_cfg_jtag_addr_esto[0];
  cgra_cfg_jtag_data_wsti[1] = cgra_cfg_jtag_data_esto[0];
  cgra_cfg_jtag_rd_en_bypass_wsti[1] = cgra_cfg_jtag_rd_en_bypass_esto[0];
  cgra_cfg_jtag_addr_bypass_wsti[1] = cgra_cfg_jtag_addr_bypass_esto[0];
  cgra_cfg_pcfg_rd_en_wsti[1] = cgra_cfg_pcfg_rd_en_esto[0];
  cgra_cfg_pcfg_wr_en_wsti[1] = cgra_cfg_pcfg_wr_en_esto[0];
  cgra_cfg_pcfg_addr_wsti[1] = cgra_cfg_pcfg_addr_esto[0];
  cgra_cfg_pcfg_data_wsti[1] = cgra_cfg_pcfg_data_esto[0];
end
always_comb begin
  cgra_cfg_pcfg_rd_en_esti[0] = cgra_cfg_pcfg_rd_en_wsto[1];
  cgra_cfg_pcfg_wr_en_esti[0] = cgra_cfg_pcfg_wr_en_wsto[1];
  cgra_cfg_pcfg_addr_esti[0] = cgra_cfg_pcfg_addr_wsto[1];
  cgra_cfg_pcfg_data_esti[0] = cgra_cfg_pcfg_data_wsto[1];
  cgra_cfg_pcfg_rd_en_esti[1] = 1'h0;
  cgra_cfg_pcfg_wr_en_esti[1] = 1'h0;
  cgra_cfg_pcfg_addr_esti[1] = 32'h0;
  cgra_cfg_pcfg_data_esti[1] = 32'h0;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    for (int unsigned i = 0; i < 2; i += 1) begin
        strm_f2g_interrupt_pulse_d[1'(i)] <= 1'h0;
        strm_g2f_interrupt_pulse_d[1'(i)] <= 1'h0;
        pcfg_g2f_interrupt_pulse_d[1'(i)] <= 1'h0;
      end
  end
  else begin
    for (int unsigned i = 0; i < 2; i += 1) begin
        strm_f2g_interrupt_pulse_d[1'(i)] <= strm_f2g_interrupt_pulse_w[1'(i)];
        strm_g2f_interrupt_pulse_d[1'(i)] <= strm_g2f_interrupt_pulse_w[1'(i)];
        pcfg_g2f_interrupt_pulse_d[1'(i)] <= pcfg_g2f_interrupt_pulse_w[1'(i)];
      end
  end
end
assign if_cfg_rd_data = if_cfg_tile2tile_0.rd_data;
assign if_cfg_rd_data_valid = if_cfg_tile2tile_0.rd_data_valid;
assign flush_crossbar_in[0] = data_flush_d[0];
assign flush_crossbar_in[1] = data_flush_d[1];
assign flush_crossbar_sel_w = flush_crossbar_sel;
glb_tile glb_tile_gen_0 (
  .cfg_pcfg_tile_connected_wsti(cfg_pcfg_tile_connected[0]),
  .cfg_tile_connected_wsti(cfg_tile_connected[0]),
  .cgra_cfg_jtag_addr_bypass_wsti(cgra_cfg_jtag_addr_bypass_wsti[0]),
  .cgra_cfg_jtag_addr_wsti(cgra_cfg_jtag_addr_wsti[0]),
  .cgra_cfg_jtag_data_wsti(cgra_cfg_jtag_data_wsti[0]),
  .cgra_cfg_jtag_rd_en_bypass_wsti(cgra_cfg_jtag_rd_en_bypass_wsti[0]),
  .cgra_cfg_jtag_rd_en_wsti(cgra_cfg_jtag_rd_en_wsti[0]),
  .cgra_cfg_jtag_wr_en_wsti(cgra_cfg_jtag_wr_en_wsti[0]),
  .cgra_cfg_pcfg_addr_e2w_esti(cgra_cfg_pcfg_addr_esti[0]),
  .cgra_cfg_pcfg_addr_w2e_wsti(cgra_cfg_pcfg_addr_wsti[0]),
  .cgra_cfg_pcfg_data_e2w_esti(cgra_cfg_pcfg_data_esti[0]),
  .cgra_cfg_pcfg_data_w2e_wsti(cgra_cfg_pcfg_data_wsti[0]),
  .cgra_cfg_pcfg_rd_en_e2w_esti(cgra_cfg_pcfg_rd_en_esti[0]),
  .cgra_cfg_pcfg_rd_en_w2e_wsti(cgra_cfg_pcfg_rd_en_wsti[0]),
  .cgra_cfg_pcfg_wr_en_e2w_esti(cgra_cfg_pcfg_wr_en_esti[0]),
  .cgra_cfg_pcfg_wr_en_w2e_wsti(cgra_cfg_pcfg_wr_en_wsti[0]),
  .clk(clk),
  .clk_en_bank_master(glb_tile_gen_0_clk_en_bank_master),
  .clk_en_master(glb_tile_gen_0_clk_en_master),
  .clk_en_pcfg_broadcast(glb_tile_gen_0_clk_en_pcfg_broadcast),
  .glb_tile_id(1'h0),
  .if_cfg_est_m_rd_data(if_cfg_tile2tile_1.rd_data),
  .if_cfg_est_m_rd_data_valid(if_cfg_tile2tile_1.rd_data_valid),
  .if_cfg_wst_s_rd_addr(if_cfg_tile2tile_0.rd_addr),
  .if_cfg_wst_s_rd_clk_en(if_cfg_tile2tile_0.rd_clk_en),
  .if_cfg_wst_s_rd_en(if_cfg_tile2tile_0.rd_en),
  .if_cfg_wst_s_wr_addr(if_cfg_tile2tile_0.wr_addr),
  .if_cfg_wst_s_wr_clk_en(if_cfg_tile2tile_0.wr_clk_en),
  .if_cfg_wst_s_wr_data(if_cfg_tile2tile_0.wr_data),
  .if_cfg_wst_s_wr_en(if_cfg_tile2tile_0.wr_en),
  .if_proc_est_m_rd_data(if_proc_tile2tile_1.rd_data),
  .if_proc_est_m_rd_data_valid(if_proc_tile2tile_1.rd_data_valid),
  .if_proc_wst_s_rd_addr(if_proc_tile2tile_0.rd_addr),
  .if_proc_wst_s_rd_clk_en(if_proc_tile2tile_0.rd_clk_en),
  .if_proc_wst_s_rd_en(if_proc_tile2tile_0.rd_en),
  .if_proc_wst_s_wr_addr(if_proc_tile2tile_0.wr_addr),
  .if_proc_wst_s_wr_clk_en(if_proc_tile2tile_0.wr_clk_en),
  .if_proc_wst_s_wr_data(if_proc_tile2tile_0.wr_data),
  .if_proc_wst_s_wr_en(if_proc_tile2tile_0.wr_en),
  .if_proc_wst_s_wr_strb(if_proc_tile2tile_0.wr_strb),
  .pcfg_rd_addr_e2w_esti(pcfg_packet_e2w_esti[0].rdrq.rd_addr),
  .pcfg_rd_addr_w2e_wsti(pcfg_packet_w2e_wsti[0].rdrq.rd_addr),
  .pcfg_rd_data_e2w_esti(pcfg_packet_e2w_esti[0].rdrs.rd_data),
  .pcfg_rd_data_valid_e2w_esti(pcfg_packet_e2w_esti[0].rdrs.rd_data_valid),
  .pcfg_rd_data_valid_w2e_wsti(pcfg_packet_w2e_wsti[0].rdrs.rd_data_valid),
  .pcfg_rd_data_w2e_wsti(pcfg_packet_w2e_wsti[0].rdrs.rd_data),
  .pcfg_rd_en_e2w_esti(pcfg_packet_e2w_esti[0].rdrq.rd_en),
  .pcfg_rd_en_w2e_wsti(pcfg_packet_w2e_wsti[0].rdrq.rd_en),
  .pcfg_start_pulse(pcfg_start_pulse[0]),
  .reset(reset),
  .strm_data_f2g(strm_data_f2g[0]),
  .strm_data_valid_f2g(strm_data_valid_f2g[0]),
  .strm_f2g_start_pulse(strm_f2g_start_pulse[0]),
  .strm_g2f_start_pulse(strm_g2f_start_pulse[0]),
  .strm_rd_addr_e2w_esti(strm_packet_e2w_esti[0].rdrq.rd_addr),
  .strm_rd_addr_w2e_wsti(strm_packet_w2e_wsti[0].rdrq.rd_addr),
  .strm_rd_data_e2w_esti(strm_packet_e2w_esti[0].rdrs.rd_data),
  .strm_rd_data_valid_e2w_esti(strm_packet_e2w_esti[0].rdrs.rd_data_valid),
  .strm_rd_data_valid_w2e_wsti(strm_packet_w2e_wsti[0].rdrs.rd_data_valid),
  .strm_rd_data_w2e_wsti(strm_packet_w2e_wsti[0].rdrs.rd_data),
  .strm_rd_en_e2w_esti(strm_packet_e2w_esti[0].rdrq.rd_en),
  .strm_rd_en_w2e_wsti(strm_packet_w2e_wsti[0].rdrq.rd_en),
  .strm_wr_addr_e2w_esti(strm_packet_e2w_esti[0].wr.wr_addr),
  .strm_wr_addr_w2e_wsti(strm_packet_w2e_wsti[0].wr.wr_addr),
  .strm_wr_data_e2w_esti(strm_packet_e2w_esti[0].wr.wr_data),
  .strm_wr_data_w2e_wsti(strm_packet_w2e_wsti[0].wr.wr_data),
  .strm_wr_en_e2w_esti(strm_packet_e2w_esti[0].wr.wr_en),
  .strm_wr_en_w2e_wsti(strm_packet_w2e_wsti[0].wr.wr_en),
  .strm_wr_strb_e2w_esti(strm_packet_e2w_esti[0].wr.wr_strb),
  .strm_wr_strb_w2e_wsti(strm_packet_w2e_wsti[0].wr.wr_strb),
  .cfg_pcfg_tile_connected_esto(glb_tile_gen_0_cfg_pcfg_tile_connected_esto),
  .cfg_tile_connected_esto(glb_tile_gen_0_cfg_tile_connected_esto),
  .cgra_cfg_g2f_cfg_addr(glb_tile_gen_0_cgra_cfg_g2f_cfg_addr),
  .cgra_cfg_g2f_cfg_data(glb_tile_gen_0_cgra_cfg_g2f_cfg_data),
  .cgra_cfg_g2f_cfg_rd_en(glb_tile_gen_0_cgra_cfg_g2f_cfg_rd_en),
  .cgra_cfg_g2f_cfg_wr_en(glb_tile_gen_0_cgra_cfg_g2f_cfg_wr_en),
  .cgra_cfg_jtag_addr_bypass_esto(glb_tile_gen_0_cgra_cfg_jtag_addr_bypass_esto),
  .cgra_cfg_jtag_addr_esto(glb_tile_gen_0_cgra_cfg_jtag_addr_esto),
  .cgra_cfg_jtag_data_esto(glb_tile_gen_0_cgra_cfg_jtag_data_esto),
  .cgra_cfg_jtag_rd_en_bypass_esto(glb_tile_gen_0_cgra_cfg_jtag_rd_en_bypass_esto),
  .cgra_cfg_jtag_rd_en_esto(glb_tile_gen_0_cgra_cfg_jtag_rd_en_esto),
  .cgra_cfg_jtag_wr_en_esto(glb_tile_gen_0_cgra_cfg_jtag_wr_en_esto),
  .cgra_cfg_pcfg_addr_e2w_wsto(glb_tile_gen_0_cgra_cfg_pcfg_addr_e2w_wsto),
  .cgra_cfg_pcfg_addr_w2e_esto(glb_tile_gen_0_cgra_cfg_pcfg_addr_w2e_esto),
  .cgra_cfg_pcfg_data_e2w_wsto(glb_tile_gen_0_cgra_cfg_pcfg_data_e2w_wsto),
  .cgra_cfg_pcfg_data_w2e_esto(glb_tile_gen_0_cgra_cfg_pcfg_data_w2e_esto),
  .cgra_cfg_pcfg_rd_en_e2w_wsto(glb_tile_gen_0_cgra_cfg_pcfg_rd_en_e2w_wsto),
  .cgra_cfg_pcfg_rd_en_w2e_esto(glb_tile_gen_0_cgra_cfg_pcfg_rd_en_w2e_esto),
  .cgra_cfg_pcfg_wr_en_e2w_wsto(glb_tile_gen_0_cgra_cfg_pcfg_wr_en_e2w_wsto),
  .cgra_cfg_pcfg_wr_en_w2e_esto(glb_tile_gen_0_cgra_cfg_pcfg_wr_en_w2e_esto),
  .data_flush(glb_tile_gen_0_data_flush),
  .if_cfg_est_m_rd_addr(if_cfg_tile2tile_1.rd_addr),
  .if_cfg_est_m_rd_clk_en(if_cfg_tile2tile_1.rd_clk_en),
  .if_cfg_est_m_rd_en(if_cfg_tile2tile_1.rd_en),
  .if_cfg_est_m_wr_addr(if_cfg_tile2tile_1.wr_addr),
  .if_cfg_est_m_wr_clk_en(if_cfg_tile2tile_1.wr_clk_en),
  .if_cfg_est_m_wr_data(if_cfg_tile2tile_1.wr_data),
  .if_cfg_est_m_wr_en(if_cfg_tile2tile_1.wr_en),
  .if_cfg_wst_s_rd_data(if_cfg_tile2tile_0.rd_data),
  .if_cfg_wst_s_rd_data_valid(if_cfg_tile2tile_0.rd_data_valid),
  .if_proc_est_m_rd_addr(if_proc_tile2tile_1.rd_addr),
  .if_proc_est_m_rd_clk_en(if_proc_tile2tile_1.rd_clk_en),
  .if_proc_est_m_rd_en(if_proc_tile2tile_1.rd_en),
  .if_proc_est_m_wr_addr(if_proc_tile2tile_1.wr_addr),
  .if_proc_est_m_wr_clk_en(if_proc_tile2tile_1.wr_clk_en),
  .if_proc_est_m_wr_data(if_proc_tile2tile_1.wr_data),
  .if_proc_est_m_wr_en(if_proc_tile2tile_1.wr_en),
  .if_proc_est_m_wr_strb(if_proc_tile2tile_1.wr_strb),
  .if_proc_wst_s_rd_data(if_proc_tile2tile_0.rd_data),
  .if_proc_wst_s_rd_data_valid(if_proc_tile2tile_0.rd_data_valid),
  .pcfg_g2f_interrupt_pulse(glb_tile_gen_0_pcfg_g2f_interrupt_pulse),
  .pcfg_rd_addr_e2w_wsto(glb_tile_gen_0_pcfg_rd_addr_e2w_wsto),
  .pcfg_rd_addr_w2e_esto(glb_tile_gen_0_pcfg_rd_addr_w2e_esto),
  .pcfg_rd_data_e2w_wsto(glb_tile_gen_0_pcfg_rd_data_e2w_wsto),
  .pcfg_rd_data_valid_e2w_wsto(glb_tile_gen_0_pcfg_rd_data_valid_e2w_wsto),
  .pcfg_rd_data_valid_w2e_esto(glb_tile_gen_0_pcfg_rd_data_valid_w2e_esto),
  .pcfg_rd_data_w2e_esto(glb_tile_gen_0_pcfg_rd_data_w2e_esto),
  .pcfg_rd_en_e2w_wsto(glb_tile_gen_0_pcfg_rd_en_e2w_wsto),
  .pcfg_rd_en_w2e_esto(glb_tile_gen_0_pcfg_rd_en_w2e_esto),
  .strm_data_g2f(glb_tile_gen_0_strm_data_g2f),
  .strm_data_valid_g2f(glb_tile_gen_0_strm_data_valid_g2f),
  .strm_f2g_interrupt_pulse(glb_tile_gen_0_strm_f2g_interrupt_pulse),
  .strm_g2f_interrupt_pulse(glb_tile_gen_0_strm_g2f_interrupt_pulse),
  .strm_rd_addr_e2w_wsto(glb_tile_gen_0_strm_rd_addr_e2w_wsto),
  .strm_rd_addr_w2e_esto(glb_tile_gen_0_strm_rd_addr_w2e_esto),
  .strm_rd_data_e2w_wsto(glb_tile_gen_0_strm_rd_data_e2w_wsto),
  .strm_rd_data_valid_e2w_wsto(glb_tile_gen_0_strm_rd_data_valid_e2w_wsto),
  .strm_rd_data_valid_w2e_esto(glb_tile_gen_0_strm_rd_data_valid_w2e_esto),
  .strm_rd_data_w2e_esto(glb_tile_gen_0_strm_rd_data_w2e_esto),
  .strm_rd_en_e2w_wsto(glb_tile_gen_0_strm_rd_en_e2w_wsto),
  .strm_rd_en_w2e_esto(glb_tile_gen_0_strm_rd_en_w2e_esto),
  .strm_wr_addr_e2w_wsto(glb_tile_gen_0_strm_wr_addr_e2w_wsto),
  .strm_wr_addr_w2e_esto(glb_tile_gen_0_strm_wr_addr_w2e_esto),
  .strm_wr_data_e2w_wsto(glb_tile_gen_0_strm_wr_data_e2w_wsto),
  .strm_wr_data_w2e_esto(glb_tile_gen_0_strm_wr_data_w2e_esto),
  .strm_wr_en_e2w_wsto(glb_tile_gen_0_strm_wr_en_e2w_wsto),
  .strm_wr_en_w2e_esto(glb_tile_gen_0_strm_wr_en_w2e_esto),
  .strm_wr_strb_e2w_wsto(glb_tile_gen_0_strm_wr_strb_e2w_wsto),
  .strm_wr_strb_w2e_esto(glb_tile_gen_0_strm_wr_strb_w2e_esto)
);

glb_tile glb_tile_gen_1 (
  .cfg_pcfg_tile_connected_wsti(cfg_pcfg_tile_connected[1]),
  .cfg_tile_connected_wsti(cfg_tile_connected[1]),
  .cgra_cfg_jtag_addr_bypass_wsti(cgra_cfg_jtag_addr_bypass_wsti[1]),
  .cgra_cfg_jtag_addr_wsti(cgra_cfg_jtag_addr_wsti[1]),
  .cgra_cfg_jtag_data_wsti(cgra_cfg_jtag_data_wsti[1]),
  .cgra_cfg_jtag_rd_en_bypass_wsti(cgra_cfg_jtag_rd_en_bypass_wsti[1]),
  .cgra_cfg_jtag_rd_en_wsti(cgra_cfg_jtag_rd_en_wsti[1]),
  .cgra_cfg_jtag_wr_en_wsti(cgra_cfg_jtag_wr_en_wsti[1]),
  .cgra_cfg_pcfg_addr_e2w_esti(cgra_cfg_pcfg_addr_esti[1]),
  .cgra_cfg_pcfg_addr_w2e_wsti(cgra_cfg_pcfg_addr_wsti[1]),
  .cgra_cfg_pcfg_data_e2w_esti(cgra_cfg_pcfg_data_esti[1]),
  .cgra_cfg_pcfg_data_w2e_wsti(cgra_cfg_pcfg_data_wsti[1]),
  .cgra_cfg_pcfg_rd_en_e2w_esti(cgra_cfg_pcfg_rd_en_esti[1]),
  .cgra_cfg_pcfg_rd_en_w2e_wsti(cgra_cfg_pcfg_rd_en_wsti[1]),
  .cgra_cfg_pcfg_wr_en_e2w_esti(cgra_cfg_pcfg_wr_en_esti[1]),
  .cgra_cfg_pcfg_wr_en_w2e_wsti(cgra_cfg_pcfg_wr_en_wsti[1]),
  .clk(clk),
  .clk_en_bank_master(glb_tile_gen_1_clk_en_bank_master),
  .clk_en_master(glb_tile_gen_1_clk_en_master),
  .clk_en_pcfg_broadcast(glb_tile_gen_1_clk_en_pcfg_broadcast),
  .glb_tile_id(1'h1),
  .if_cfg_est_m_rd_data(32'h0),
  .if_cfg_est_m_rd_data_valid(1'h0),
  .if_cfg_wst_s_rd_addr(if_cfg_tile2tile_1.rd_addr),
  .if_cfg_wst_s_rd_clk_en(if_cfg_tile2tile_1.rd_clk_en),
  .if_cfg_wst_s_rd_en(if_cfg_tile2tile_1.rd_en),
  .if_cfg_wst_s_wr_addr(if_cfg_tile2tile_1.wr_addr),
  .if_cfg_wst_s_wr_clk_en(if_cfg_tile2tile_1.wr_clk_en),
  .if_cfg_wst_s_wr_data(if_cfg_tile2tile_1.wr_data),
  .if_cfg_wst_s_wr_en(if_cfg_tile2tile_1.wr_en),
  .if_proc_est_m_rd_data(64'h0),
  .if_proc_est_m_rd_data_valid(1'h0),
  .if_proc_wst_s_rd_addr(if_proc_tile2tile_1.rd_addr),
  .if_proc_wst_s_rd_clk_en(if_proc_tile2tile_1.rd_clk_en),
  .if_proc_wst_s_rd_en(if_proc_tile2tile_1.rd_en),
  .if_proc_wst_s_wr_addr(if_proc_tile2tile_1.wr_addr),
  .if_proc_wst_s_wr_clk_en(if_proc_tile2tile_1.wr_clk_en),
  .if_proc_wst_s_wr_data(if_proc_tile2tile_1.wr_data),
  .if_proc_wst_s_wr_en(if_proc_tile2tile_1.wr_en),
  .if_proc_wst_s_wr_strb(if_proc_tile2tile_1.wr_strb),
  .pcfg_rd_addr_e2w_esti(pcfg_packet_e2w_esti[1].rdrq.rd_addr),
  .pcfg_rd_addr_w2e_wsti(pcfg_packet_w2e_wsti[1].rdrq.rd_addr),
  .pcfg_rd_data_e2w_esti(pcfg_packet_e2w_esti[1].rdrs.rd_data),
  .pcfg_rd_data_valid_e2w_esti(pcfg_packet_e2w_esti[1].rdrs.rd_data_valid),
  .pcfg_rd_data_valid_w2e_wsti(pcfg_packet_w2e_wsti[1].rdrs.rd_data_valid),
  .pcfg_rd_data_w2e_wsti(pcfg_packet_w2e_wsti[1].rdrs.rd_data),
  .pcfg_rd_en_e2w_esti(pcfg_packet_e2w_esti[1].rdrq.rd_en),
  .pcfg_rd_en_w2e_wsti(pcfg_packet_w2e_wsti[1].rdrq.rd_en),
  .pcfg_start_pulse(pcfg_start_pulse[1]),
  .reset(reset),
  .strm_data_f2g(strm_data_f2g[1]),
  .strm_data_valid_f2g(strm_data_valid_f2g[1]),
  .strm_f2g_start_pulse(strm_f2g_start_pulse[1]),
  .strm_g2f_start_pulse(strm_g2f_start_pulse[1]),
  .strm_rd_addr_e2w_esti(strm_packet_e2w_esti[1].rdrq.rd_addr),
  .strm_rd_addr_w2e_wsti(strm_packet_w2e_wsti[1].rdrq.rd_addr),
  .strm_rd_data_e2w_esti(strm_packet_e2w_esti[1].rdrs.rd_data),
  .strm_rd_data_valid_e2w_esti(strm_packet_e2w_esti[1].rdrs.rd_data_valid),
  .strm_rd_data_valid_w2e_wsti(strm_packet_w2e_wsti[1].rdrs.rd_data_valid),
  .strm_rd_data_w2e_wsti(strm_packet_w2e_wsti[1].rdrs.rd_data),
  .strm_rd_en_e2w_esti(strm_packet_e2w_esti[1].rdrq.rd_en),
  .strm_rd_en_w2e_wsti(strm_packet_w2e_wsti[1].rdrq.rd_en),
  .strm_wr_addr_e2w_esti(strm_packet_e2w_esti[1].wr.wr_addr),
  .strm_wr_addr_w2e_wsti(strm_packet_w2e_wsti[1].wr.wr_addr),
  .strm_wr_data_e2w_esti(strm_packet_e2w_esti[1].wr.wr_data),
  .strm_wr_data_w2e_wsti(strm_packet_w2e_wsti[1].wr.wr_data),
  .strm_wr_en_e2w_esti(strm_packet_e2w_esti[1].wr.wr_en),
  .strm_wr_en_w2e_wsti(strm_packet_w2e_wsti[1].wr.wr_en),
  .strm_wr_strb_e2w_esti(strm_packet_e2w_esti[1].wr.wr_strb),
  .strm_wr_strb_w2e_wsti(strm_packet_w2e_wsti[1].wr.wr_strb),
  .cfg_pcfg_tile_connected_esto(glb_tile_gen_1_cfg_pcfg_tile_connected_esto),
  .cfg_tile_connected_esto(glb_tile_gen_1_cfg_tile_connected_esto),
  .cgra_cfg_g2f_cfg_addr(glb_tile_gen_1_cgra_cfg_g2f_cfg_addr),
  .cgra_cfg_g2f_cfg_data(glb_tile_gen_1_cgra_cfg_g2f_cfg_data),
  .cgra_cfg_g2f_cfg_rd_en(glb_tile_gen_1_cgra_cfg_g2f_cfg_rd_en),
  .cgra_cfg_g2f_cfg_wr_en(glb_tile_gen_1_cgra_cfg_g2f_cfg_wr_en),
  .cgra_cfg_jtag_addr_bypass_esto(glb_tile_gen_1_cgra_cfg_jtag_addr_bypass_esto),
  .cgra_cfg_jtag_addr_esto(glb_tile_gen_1_cgra_cfg_jtag_addr_esto),
  .cgra_cfg_jtag_data_esto(glb_tile_gen_1_cgra_cfg_jtag_data_esto),
  .cgra_cfg_jtag_rd_en_bypass_esto(glb_tile_gen_1_cgra_cfg_jtag_rd_en_bypass_esto),
  .cgra_cfg_jtag_rd_en_esto(glb_tile_gen_1_cgra_cfg_jtag_rd_en_esto),
  .cgra_cfg_jtag_wr_en_esto(glb_tile_gen_1_cgra_cfg_jtag_wr_en_esto),
  .cgra_cfg_pcfg_addr_e2w_wsto(glb_tile_gen_1_cgra_cfg_pcfg_addr_e2w_wsto),
  .cgra_cfg_pcfg_addr_w2e_esto(glb_tile_gen_1_cgra_cfg_pcfg_addr_w2e_esto),
  .cgra_cfg_pcfg_data_e2w_wsto(glb_tile_gen_1_cgra_cfg_pcfg_data_e2w_wsto),
  .cgra_cfg_pcfg_data_w2e_esto(glb_tile_gen_1_cgra_cfg_pcfg_data_w2e_esto),
  .cgra_cfg_pcfg_rd_en_e2w_wsto(glb_tile_gen_1_cgra_cfg_pcfg_rd_en_e2w_wsto),
  .cgra_cfg_pcfg_rd_en_w2e_esto(glb_tile_gen_1_cgra_cfg_pcfg_rd_en_w2e_esto),
  .cgra_cfg_pcfg_wr_en_e2w_wsto(glb_tile_gen_1_cgra_cfg_pcfg_wr_en_e2w_wsto),
  .cgra_cfg_pcfg_wr_en_w2e_esto(glb_tile_gen_1_cgra_cfg_pcfg_wr_en_w2e_esto),
  .data_flush(glb_tile_gen_1_data_flush),
  .if_cfg_est_m_rd_addr(if_cfg_tile2tile_2.rd_addr),
  .if_cfg_est_m_rd_clk_en(if_cfg_tile2tile_2.rd_clk_en),
  .if_cfg_est_m_rd_en(if_cfg_tile2tile_2.rd_en),
  .if_cfg_est_m_wr_addr(if_cfg_tile2tile_2.wr_addr),
  .if_cfg_est_m_wr_clk_en(if_cfg_tile2tile_2.wr_clk_en),
  .if_cfg_est_m_wr_data(if_cfg_tile2tile_2.wr_data),
  .if_cfg_est_m_wr_en(if_cfg_tile2tile_2.wr_en),
  .if_cfg_wst_s_rd_data(if_cfg_tile2tile_1.rd_data),
  .if_cfg_wst_s_rd_data_valid(if_cfg_tile2tile_1.rd_data_valid),
  .if_proc_est_m_rd_addr(if_proc_tile2tile_2.rd_addr),
  .if_proc_est_m_rd_clk_en(if_proc_tile2tile_2.rd_clk_en),
  .if_proc_est_m_rd_en(if_proc_tile2tile_2.rd_en),
  .if_proc_est_m_wr_addr(if_proc_tile2tile_2.wr_addr),
  .if_proc_est_m_wr_clk_en(if_proc_tile2tile_2.wr_clk_en),
  .if_proc_est_m_wr_data(if_proc_tile2tile_2.wr_data),
  .if_proc_est_m_wr_en(if_proc_tile2tile_2.wr_en),
  .if_proc_est_m_wr_strb(if_proc_tile2tile_2.wr_strb),
  .if_proc_wst_s_rd_data(if_proc_tile2tile_1.rd_data),
  .if_proc_wst_s_rd_data_valid(if_proc_tile2tile_1.rd_data_valid),
  .pcfg_g2f_interrupt_pulse(glb_tile_gen_1_pcfg_g2f_interrupt_pulse),
  .pcfg_rd_addr_e2w_wsto(glb_tile_gen_1_pcfg_rd_addr_e2w_wsto),
  .pcfg_rd_addr_w2e_esto(glb_tile_gen_1_pcfg_rd_addr_w2e_esto),
  .pcfg_rd_data_e2w_wsto(glb_tile_gen_1_pcfg_rd_data_e2w_wsto),
  .pcfg_rd_data_valid_e2w_wsto(glb_tile_gen_1_pcfg_rd_data_valid_e2w_wsto),
  .pcfg_rd_data_valid_w2e_esto(glb_tile_gen_1_pcfg_rd_data_valid_w2e_esto),
  .pcfg_rd_data_w2e_esto(glb_tile_gen_1_pcfg_rd_data_w2e_esto),
  .pcfg_rd_en_e2w_wsto(glb_tile_gen_1_pcfg_rd_en_e2w_wsto),
  .pcfg_rd_en_w2e_esto(glb_tile_gen_1_pcfg_rd_en_w2e_esto),
  .strm_data_g2f(glb_tile_gen_1_strm_data_g2f),
  .strm_data_valid_g2f(glb_tile_gen_1_strm_data_valid_g2f),
  .strm_f2g_interrupt_pulse(glb_tile_gen_1_strm_f2g_interrupt_pulse),
  .strm_g2f_interrupt_pulse(glb_tile_gen_1_strm_g2f_interrupt_pulse),
  .strm_rd_addr_e2w_wsto(glb_tile_gen_1_strm_rd_addr_e2w_wsto),
  .strm_rd_addr_w2e_esto(glb_tile_gen_1_strm_rd_addr_w2e_esto),
  .strm_rd_data_e2w_wsto(glb_tile_gen_1_strm_rd_data_e2w_wsto),
  .strm_rd_data_valid_e2w_wsto(glb_tile_gen_1_strm_rd_data_valid_e2w_wsto),
  .strm_rd_data_valid_w2e_esto(glb_tile_gen_1_strm_rd_data_valid_w2e_esto),
  .strm_rd_data_w2e_esto(glb_tile_gen_1_strm_rd_data_w2e_esto),
  .strm_rd_en_e2w_wsto(glb_tile_gen_1_strm_rd_en_e2w_wsto),
  .strm_rd_en_w2e_esto(glb_tile_gen_1_strm_rd_en_w2e_esto),
  .strm_wr_addr_e2w_wsto(glb_tile_gen_1_strm_wr_addr_e2w_wsto),
  .strm_wr_addr_w2e_esto(glb_tile_gen_1_strm_wr_addr_w2e_esto),
  .strm_wr_data_e2w_wsto(glb_tile_gen_1_strm_wr_data_e2w_wsto),
  .strm_wr_data_w2e_esto(glb_tile_gen_1_strm_wr_data_w2e_esto),
  .strm_wr_en_e2w_wsto(glb_tile_gen_1_strm_wr_en_e2w_wsto),
  .strm_wr_en_w2e_esto(glb_tile_gen_1_strm_wr_en_w2e_esto),
  .strm_wr_strb_e2w_wsto(glb_tile_gen_1_strm_wr_strb_e2w_wsto),
  .strm_wr_strb_w2e_esto(glb_tile_gen_1_strm_wr_strb_w2e_esto)
);

glb_clk_en_gen_unq1 proc_wr_clk_en_gen (
  .clk(clk),
  .enable(proc_wr_clk_en_gen_enable),
  .reset(reset),
  .clk_en(proc_wr_clk_en)
);

glb_clk_en_gen_unq2 proc_rd_clk_en_gen (
  .clk(clk),
  .enable(proc_rd_clk_en_gen_enable),
  .reset(reset),
  .clk_en(proc_rd_clk_en)
);

pipeline_w_2_d_1 flush_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(data_flush),
  .reset(reset),
  .out_(data_flush_d)
);

glb_crossbar_I_2_O_1_W_1 flush_crossbar (
  .in_(flush_crossbar_in),
  .sel_(flush_crossbar_sel_w),
  .out_(strm_data_flush_g2f)
);

endmodule   // global_buffer

module global_buffer_W (
  input logic [31:0] cgra_cfg_jtag_gc2glb_addr,
  input logic [31:0] cgra_cfg_jtag_gc2glb_data,
  input logic cgra_cfg_jtag_gc2glb_rd_en,
  input logic cgra_cfg_jtag_gc2glb_wr_en,
  input logic [3:0] cgra_stall_in,
  input logic clk,
  input logic flush_crossbar_sel,
  input logic [1:0] glb_clk_en_bank_master,
  input logic [1:0] glb_clk_en_master,
  input logic [11:0] if_cfg_rd_addr,
  input logic if_cfg_rd_clk_en,
  input logic if_cfg_rd_en,
  input logic [11:0] if_cfg_wr_addr,
  input logic if_cfg_wr_clk_en,
  input logic [31:0] if_cfg_wr_data,
  input logic if_cfg_wr_en,
  input logic [18:0] if_sram_cfg_rd_addr,
  input logic if_sram_cfg_rd_en,
  input logic [18:0] if_sram_cfg_wr_addr,
  input logic [31:0] if_sram_cfg_wr_data,
  input logic if_sram_cfg_wr_en,
  input logic [1:0] pcfg_broadcast_stall,
  input logic [1:0] pcfg_start_pulse,
  input logic [18:0] proc_rd_addr,
  input logic proc_rd_en,
  input logic [18:0] proc_wr_addr,
  input logic [63:0] proc_wr_data,
  input logic proc_wr_en,
  input logic [7:0] proc_wr_strb,
  input logic reset,
  input logic [15:0] strm_data_f2g_0_0,
  input logic [15:0] strm_data_f2g_0_1,
  input logic [15:0] strm_data_f2g_1_0,
  input logic [15:0] strm_data_f2g_1_1,
  input logic strm_data_valid_f2g_0_0,
  input logic strm_data_valid_f2g_0_1,
  input logic strm_data_valid_f2g_1_0,
  input logic strm_data_valid_f2g_1_1,
  input logic [1:0] strm_f2g_start_pulse,
  input logic [1:0] strm_g2f_start_pulse,
  output logic [31:0] cgra_cfg_g2f_cfg_addr_0_0,
  output logic [31:0] cgra_cfg_g2f_cfg_addr_0_1,
  output logic [31:0] cgra_cfg_g2f_cfg_addr_1_0,
  output logic [31:0] cgra_cfg_g2f_cfg_addr_1_1,
  output logic [31:0] cgra_cfg_g2f_cfg_data_0_0,
  output logic [31:0] cgra_cfg_g2f_cfg_data_0_1,
  output logic [31:0] cgra_cfg_g2f_cfg_data_1_0,
  output logic [31:0] cgra_cfg_g2f_cfg_data_1_1,
  output logic cgra_cfg_g2f_cfg_rd_en_0_0,
  output logic cgra_cfg_g2f_cfg_rd_en_0_1,
  output logic cgra_cfg_g2f_cfg_rd_en_1_0,
  output logic cgra_cfg_g2f_cfg_rd_en_1_1,
  output logic cgra_cfg_g2f_cfg_wr_en_0_0,
  output logic cgra_cfg_g2f_cfg_wr_en_0_1,
  output logic cgra_cfg_g2f_cfg_wr_en_1_0,
  output logic cgra_cfg_g2f_cfg_wr_en_1_1,
  output logic [3:0] cgra_stall,
  output logic [31:0] if_cfg_rd_data,
  output logic if_cfg_rd_data_valid,
  output logic [31:0] if_sram_cfg_rd_data,
  output logic if_sram_cfg_rd_data_valid,
  output logic [1:0] pcfg_g2f_interrupt_pulse,
  output logic [63:0] proc_rd_data,
  output logic proc_rd_data_valid,
  output logic strm_data_flush_g2f,
  output logic [15:0] strm_data_g2f_0_0,
  output logic [15:0] strm_data_g2f_0_1,
  output logic [15:0] strm_data_g2f_1_0,
  output logic [15:0] strm_data_g2f_1_1,
  output logic strm_data_valid_g2f_0_0,
  output logic strm_data_valid_g2f_0_1,
  output logic strm_data_valid_g2f_1_0,
  output logic strm_data_valid_g2f_1_1,
  output logic [1:0] strm_f2g_interrupt_pulse,
  output logic [1:0] strm_g2f_interrupt_pulse
);

logic [1:0][1:0][31:0] global_buffer_cgra_cfg_g2f_cfg_addr;
logic [1:0][1:0][31:0] global_buffer_cgra_cfg_g2f_cfg_data;
logic [1:0][1:0] global_buffer_cgra_cfg_g2f_cfg_rd_en;
logic [1:0][1:0] global_buffer_cgra_cfg_g2f_cfg_wr_en;
logic [1:0][1:0][15:0] global_buffer_strm_data_f2g;
logic [1:0][1:0][15:0] global_buffer_strm_data_g2f;
logic [1:0][1:0] global_buffer_strm_data_valid_f2g;
logic [1:0][1:0] global_buffer_strm_data_valid_g2f;
assign cgra_cfg_g2f_cfg_addr_0_0 = global_buffer_cgra_cfg_g2f_cfg_addr[0][0];
assign cgra_cfg_g2f_cfg_addr_0_1 = global_buffer_cgra_cfg_g2f_cfg_addr[0][1];
assign cgra_cfg_g2f_cfg_addr_1_0 = global_buffer_cgra_cfg_g2f_cfg_addr[1][0];
assign cgra_cfg_g2f_cfg_addr_1_1 = global_buffer_cgra_cfg_g2f_cfg_addr[1][1];
assign cgra_cfg_g2f_cfg_data_0_0 = global_buffer_cgra_cfg_g2f_cfg_data[0][0];
assign cgra_cfg_g2f_cfg_data_0_1 = global_buffer_cgra_cfg_g2f_cfg_data[0][1];
assign cgra_cfg_g2f_cfg_data_1_0 = global_buffer_cgra_cfg_g2f_cfg_data[1][0];
assign cgra_cfg_g2f_cfg_data_1_1 = global_buffer_cgra_cfg_g2f_cfg_data[1][1];
assign cgra_cfg_g2f_cfg_rd_en_0_0 = global_buffer_cgra_cfg_g2f_cfg_rd_en[0][0];
assign cgra_cfg_g2f_cfg_rd_en_0_1 = global_buffer_cgra_cfg_g2f_cfg_rd_en[0][1];
assign cgra_cfg_g2f_cfg_rd_en_1_0 = global_buffer_cgra_cfg_g2f_cfg_rd_en[1][0];
assign cgra_cfg_g2f_cfg_rd_en_1_1 = global_buffer_cgra_cfg_g2f_cfg_rd_en[1][1];
assign cgra_cfg_g2f_cfg_wr_en_0_0 = global_buffer_cgra_cfg_g2f_cfg_wr_en[0][0];
assign cgra_cfg_g2f_cfg_wr_en_0_1 = global_buffer_cgra_cfg_g2f_cfg_wr_en[0][1];
assign cgra_cfg_g2f_cfg_wr_en_1_0 = global_buffer_cgra_cfg_g2f_cfg_wr_en[1][0];
assign cgra_cfg_g2f_cfg_wr_en_1_1 = global_buffer_cgra_cfg_g2f_cfg_wr_en[1][1];
assign global_buffer_strm_data_f2g[0][0] = strm_data_f2g_0_0;
assign global_buffer_strm_data_f2g[0][1] = strm_data_f2g_0_1;
assign global_buffer_strm_data_f2g[1][0] = strm_data_f2g_1_0;
assign global_buffer_strm_data_f2g[1][1] = strm_data_f2g_1_1;
assign strm_data_g2f_0_0 = global_buffer_strm_data_g2f[0][0];
assign strm_data_g2f_0_1 = global_buffer_strm_data_g2f[0][1];
assign strm_data_g2f_1_0 = global_buffer_strm_data_g2f[1][0];
assign strm_data_g2f_1_1 = global_buffer_strm_data_g2f[1][1];
assign global_buffer_strm_data_valid_f2g[0][0] = strm_data_valid_f2g_0_0;
assign global_buffer_strm_data_valid_f2g[0][1] = strm_data_valid_f2g_0_1;
assign global_buffer_strm_data_valid_f2g[1][0] = strm_data_valid_f2g_1_0;
assign global_buffer_strm_data_valid_f2g[1][1] = strm_data_valid_f2g_1_1;
assign strm_data_valid_g2f_0_0 = global_buffer_strm_data_valid_g2f[0][0];
assign strm_data_valid_g2f_0_1 = global_buffer_strm_data_valid_g2f[0][1];
assign strm_data_valid_g2f_1_0 = global_buffer_strm_data_valid_g2f[1][0];
assign strm_data_valid_g2f_1_1 = global_buffer_strm_data_valid_g2f[1][1];
global_buffer global_buffer (
  .cgra_cfg_jtag_gc2glb_addr(cgra_cfg_jtag_gc2glb_addr),
  .cgra_cfg_jtag_gc2glb_data(cgra_cfg_jtag_gc2glb_data),
  .cgra_cfg_jtag_gc2glb_rd_en(cgra_cfg_jtag_gc2glb_rd_en),
  .cgra_cfg_jtag_gc2glb_wr_en(cgra_cfg_jtag_gc2glb_wr_en),
  .cgra_stall_in(cgra_stall_in),
  .clk(clk),
  .flush_crossbar_sel(flush_crossbar_sel),
  .glb_clk_en_bank_master(glb_clk_en_bank_master),
  .glb_clk_en_master(glb_clk_en_master),
  .if_cfg_rd_addr(if_cfg_rd_addr),
  .if_cfg_rd_clk_en(if_cfg_rd_clk_en),
  .if_cfg_rd_en(if_cfg_rd_en),
  .if_cfg_wr_addr(if_cfg_wr_addr),
  .if_cfg_wr_clk_en(if_cfg_wr_clk_en),
  .if_cfg_wr_data(if_cfg_wr_data),
  .if_cfg_wr_en(if_cfg_wr_en),
  .if_sram_cfg_rd_addr(if_sram_cfg_rd_addr),
  .if_sram_cfg_rd_en(if_sram_cfg_rd_en),
  .if_sram_cfg_wr_addr(if_sram_cfg_wr_addr),
  .if_sram_cfg_wr_data(if_sram_cfg_wr_data),
  .if_sram_cfg_wr_en(if_sram_cfg_wr_en),
  .pcfg_broadcast_stall(pcfg_broadcast_stall),
  .pcfg_start_pulse(pcfg_start_pulse),
  .proc_rd_addr(proc_rd_addr),
  .proc_rd_en(proc_rd_en),
  .proc_wr_addr(proc_wr_addr),
  .proc_wr_data(proc_wr_data),
  .proc_wr_en(proc_wr_en),
  .proc_wr_strb(proc_wr_strb),
  .reset(reset),
  .strm_data_f2g(global_buffer_strm_data_f2g),
  .strm_data_valid_f2g(global_buffer_strm_data_valid_f2g),
  .strm_f2g_start_pulse(strm_f2g_start_pulse),
  .strm_g2f_start_pulse(strm_g2f_start_pulse),
  .cgra_cfg_g2f_cfg_addr(global_buffer_cgra_cfg_g2f_cfg_addr),
  .cgra_cfg_g2f_cfg_data(global_buffer_cgra_cfg_g2f_cfg_data),
  .cgra_cfg_g2f_cfg_rd_en(global_buffer_cgra_cfg_g2f_cfg_rd_en),
  .cgra_cfg_g2f_cfg_wr_en(global_buffer_cgra_cfg_g2f_cfg_wr_en),
  .cgra_stall(cgra_stall),
  .if_cfg_rd_data(if_cfg_rd_data),
  .if_cfg_rd_data_valid(if_cfg_rd_data_valid),
  .if_sram_cfg_rd_data(if_sram_cfg_rd_data),
  .if_sram_cfg_rd_data_valid(if_sram_cfg_rd_data_valid),
  .pcfg_g2f_interrupt_pulse(pcfg_g2f_interrupt_pulse),
  .proc_rd_data(proc_rd_data),
  .proc_rd_data_valid(proc_rd_data_valid),
  .strm_data_flush_g2f(strm_data_flush_g2f),
  .strm_data_g2f(global_buffer_strm_data_g2f),
  .strm_data_valid_g2f(global_buffer_strm_data_valid_g2f),
  .strm_f2g_interrupt_pulse(strm_f2g_interrupt_pulse),
  .strm_g2f_interrupt_pulse(strm_g2f_interrupt_pulse)
);

endmodule   // global_buffer_W

module pipeline_w_144_d_0 (
  input logic clk,
  input logic clk_en,
  input logic [143:0] in_,
  input logic reset,
  output logic [143:0] out_
);

assign out_ = in_;
endmodule   // pipeline_w_144_d_0

module pipeline_w_18_d_0 (
  input logic clk,
  input logic clk_en,
  input logic [17:0] in_,
  input logic reset,
  output logic [17:0] out_
);

assign out_ = in_;
endmodule   // pipeline_w_18_d_0

module pipeline_w_1_d_1 (
  input logic clk,
  input logic clk_en,
  input logic in_,
  input logic reset,
  output logic out_
);

logic pipeline_r;
assign out_ = pipeline_r;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    pipeline_r <= 1'h0;
  end
  else if (clk_en) begin
    pipeline_r <= in_;
  end
end
endmodule   // pipeline_w_1_d_1

module pipeline_w_1_d_10_array (
  input logic clk,
  input logic clk_en,
  input logic in_,
  input logic reset,
  output logic out_ [9:0]
);

logic pipeline_r [9:0];
assign out_ = pipeline_r;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    pipeline_r[0] <= 1'h0;
    pipeline_r[1] <= 1'h0;
    pipeline_r[2] <= 1'h0;
    pipeline_r[3] <= 1'h0;
    pipeline_r[4] <= 1'h0;
    pipeline_r[5] <= 1'h0;
    pipeline_r[6] <= 1'h0;
    pipeline_r[7] <= 1'h0;
    pipeline_r[8] <= 1'h0;
    pipeline_r[9] <= 1'h0;
  end
  else if (clk_en) begin
    pipeline_r[0] <= in_;
    pipeline_r[1] <= pipeline_r[4'h0];
    pipeline_r[2] <= pipeline_r[4'h1];
    pipeline_r[3] <= pipeline_r[4'h2];
    pipeline_r[4] <= pipeline_r[4'h3];
    pipeline_r[5] <= pipeline_r[4'h4];
    pipeline_r[6] <= pipeline_r[4'h5];
    pipeline_r[7] <= pipeline_r[4'h6];
    pipeline_r[8] <= pipeline_r[4'h7];
    pipeline_r[9] <= pipeline_r[4'h8];
  end
end
endmodule   // pipeline_w_1_d_10_array

module pipeline_w_1_d_11_array (
  input logic clk,
  input logic clk_en,
  input logic in_,
  input logic reset,
  output logic out_ [10:0]
);

logic pipeline_r [10:0];
assign out_ = pipeline_r;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    pipeline_r[0] <= 1'h0;
    pipeline_r[1] <= 1'h0;
    pipeline_r[2] <= 1'h0;
    pipeline_r[3] <= 1'h0;
    pipeline_r[4] <= 1'h0;
    pipeline_r[5] <= 1'h0;
    pipeline_r[6] <= 1'h0;
    pipeline_r[7] <= 1'h0;
    pipeline_r[8] <= 1'h0;
    pipeline_r[9] <= 1'h0;
    pipeline_r[10] <= 1'h0;
  end
  else if (clk_en) begin
    pipeline_r[0] <= in_;
    pipeline_r[1] <= pipeline_r[4'h0];
    pipeline_r[2] <= pipeline_r[4'h1];
    pipeline_r[3] <= pipeline_r[4'h2];
    pipeline_r[4] <= pipeline_r[4'h3];
    pipeline_r[5] <= pipeline_r[4'h4];
    pipeline_r[6] <= pipeline_r[4'h5];
    pipeline_r[7] <= pipeline_r[4'h6];
    pipeline_r[8] <= pipeline_r[4'h7];
    pipeline_r[9] <= pipeline_r[4'h8];
    pipeline_r[10] <= pipeline_r[4'h9];
  end
end
endmodule   // pipeline_w_1_d_11_array

module pipeline_w_1_d_12_array (
  input logic clk,
  input logic clk_en,
  input logic in_,
  input logic reset,
  output logic out_ [11:0]
);

logic pipeline_r [11:0];
assign out_ = pipeline_r;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    pipeline_r[0] <= 1'h0;
    pipeline_r[1] <= 1'h0;
    pipeline_r[2] <= 1'h0;
    pipeline_r[3] <= 1'h0;
    pipeline_r[4] <= 1'h0;
    pipeline_r[5] <= 1'h0;
    pipeline_r[6] <= 1'h0;
    pipeline_r[7] <= 1'h0;
    pipeline_r[8] <= 1'h0;
    pipeline_r[9] <= 1'h0;
    pipeline_r[10] <= 1'h0;
    pipeline_r[11] <= 1'h0;
  end
  else if (clk_en) begin
    pipeline_r[0] <= in_;
    pipeline_r[1] <= pipeline_r[4'h0];
    pipeline_r[2] <= pipeline_r[4'h1];
    pipeline_r[3] <= pipeline_r[4'h2];
    pipeline_r[4] <= pipeline_r[4'h3];
    pipeline_r[5] <= pipeline_r[4'h4];
    pipeline_r[6] <= pipeline_r[4'h5];
    pipeline_r[7] <= pipeline_r[4'h6];
    pipeline_r[8] <= pipeline_r[4'h7];
    pipeline_r[9] <= pipeline_r[4'h8];
    pipeline_r[10] <= pipeline_r[4'h9];
    pipeline_r[11] <= pipeline_r[4'hA];
  end
end
endmodule   // pipeline_w_1_d_12_array

module pipeline_w_1_d_5 (
  input logic clk,
  input logic clk_en,
  input logic in_,
  input logic reset,
  output logic out_
);

logic pipeline_r [4:0];
assign out_ = pipeline_r[4];

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    pipeline_r[0] <= 1'h0;
    pipeline_r[1] <= 1'h0;
    pipeline_r[2] <= 1'h0;
    pipeline_r[3] <= 1'h0;
    pipeline_r[4] <= 1'h0;
  end
  else if (clk_en) begin
    pipeline_r[0] <= in_;
    pipeline_r[1] <= pipeline_r[3'h0];
    pipeline_r[2] <= pipeline_r[3'h1];
    pipeline_r[3] <= pipeline_r[3'h2];
    pipeline_r[4] <= pipeline_r[3'h3];
  end
end
endmodule   // pipeline_w_1_d_5

module pipeline_w_1_d_8_array (
  input logic clk,
  input logic clk_en,
  input logic in_,
  input logic reset,
  output logic out_ [7:0]
);

logic pipeline_r [7:0];
assign out_ = pipeline_r;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    pipeline_r[0] <= 1'h0;
    pipeline_r[1] <= 1'h0;
    pipeline_r[2] <= 1'h0;
    pipeline_r[3] <= 1'h0;
    pipeline_r[4] <= 1'h0;
    pipeline_r[5] <= 1'h0;
    pipeline_r[6] <= 1'h0;
    pipeline_r[7] <= 1'h0;
  end
  else if (clk_en) begin
    pipeline_r[0] <= in_;
    pipeline_r[1] <= pipeline_r[3'h0];
    pipeline_r[2] <= pipeline_r[3'h1];
    pipeline_r[3] <= pipeline_r[3'h2];
    pipeline_r[4] <= pipeline_r[3'h3];
    pipeline_r[5] <= pipeline_r[3'h4];
    pipeline_r[6] <= pipeline_r[3'h5];
    pipeline_r[7] <= pipeline_r[3'h6];
  end
end
endmodule   // pipeline_w_1_d_8_array

module pipeline_w_2_d_1 (
  input logic clk,
  input logic clk_en,
  input logic [1:0] in_,
  input logic reset,
  output logic [1:0] out_
);

logic [1:0] pipeline_r [0:0];
assign out_ = pipeline_r[0];

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    for (int unsigned i = 0; i < 1; i += 1) begin
        pipeline_r[1'(i)] <= 2'h0;
      end
  end
  else if (clk_en) begin
    for (int unsigned i = 0; i < 1; i += 1) begin
        if (i == 32'h0) begin
          pipeline_r[1'(i)] <= in_;
        end
        else pipeline_r[1'(i)] <= pipeline_r[1'(i - 32'h1)];
      end
  end
end
endmodule   // pipeline_w_2_d_1

module pipeline_w_2_d_10_array (
  input logic clk,
  input logic clk_en,
  input logic [1:0] in_,
  input logic reset,
  output logic [1:0] out_ [9:0]
);

logic [1:0] pipeline_r [9:0];
assign out_ = pipeline_r;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    for (int unsigned i = 0; i < 10; i += 1) begin
        pipeline_r[4'(i)] <= 2'h0;
      end
  end
  else if (clk_en) begin
    for (int unsigned i = 0; i < 10; i += 1) begin
        if (i == 32'h0) begin
          pipeline_r[4'(i)] <= in_;
        end
        else pipeline_r[4'(i)] <= pipeline_r[4'(i - 32'h1)];
      end
  end
end
endmodule   // pipeline_w_2_d_10_array

module pipeline_w_4_d_2 (
  input logic clk,
  input logic clk_en,
  input logic [3:0] in_,
  input logic reset,
  output logic [3:0] out_
);

logic [3:0] pipeline_r [1:0];
assign out_ = pipeline_r[1];

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    for (int unsigned i = 0; i < 2; i += 1) begin
        pipeline_r[1'(i)] <= 4'h0;
      end
  end
  else if (clk_en) begin
    for (int unsigned i = 0; i < 2; i += 1) begin
        if (i == 32'h0) begin
          pipeline_r[1'(i)] <= in_;
        end
        else pipeline_r[1'(i)] <= pipeline_r[1'(i - 32'h1)];
      end
  end
end
endmodule   // pipeline_w_4_d_2

module pipeline_w_64_d_0 (
  input logic clk,
  input logic clk_en,
  input logic [63:0] in_,
  input logic reset,
  output logic [63:0] out_
);

assign out_ = in_;
endmodule   // pipeline_w_64_d_0

module pipeline_w_65_d_1 (
  input logic clk,
  input logic clk_en,
  input logic [64:0] in_,
  input logic reset,
  output logic [64:0] out_
);

logic [64:0] pipeline_r [0:0];
assign out_ = pipeline_r[0];

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    for (int unsigned i = 0; i < 1; i += 1) begin
        pipeline_r[1'(i)] <= 65'h0;
      end
  end
  else if (clk_en) begin
    for (int unsigned i = 0; i < 1; i += 1) begin
        if (i == 32'h0) begin
          pipeline_r[1'(i)] <= in_;
        end
        else pipeline_r[1'(i)] <= pipeline_r[1'(i - 32'h1)];
      end
  end
end
endmodule   // pipeline_w_65_d_1

module pipeline_w_74_d_0_reset_high (
  input logic clk,
  input logic clk_en,
  input logic [73:0] in_,
  input logic reset,
  output logic [73:0] out_
);

assign out_ = in_;
endmodule   // pipeline_w_74_d_0_reset_high

module pipeline_w_78_d_0 (
  input logic clk,
  input logic clk_en,
  input logic [77:0] in_,
  input logic reset,
  output logic [77:0] out_
);

assign out_ = in_;
endmodule   // pipeline_w_78_d_0

module pipeline_w_90_d_0 (
  input logic clk,
  input logic clk_en,
  input logic [89:0] in_,
  input logic reset,
  output logic [89:0] out_
);

assign out_ = in_;
endmodule   // pipeline_w_90_d_0


module flush_mux_sel_unq1 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[0:0];
endmodule

module flush_mux_sel (
    input [23:0] I,
    output [0:0] O
);
assign O = I[0:0];
endmodule

module coreir_wrap (
    input in,
    output out
);
  assign out = in;
endmodule

module coreir_ult #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = in0 < in1;
endmodule

module coreir_ule #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = in0 <= in1;
endmodule

module coreir_uge #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = in0 >= in1;
endmodule

module coreir_slice #(
    parameter hi = 1,
    parameter lo = 0,
    parameter width = 1
) (
    input [width-1:0] in,
    output [hi-lo-1:0] out
);
  assign out = in[hi-1:lo];
endmodule

module coreir_sle #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = $signed(in0) <= $signed(in1);
endmodule

module coreir_sgt #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = $signed(in0) > $signed(in1);
endmodule

module coreir_sge #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = $signed(in0) >= $signed(in1);
endmodule

module coreir_orr #(
    parameter width = 1
) (
    input [width-1:0] in,
    output out
);
  assign out = |in;
endmodule

module coreir_or #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 | in1;
endmodule

module coreir_not #(
    parameter width = 1
) (
    input [width-1:0] in,
    output [width-1:0] out
);
  assign out = ~in;
endmodule

module coreir_neg #(
    parameter width = 1
) (
    input [width-1:0] in,
    output [width-1:0] out
);
  assign out = -in;
endmodule

module coreir_mux #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    input sel,
    output [width-1:0] out
);
  assign out = sel ? in1 : in0;
endmodule

module coreir_mul #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 * in1;
endmodule

module coreir_lshr #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 >> in1;
endmodule

module coreir_eq #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = in0 == in1;
endmodule

module coreir_const #(
    parameter width = 1,
    parameter value = 1
) (
    output [width-1:0] out
);
  assign out = value;
endmodule

module coreir_ashr #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = $signed(in0) >>> in1;
endmodule

module coreir_and #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 & in1;
endmodule

module coreir_add #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 + in1;
endmodule

module corebit_xor (
    input in0,
    input in1,
    output out
);
  assign out = in0 ^ in1;
endmodule

module corebit_term (
    input in
);

endmodule

module corebit_or (
    input in0,
    input in1,
    output out
);
  assign out = in0 | in1;
endmodule

module corebit_not (
    input in,
    output out
);
  assign out = ~in;
endmodule

module corebit_const #(
    parameter value = 1
) (
    output out
);
  assign out = value;
endmodule

module corebit_and (
    input in0,
    input in1,
    output out
);
  assign out = in0 & in1;
endmodule

module commonlib_muxn__N2__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [0:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(in_data_0),
    .in1(in_data_1),
    .sel(in_sel[0]),
    .out(_join_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N4__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_2,
    input [31:0] in_data_3,
    input [1:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [0:0] sel_slice0_out;
wire [0:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[1]),
    .out(_join_out)
);
commonlib_muxn__N2__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N2__width32 muxN_1 (
    .in_data_0(in_data_2),
    .in_data_1(in_data_3),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(1),
    .lo(0),
    .width(2)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(1),
    .lo(0),
    .width(2)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N8__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_2,
    input [31:0] in_data_3,
    input [31:0] in_data_4,
    input [31:0] in_data_5,
    input [31:0] in_data_6,
    input [31:0] in_data_7,
    input [2:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [1:0] sel_slice0_out;
wire [1:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[2]),
    .out(_join_out)
);
commonlib_muxn__N4__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N4__width32 muxN_1 (
    .in_data_0(in_data_4),
    .in_data_1(in_data_5),
    .in_data_2(in_data_6),
    .in_data_3(in_data_7),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(2),
    .lo(0),
    .width(3)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(2),
    .lo(0),
    .width(3)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N1__width32 (
    input [31:0] in_data_0,
    input [0:0] in_sel,
    output [31:0] out
);
corebit_term term_sel (
    .in(in_sel[0])
);
assign out = in_data_0;
endmodule

module commonlib_muxn__N5__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_2,
    input [31:0] in_data_3,
    input [31:0] in_data_4,
    input [2:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [1:0] sel_slice0_out;
wire [0:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[2]),
    .out(_join_out)
);
commonlib_muxn__N4__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N1__width32 muxN_1 (
    .in_data_0(in_data_4),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(2),
    .lo(0),
    .width(3)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(1),
    .lo(0),
    .width(3)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N3__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_2,
    input [1:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [0:0] sel_slice0_out;
wire [0:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[1]),
    .out(_join_out)
);
commonlib_muxn__N2__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N1__width32 muxN_1 (
    .in_data_0(in_data_2),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(1),
    .lo(0),
    .width(2)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(1),
    .lo(0),
    .width(2)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N7__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_2,
    input [31:0] in_data_3,
    input [31:0] in_data_4,
    input [31:0] in_data_5,
    input [31:0] in_data_6,
    input [2:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [1:0] sel_slice0_out;
wire [1:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[2]),
    .out(_join_out)
);
commonlib_muxn__N4__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N3__width32 muxN_1 (
    .in_data_0(in_data_4),
    .in_data_1(in_data_5),
    .in_data_2(in_data_6),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(2),
    .lo(0),
    .width(3)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(2),
    .lo(0),
    .width(3)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N16__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_10,
    input [31:0] in_data_11,
    input [31:0] in_data_12,
    input [31:0] in_data_13,
    input [31:0] in_data_14,
    input [31:0] in_data_15,
    input [31:0] in_data_2,
    input [31:0] in_data_3,
    input [31:0] in_data_4,
    input [31:0] in_data_5,
    input [31:0] in_data_6,
    input [31:0] in_data_7,
    input [31:0] in_data_8,
    input [31:0] in_data_9,
    input [3:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [2:0] sel_slice0_out;
wire [2:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[3]),
    .out(_join_out)
);
commonlib_muxn__N8__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_data_4(in_data_4),
    .in_data_5(in_data_5),
    .in_data_6(in_data_6),
    .in_data_7(in_data_7),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N8__width32 muxN_1 (
    .in_data_0(in_data_8),
    .in_data_1(in_data_9),
    .in_data_2(in_data_10),
    .in_data_3(in_data_11),
    .in_data_4(in_data_12),
    .in_data_5(in_data_13),
    .in_data_6(in_data_14),
    .in_data_7(in_data_15),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(3),
    .lo(0),
    .width(4)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(3),
    .lo(0),
    .width(4)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N32__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_10,
    input [31:0] in_data_11,
    input [31:0] in_data_12,
    input [31:0] in_data_13,
    input [31:0] in_data_14,
    input [31:0] in_data_15,
    input [31:0] in_data_16,
    input [31:0] in_data_17,
    input [31:0] in_data_18,
    input [31:0] in_data_19,
    input [31:0] in_data_2,
    input [31:0] in_data_20,
    input [31:0] in_data_21,
    input [31:0] in_data_22,
    input [31:0] in_data_23,
    input [31:0] in_data_24,
    input [31:0] in_data_25,
    input [31:0] in_data_26,
    input [31:0] in_data_27,
    input [31:0] in_data_28,
    input [31:0] in_data_29,
    input [31:0] in_data_3,
    input [31:0] in_data_30,
    input [31:0] in_data_31,
    input [31:0] in_data_4,
    input [31:0] in_data_5,
    input [31:0] in_data_6,
    input [31:0] in_data_7,
    input [31:0] in_data_8,
    input [31:0] in_data_9,
    input [4:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [3:0] sel_slice0_out;
wire [3:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[4]),
    .out(_join_out)
);
commonlib_muxn__N16__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_10(in_data_10),
    .in_data_11(in_data_11),
    .in_data_12(in_data_12),
    .in_data_13(in_data_13),
    .in_data_14(in_data_14),
    .in_data_15(in_data_15),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_data_4(in_data_4),
    .in_data_5(in_data_5),
    .in_data_6(in_data_6),
    .in_data_7(in_data_7),
    .in_data_8(in_data_8),
    .in_data_9(in_data_9),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N16__width32 muxN_1 (
    .in_data_0(in_data_16),
    .in_data_1(in_data_17),
    .in_data_10(in_data_26),
    .in_data_11(in_data_27),
    .in_data_12(in_data_28),
    .in_data_13(in_data_29),
    .in_data_14(in_data_30),
    .in_data_15(in_data_31),
    .in_data_2(in_data_18),
    .in_data_3(in_data_19),
    .in_data_4(in_data_20),
    .in_data_5(in_data_21),
    .in_data_6(in_data_22),
    .in_data_7(in_data_23),
    .in_data_8(in_data_24),
    .in_data_9(in_data_25),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(4),
    .lo(0),
    .width(5)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(4),
    .lo(0),
    .width(5)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N64__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_10,
    input [31:0] in_data_11,
    input [31:0] in_data_12,
    input [31:0] in_data_13,
    input [31:0] in_data_14,
    input [31:0] in_data_15,
    input [31:0] in_data_16,
    input [31:0] in_data_17,
    input [31:0] in_data_18,
    input [31:0] in_data_19,
    input [31:0] in_data_2,
    input [31:0] in_data_20,
    input [31:0] in_data_21,
    input [31:0] in_data_22,
    input [31:0] in_data_23,
    input [31:0] in_data_24,
    input [31:0] in_data_25,
    input [31:0] in_data_26,
    input [31:0] in_data_27,
    input [31:0] in_data_28,
    input [31:0] in_data_29,
    input [31:0] in_data_3,
    input [31:0] in_data_30,
    input [31:0] in_data_31,
    input [31:0] in_data_32,
    input [31:0] in_data_33,
    input [31:0] in_data_34,
    input [31:0] in_data_35,
    input [31:0] in_data_36,
    input [31:0] in_data_37,
    input [31:0] in_data_38,
    input [31:0] in_data_39,
    input [31:0] in_data_4,
    input [31:0] in_data_40,
    input [31:0] in_data_41,
    input [31:0] in_data_42,
    input [31:0] in_data_43,
    input [31:0] in_data_44,
    input [31:0] in_data_45,
    input [31:0] in_data_46,
    input [31:0] in_data_47,
    input [31:0] in_data_48,
    input [31:0] in_data_49,
    input [31:0] in_data_5,
    input [31:0] in_data_50,
    input [31:0] in_data_51,
    input [31:0] in_data_52,
    input [31:0] in_data_53,
    input [31:0] in_data_54,
    input [31:0] in_data_55,
    input [31:0] in_data_56,
    input [31:0] in_data_57,
    input [31:0] in_data_58,
    input [31:0] in_data_59,
    input [31:0] in_data_6,
    input [31:0] in_data_60,
    input [31:0] in_data_61,
    input [31:0] in_data_62,
    input [31:0] in_data_63,
    input [31:0] in_data_7,
    input [31:0] in_data_8,
    input [31:0] in_data_9,
    input [5:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [4:0] sel_slice0_out;
wire [4:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[5]),
    .out(_join_out)
);
commonlib_muxn__N32__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_10(in_data_10),
    .in_data_11(in_data_11),
    .in_data_12(in_data_12),
    .in_data_13(in_data_13),
    .in_data_14(in_data_14),
    .in_data_15(in_data_15),
    .in_data_16(in_data_16),
    .in_data_17(in_data_17),
    .in_data_18(in_data_18),
    .in_data_19(in_data_19),
    .in_data_2(in_data_2),
    .in_data_20(in_data_20),
    .in_data_21(in_data_21),
    .in_data_22(in_data_22),
    .in_data_23(in_data_23),
    .in_data_24(in_data_24),
    .in_data_25(in_data_25),
    .in_data_26(in_data_26),
    .in_data_27(in_data_27),
    .in_data_28(in_data_28),
    .in_data_29(in_data_29),
    .in_data_3(in_data_3),
    .in_data_30(in_data_30),
    .in_data_31(in_data_31),
    .in_data_4(in_data_4),
    .in_data_5(in_data_5),
    .in_data_6(in_data_6),
    .in_data_7(in_data_7),
    .in_data_8(in_data_8),
    .in_data_9(in_data_9),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N32__width32 muxN_1 (
    .in_data_0(in_data_32),
    .in_data_1(in_data_33),
    .in_data_10(in_data_42),
    .in_data_11(in_data_43),
    .in_data_12(in_data_44),
    .in_data_13(in_data_45),
    .in_data_14(in_data_46),
    .in_data_15(in_data_47),
    .in_data_16(in_data_48),
    .in_data_17(in_data_49),
    .in_data_18(in_data_50),
    .in_data_19(in_data_51),
    .in_data_2(in_data_34),
    .in_data_20(in_data_52),
    .in_data_21(in_data_53),
    .in_data_22(in_data_54),
    .in_data_23(in_data_55),
    .in_data_24(in_data_56),
    .in_data_25(in_data_57),
    .in_data_26(in_data_58),
    .in_data_27(in_data_59),
    .in_data_28(in_data_60),
    .in_data_29(in_data_61),
    .in_data_3(in_data_35),
    .in_data_30(in_data_62),
    .in_data_31(in_data_63),
    .in_data_4(in_data_36),
    .in_data_5(in_data_37),
    .in_data_6(in_data_38),
    .in_data_7(in_data_39),
    .in_data_8(in_data_40),
    .in_data_9(in_data_41),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(5),
    .lo(0),
    .width(6)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(5),
    .lo(0),
    .width(6)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N20__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_10,
    input [31:0] in_data_11,
    input [31:0] in_data_12,
    input [31:0] in_data_13,
    input [31:0] in_data_14,
    input [31:0] in_data_15,
    input [31:0] in_data_16,
    input [31:0] in_data_17,
    input [31:0] in_data_18,
    input [31:0] in_data_19,
    input [31:0] in_data_2,
    input [31:0] in_data_3,
    input [31:0] in_data_4,
    input [31:0] in_data_5,
    input [31:0] in_data_6,
    input [31:0] in_data_7,
    input [31:0] in_data_8,
    input [31:0] in_data_9,
    input [4:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [3:0] sel_slice0_out;
wire [1:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[4]),
    .out(_join_out)
);
commonlib_muxn__N16__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_10(in_data_10),
    .in_data_11(in_data_11),
    .in_data_12(in_data_12),
    .in_data_13(in_data_13),
    .in_data_14(in_data_14),
    .in_data_15(in_data_15),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_data_4(in_data_4),
    .in_data_5(in_data_5),
    .in_data_6(in_data_6),
    .in_data_7(in_data_7),
    .in_data_8(in_data_8),
    .in_data_9(in_data_9),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N4__width32 muxN_1 (
    .in_data_0(in_data_16),
    .in_data_1(in_data_17),
    .in_data_2(in_data_18),
    .in_data_3(in_data_19),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(4),
    .lo(0),
    .width(5)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(2),
    .lo(0),
    .width(5)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N84__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_10,
    input [31:0] in_data_11,
    input [31:0] in_data_12,
    input [31:0] in_data_13,
    input [31:0] in_data_14,
    input [31:0] in_data_15,
    input [31:0] in_data_16,
    input [31:0] in_data_17,
    input [31:0] in_data_18,
    input [31:0] in_data_19,
    input [31:0] in_data_2,
    input [31:0] in_data_20,
    input [31:0] in_data_21,
    input [31:0] in_data_22,
    input [31:0] in_data_23,
    input [31:0] in_data_24,
    input [31:0] in_data_25,
    input [31:0] in_data_26,
    input [31:0] in_data_27,
    input [31:0] in_data_28,
    input [31:0] in_data_29,
    input [31:0] in_data_3,
    input [31:0] in_data_30,
    input [31:0] in_data_31,
    input [31:0] in_data_32,
    input [31:0] in_data_33,
    input [31:0] in_data_34,
    input [31:0] in_data_35,
    input [31:0] in_data_36,
    input [31:0] in_data_37,
    input [31:0] in_data_38,
    input [31:0] in_data_39,
    input [31:0] in_data_4,
    input [31:0] in_data_40,
    input [31:0] in_data_41,
    input [31:0] in_data_42,
    input [31:0] in_data_43,
    input [31:0] in_data_44,
    input [31:0] in_data_45,
    input [31:0] in_data_46,
    input [31:0] in_data_47,
    input [31:0] in_data_48,
    input [31:0] in_data_49,
    input [31:0] in_data_5,
    input [31:0] in_data_50,
    input [31:0] in_data_51,
    input [31:0] in_data_52,
    input [31:0] in_data_53,
    input [31:0] in_data_54,
    input [31:0] in_data_55,
    input [31:0] in_data_56,
    input [31:0] in_data_57,
    input [31:0] in_data_58,
    input [31:0] in_data_59,
    input [31:0] in_data_6,
    input [31:0] in_data_60,
    input [31:0] in_data_61,
    input [31:0] in_data_62,
    input [31:0] in_data_63,
    input [31:0] in_data_64,
    input [31:0] in_data_65,
    input [31:0] in_data_66,
    input [31:0] in_data_67,
    input [31:0] in_data_68,
    input [31:0] in_data_69,
    input [31:0] in_data_7,
    input [31:0] in_data_70,
    input [31:0] in_data_71,
    input [31:0] in_data_72,
    input [31:0] in_data_73,
    input [31:0] in_data_74,
    input [31:0] in_data_75,
    input [31:0] in_data_76,
    input [31:0] in_data_77,
    input [31:0] in_data_78,
    input [31:0] in_data_79,
    input [31:0] in_data_8,
    input [31:0] in_data_80,
    input [31:0] in_data_81,
    input [31:0] in_data_82,
    input [31:0] in_data_83,
    input [31:0] in_data_9,
    input [6:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [5:0] sel_slice0_out;
wire [4:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[6]),
    .out(_join_out)
);
commonlib_muxn__N64__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_10(in_data_10),
    .in_data_11(in_data_11),
    .in_data_12(in_data_12),
    .in_data_13(in_data_13),
    .in_data_14(in_data_14),
    .in_data_15(in_data_15),
    .in_data_16(in_data_16),
    .in_data_17(in_data_17),
    .in_data_18(in_data_18),
    .in_data_19(in_data_19),
    .in_data_2(in_data_2),
    .in_data_20(in_data_20),
    .in_data_21(in_data_21),
    .in_data_22(in_data_22),
    .in_data_23(in_data_23),
    .in_data_24(in_data_24),
    .in_data_25(in_data_25),
    .in_data_26(in_data_26),
    .in_data_27(in_data_27),
    .in_data_28(in_data_28),
    .in_data_29(in_data_29),
    .in_data_3(in_data_3),
    .in_data_30(in_data_30),
    .in_data_31(in_data_31),
    .in_data_32(in_data_32),
    .in_data_33(in_data_33),
    .in_data_34(in_data_34),
    .in_data_35(in_data_35),
    .in_data_36(in_data_36),
    .in_data_37(in_data_37),
    .in_data_38(in_data_38),
    .in_data_39(in_data_39),
    .in_data_4(in_data_4),
    .in_data_40(in_data_40),
    .in_data_41(in_data_41),
    .in_data_42(in_data_42),
    .in_data_43(in_data_43),
    .in_data_44(in_data_44),
    .in_data_45(in_data_45),
    .in_data_46(in_data_46),
    .in_data_47(in_data_47),
    .in_data_48(in_data_48),
    .in_data_49(in_data_49),
    .in_data_5(in_data_5),
    .in_data_50(in_data_50),
    .in_data_51(in_data_51),
    .in_data_52(in_data_52),
    .in_data_53(in_data_53),
    .in_data_54(in_data_54),
    .in_data_55(in_data_55),
    .in_data_56(in_data_56),
    .in_data_57(in_data_57),
    .in_data_58(in_data_58),
    .in_data_59(in_data_59),
    .in_data_6(in_data_6),
    .in_data_60(in_data_60),
    .in_data_61(in_data_61),
    .in_data_62(in_data_62),
    .in_data_63(in_data_63),
    .in_data_7(in_data_7),
    .in_data_8(in_data_8),
    .in_data_9(in_data_9),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N20__width32 muxN_1 (
    .in_data_0(in_data_64),
    .in_data_1(in_data_65),
    .in_data_10(in_data_74),
    .in_data_11(in_data_75),
    .in_data_12(in_data_76),
    .in_data_13(in_data_77),
    .in_data_14(in_data_78),
    .in_data_15(in_data_79),
    .in_data_16(in_data_80),
    .in_data_17(in_data_81),
    .in_data_18(in_data_82),
    .in_data_19(in_data_83),
    .in_data_2(in_data_66),
    .in_data_3(in_data_67),
    .in_data_4(in_data_68),
    .in_data_5(in_data_69),
    .in_data_6(in_data_70),
    .in_data_7(in_data_71),
    .in_data_8(in_data_72),
    .in_data_9(in_data_73),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(6),
    .lo(0),
    .width(7)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(5),
    .lo(0),
    .width(7)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N15__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_10,
    input [31:0] in_data_11,
    input [31:0] in_data_12,
    input [31:0] in_data_13,
    input [31:0] in_data_14,
    input [31:0] in_data_2,
    input [31:0] in_data_3,
    input [31:0] in_data_4,
    input [31:0] in_data_5,
    input [31:0] in_data_6,
    input [31:0] in_data_7,
    input [31:0] in_data_8,
    input [31:0] in_data_9,
    input [3:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [2:0] sel_slice0_out;
wire [2:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[3]),
    .out(_join_out)
);
commonlib_muxn__N8__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_data_4(in_data_4),
    .in_data_5(in_data_5),
    .in_data_6(in_data_6),
    .in_data_7(in_data_7),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N7__width32 muxN_1 (
    .in_data_0(in_data_8),
    .in_data_1(in_data_9),
    .in_data_2(in_data_10),
    .in_data_3(in_data_11),
    .in_data_4(in_data_12),
    .in_data_5(in_data_13),
    .in_data_6(in_data_14),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(3),
    .lo(0),
    .width(4)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(3),
    .lo(0),
    .width(4)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N13__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_10,
    input [31:0] in_data_11,
    input [31:0] in_data_12,
    input [31:0] in_data_2,
    input [31:0] in_data_3,
    input [31:0] in_data_4,
    input [31:0] in_data_5,
    input [31:0] in_data_6,
    input [31:0] in_data_7,
    input [31:0] in_data_8,
    input [31:0] in_data_9,
    input [3:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [2:0] sel_slice0_out;
wire [2:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[3]),
    .out(_join_out)
);
commonlib_muxn__N8__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_data_4(in_data_4),
    .in_data_5(in_data_5),
    .in_data_6(in_data_6),
    .in_data_7(in_data_7),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N5__width32 muxN_1 (
    .in_data_0(in_data_8),
    .in_data_1(in_data_9),
    .in_data_2(in_data_10),
    .in_data_3(in_data_11),
    .in_data_4(in_data_12),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(3),
    .lo(0),
    .width(4)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(3),
    .lo(0),
    .width(4)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N11__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_10,
    input [31:0] in_data_2,
    input [31:0] in_data_3,
    input [31:0] in_data_4,
    input [31:0] in_data_5,
    input [31:0] in_data_6,
    input [31:0] in_data_7,
    input [31:0] in_data_8,
    input [31:0] in_data_9,
    input [3:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [2:0] sel_slice0_out;
wire [1:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[3]),
    .out(_join_out)
);
commonlib_muxn__N8__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_data_4(in_data_4),
    .in_data_5(in_data_5),
    .in_data_6(in_data_6),
    .in_data_7(in_data_7),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N3__width32 muxN_1 (
    .in_data_0(in_data_8),
    .in_data_1(in_data_9),
    .in_data_2(in_data_10),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(3),
    .lo(0),
    .width(4)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(2),
    .lo(0),
    .width(4)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module SUB (
    input [15:0] a,
    input [15:0] b,
    output [15:0] O0,
    output O1,
    output O2,
    output O3,
    output O4,
    output O5,
    input CLK,
    input ASYNCRESET
);
wire bit_const_0_None_out;
wire [15:0] const_0_16_out;
wire [16:0] const_1_17_out;
wire magma_Bit_and_inst0_out;
wire magma_Bit_and_inst1_out;
wire magma_Bit_and_inst2_out;
wire magma_Bit_and_inst3_out;
wire magma_Bit_not_inst0_out;
wire magma_Bit_not_inst1_out;
wire magma_Bit_not_inst2_out;
wire magma_Bit_or_inst0_out;
wire [15:0] magma_Bits_16_not_inst0_out;
wire magma_UInt_16_eq_inst0_out;
wire [16:0] magma_UInt_17_add_inst0_out;
wire [16:0] magma_UInt_17_add_inst1_out;
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
coreir_const #(
    .value(17'h00001),
    .width(17)
) const_1_17 (
    .out(const_1_17_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(a[15]),
    .in1(magma_Bits_16_not_inst0_out[15]),
    .out(magma_Bit_and_inst0_out)
);
corebit_and magma_Bit_and_inst1 (
    .in0(magma_Bit_and_inst0_out),
    .in1(magma_Bit_not_inst0_out),
    .out(magma_Bit_and_inst1_out)
);
corebit_and magma_Bit_and_inst2 (
    .in0(magma_Bit_not_inst1_out),
    .in1(magma_Bit_not_inst2_out),
    .out(magma_Bit_and_inst2_out)
);
corebit_and magma_Bit_and_inst3 (
    .in0(magma_Bit_and_inst2_out),
    .in1(magma_UInt_17_add_inst1_out[15]),
    .out(magma_Bit_and_inst3_out)
);
corebit_not magma_Bit_not_inst0 (
    .in(magma_UInt_17_add_inst1_out[15]),
    .out(magma_Bit_not_inst0_out)
);
corebit_not magma_Bit_not_inst1 (
    .in(a[15]),
    .out(magma_Bit_not_inst1_out)
);
corebit_not magma_Bit_not_inst2 (
    .in(magma_Bits_16_not_inst0_out[15]),
    .out(magma_Bit_not_inst2_out)
);
corebit_or magma_Bit_or_inst0 (
    .in0(magma_Bit_and_inst1_out),
    .in1(magma_Bit_and_inst3_out),
    .out(magma_Bit_or_inst0_out)
);
coreir_not #(
    .width(16)
) magma_Bits_16_not_inst0 (
    .in(b),
    .out(magma_Bits_16_not_inst0_out)
);
wire [15:0] magma_UInt_16_eq_inst0_in0;
assign magma_UInt_16_eq_inst0_in0 = {magma_UInt_17_add_inst1_out[15],magma_UInt_17_add_inst1_out[14],magma_UInt_17_add_inst1_out[13],magma_UInt_17_add_inst1_out[12],magma_UInt_17_add_inst1_out[11],magma_UInt_17_add_inst1_out[10],magma_UInt_17_add_inst1_out[9],magma_UInt_17_add_inst1_out[8],magma_UInt_17_add_inst1_out[7],magma_UInt_17_add_inst1_out[6],magma_UInt_17_add_inst1_out[5],magma_UInt_17_add_inst1_out[4],magma_UInt_17_add_inst1_out[3],magma_UInt_17_add_inst1_out[2],magma_UInt_17_add_inst1_out[1],magma_UInt_17_add_inst1_out[0]};
coreir_eq #(
    .width(16)
) magma_UInt_16_eq_inst0 (
    .in0(magma_UInt_16_eq_inst0_in0),
    .in1(const_0_16_out),
    .out(magma_UInt_16_eq_inst0_out)
);
wire [16:0] magma_UInt_17_add_inst0_in0;
assign magma_UInt_17_add_inst0_in0 = {bit_const_0_None_out,a};
wire [16:0] magma_UInt_17_add_inst0_in1;
assign magma_UInt_17_add_inst0_in1 = {bit_const_0_None_out,magma_Bits_16_not_inst0_out};
coreir_add #(
    .width(17)
) magma_UInt_17_add_inst0 (
    .in0(magma_UInt_17_add_inst0_in0),
    .in1(magma_UInt_17_add_inst0_in1),
    .out(magma_UInt_17_add_inst0_out)
);
coreir_add #(
    .width(17)
) magma_UInt_17_add_inst1 (
    .in0(magma_UInt_17_add_inst0_out),
    .in1(const_1_17_out),
    .out(magma_UInt_17_add_inst1_out)
);
assign O0 = {magma_UInt_17_add_inst1_out[15],magma_UInt_17_add_inst1_out[14],magma_UInt_17_add_inst1_out[13],magma_UInt_17_add_inst1_out[12],magma_UInt_17_add_inst1_out[11],magma_UInt_17_add_inst1_out[10],magma_UInt_17_add_inst1_out[9],magma_UInt_17_add_inst1_out[8],magma_UInt_17_add_inst1_out[7],magma_UInt_17_add_inst1_out[6],magma_UInt_17_add_inst1_out[5],magma_UInt_17_add_inst1_out[4],magma_UInt_17_add_inst1_out[3],magma_UInt_17_add_inst1_out[2],magma_UInt_17_add_inst1_out[1],magma_UInt_17_add_inst1_out[0]};
assign O1 = magma_UInt_17_add_inst1_out[16];
assign O2 = magma_UInt_16_eq_inst0_out;
assign O3 = magma_UInt_17_add_inst1_out[15];
assign O4 = magma_UInt_17_add_inst1_out[16];
assign O5 = magma_Bit_or_inst0_out;
endmodule

module SHR (
    input [0:0] signed_,
    input [15:0] a,
    input [15:0] b,
    output [15:0] O0,
    output O1,
    output O2,
    output O3,
    output O4,
    output O5,
    input CLK,
    input ASYNCRESET
);
wire [15:0] Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire bit_const_0_None_out;
wire [15:0] const_0_16_out;
wire [0:0] const_1_1_out;
wire magma_Bits_16_eq_inst0_out;
wire magma_Bits_1_eq_inst0_out;
wire [15:0] magma_SInt_16_ashr_inst0_out;
wire [15:0] magma_UInt_16_lshr_inst0_out;
coreir_mux #(
    .width(16)
) Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(magma_UInt_16_lshr_inst0_out),
    .in1(magma_SInt_16_ashr_inst0_out),
    .sel(magma_Bits_1_eq_inst0_out),
    .out(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_eq #(
    .width(16)
) magma_Bits_16_eq_inst0 (
    .in0(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(const_0_16_out),
    .out(magma_Bits_16_eq_inst0_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst0 (
    .in0(signed_),
    .in1(const_1_1_out),
    .out(magma_Bits_1_eq_inst0_out)
);
coreir_ashr #(
    .width(16)
) magma_SInt_16_ashr_inst0 (
    .in0(a),
    .in1(b),
    .out(magma_SInt_16_ashr_inst0_out)
);
coreir_lshr #(
    .width(16)
) magma_UInt_16_lshr_inst0 (
    .in0(a),
    .in1(b),
    .out(magma_UInt_16_lshr_inst0_out)
);
assign O0 = Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign O1 = bit_const_0_None_out;
assign O2 = magma_Bits_16_eq_inst0_out;
assign O3 = Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15];
assign O4 = bit_const_0_None_out;
assign O5 = bit_const_0_None_out;
endmodule

module SB_T4_WEST_SB_OUT_B1_sel (
    input [17:0] I,
    output [2:0] O
);
assign O = I[17:15];
endmodule

module SB_T4_WEST_SB_OUT_B16_sel (
    input [17:0] I,
    output [2:0] O
);
assign O = I[17:15];
endmodule

module SB_T4_SOUTH_SB_OUT_B1_sel (
    input [17:0] I,
    output [2:0] O
);
assign O = I[14:12];
endmodule

module SB_T4_SOUTH_SB_OUT_B16_sel (
    input [17:0] I,
    output [2:0] O
);
assign O = I[14:12];
endmodule

module SB_T4_NORTH_SB_OUT_B1_sel (
    input [17:0] I,
    output [2:0] O
);
assign O = I[11:9];
endmodule

module SB_T4_NORTH_SB_OUT_B16_sel (
    input [17:0] I,
    output [2:0] O
);
assign O = I[11:9];
endmodule

module SB_T4_EAST_SB_OUT_B1_sel (
    input [17:0] I,
    output [2:0] O
);
assign O = I[8:6];
endmodule

module SB_T4_EAST_SB_OUT_B16_sel (
    input [17:0] I,
    output [2:0] O
);
assign O = I[8:6];
endmodule

module SB_T3_WEST_SB_OUT_B1_sel (
    input [17:0] I,
    output [2:0] O
);
assign O = I[5:3];
endmodule

module SB_T3_WEST_SB_OUT_B16_sel (
    input [17:0] I,
    output [2:0] O
);
assign O = I[5:3];
endmodule

module SB_T3_SOUTH_SB_OUT_B1_sel (
    input [17:0] I,
    output [2:0] O
);
assign O = I[2:0];
endmodule

module SB_T3_SOUTH_SB_OUT_B16_sel (
    input [17:0] I,
    output [2:0] O
);
assign O = I[2:0];
endmodule

module SB_T3_NORTH_SB_OUT_B1_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[29:27];
endmodule

module SB_T3_NORTH_SB_OUT_B16_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[29:27];
endmodule

module SB_T3_EAST_SB_OUT_B1_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[26:24];
endmodule

module SB_T3_EAST_SB_OUT_B16_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[26:24];
endmodule

module SB_T2_WEST_SB_OUT_B1_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[23:21];
endmodule

module SB_T2_WEST_SB_OUT_B16_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[23:21];
endmodule

module SB_T2_SOUTH_SB_OUT_B1_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[20:18];
endmodule

module SB_T2_SOUTH_SB_OUT_B16_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[20:18];
endmodule

module SB_T2_NORTH_SB_OUT_B1_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[17:15];
endmodule

module SB_T2_NORTH_SB_OUT_B16_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[17:15];
endmodule

module SB_T2_EAST_SB_OUT_B1_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[14:12];
endmodule

module SB_T2_EAST_SB_OUT_B16_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[14:12];
endmodule

module SB_T1_WEST_SB_OUT_B1_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[11:9];
endmodule

module SB_T1_WEST_SB_OUT_B16_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[11:9];
endmodule

module SB_T1_SOUTH_SB_OUT_B1_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[8:6];
endmodule

module SB_T1_SOUTH_SB_OUT_B16_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[8:6];
endmodule

module SB_T1_NORTH_SB_OUT_B1_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[5:3];
endmodule

module SB_T1_NORTH_SB_OUT_B16_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[5:3];
endmodule

module SB_T1_EAST_SB_OUT_B1_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[2:0];
endmodule

module SB_T1_EAST_SB_OUT_B16_sel (
    input [29:0] I,
    output [2:0] O
);
assign O = I[2:0];
endmodule

module SB_T0_WEST_SB_OUT_B1_sel (
    input [31:0] I,
    output [2:0] O
);
assign O = I[31:29];
endmodule

module SB_T0_WEST_SB_OUT_B16_sel (
    input [31:0] I,
    output [2:0] O
);
assign O = I[31:29];
endmodule

module SB_T0_SOUTH_SB_OUT_B1_sel (
    input [31:0] I,
    output [2:0] O
);
assign O = I[28:26];
endmodule

module SB_T0_SOUTH_SB_OUT_B16_sel (
    input [31:0] I,
    output [2:0] O
);
assign O = I[28:26];
endmodule

module SB_T0_NORTH_SB_OUT_B1_sel (
    input [31:0] I,
    output [2:0] O
);
assign O = I[25:23];
endmodule

module SB_T0_NORTH_SB_OUT_B16_sel (
    input [31:0] I,
    output [2:0] O
);
assign O = I[25:23];
endmodule

module SB_T0_EAST_SB_OUT_B1_sel (
    input [31:0] I,
    output [2:0] O
);
assign O = I[22:20];
endmodule

module SB_T0_EAST_SB_OUT_B16_sel (
    input [31:0] I,
    output [2:0] O
);
assign O = I[22:20];
endmodule

module Register_unq9 (
    input [19:0] I,
    output [19:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [19:0] reg_PR20_inst0__CE_out;
regCE_arst #(
    .init(20'h00000),
    .width(20)
) reg_PR20_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR20_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR20_inst0__CE_out;
endmodule

module Register_unq8 (
    input [24:0] I,
    output [24:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [24:0] reg_PR25_inst0__CE_out;
regCE_arst #(
    .init(25'h0000000),
    .width(25)
) reg_PR25_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR25_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR25_inst0__CE_out;
endmodule

module Register_unq7 (
    input [17:0] I,
    output [17:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [17:0] reg_PR18_inst0__CE_out;
regCE_arst #(
    .init(18'h00000),
    .width(18)
) reg_PR18_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR18_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR18_inst0__CE_out;
endmodule

module Register_unq6 (
    input [29:0] I,
    output [29:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [29:0] reg_PR30_inst0__CE_out;
regCE_arst #(
    .init(30'h00000000),
    .width(30)
) reg_PR30_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR30_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR30_inst0__CE_out;
endmodule

module Register_unq5 (
    input [0:0] I,
    output [0:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [0:0] reg_PR1_inst0__CE_out;
regCE_arst #(
    .init(1'h0),
    .width(1)
) reg_PR1_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR1_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR1_inst0__CE_out;
endmodule

module Register_unq4 (
    input [22:0] I,
    output [22:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [22:0] reg_PR23_inst0__CE_out;
regCE_arst #(
    .init(23'h000000),
    .width(23)
) reg_PR23_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR23_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR23_inst0__CE_out;
endmodule

module Register_unq3 (
    input [16:0] I,
    output [16:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [16:0] reg_PR17_inst0__CE_out;
regCE_arst #(
    .init(17'h00000),
    .width(17)
) reg_PR17_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR17_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR17_inst0__CE_out;
endmodule

module Register_unq2 (
    input [23:0] I,
    output [23:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [23:0] reg_PR24_inst0__CE_out;
regCE_arst #(
    .init(24'h000000),
    .width(24)
) reg_PR24_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR24_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR24_inst0__CE_out;
endmodule

module Register_unq12 (
    input [30:0] I,
    output [30:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [30:0] reg_PR31_inst0__CE_out;
regCE_arst #(
    .init(31'h00000000),
    .width(31)
) reg_PR31_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR31_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR31_inst0__CE_out;
endmodule

module Register_unq11 (
    input [26:0] I,
    output [26:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [26:0] reg_PR27_inst0__CE_out;
regCE_arst #(
    .init(27'h0000000),
    .width(27)
) reg_PR27_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR27_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR27_inst0__CE_out;
endmodule

module Register_unq10 (
    input [25:0] I,
    output [25:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [25:0] reg_PR26_inst0__CE_out;
regCE_arst #(
    .init(26'h0000000),
    .width(26)
) reg_PR26_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR26_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR26_inst0__CE_out;
endmodule

module Register_unq1 (
    input [4:0] I,
    output [4:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [4:0] reg_PR5_inst0__CE_out;
regCE_arst #(
    .init(5'h00),
    .width(5)
) reg_PR5_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR5_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR5_inst0__CE_out;
endmodule

module Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 (
    input [15:0] I,
    output [15:0] O,
    input CLK,
    input CE
);
wire [15:0] value__CE_out;
regCE #(
    .width(16)
) value__CE (
    .in(I),
    .ce(CE),
    .out(value__CE_out),
    .clk(CLK)
);
assign O = value__CE_out;
endmodule

module Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 (
    input [0:0] I,
    output [0:0] O,
    input CLK,
    input CE
);
wire [0:0] value__CE_out;
regCE #(
    .width(1)
) value__CE (
    .in(I),
    .ce(CE),
    .out(value__CE_out),
    .clk(CLK)
);
assign O = value__CE_out;
endmodule

module Register (
    input [31:0] I,
    output [31:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [31:0] reg_PR32_inst0__CE_out;
regCE_arst #(
    .init(32'h00000000),
    .width(32)
) reg_PR32_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR32_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR32_inst0__CE_out;
endmodule

module RMUX_T4_WEST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[19:19];
endmodule

module RMUX_T4_WEST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[19:19];
endmodule

module RMUX_T4_SOUTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[18:18];
endmodule

module RMUX_T4_SOUTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[18:18];
endmodule

module RMUX_T4_NORTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[17:17];
endmodule

module RMUX_T4_NORTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[17:17];
endmodule

module RMUX_T4_EAST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[16:16];
endmodule

module RMUX_T4_EAST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[16:16];
endmodule

module RMUX_T3_WEST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[15:15];
endmodule

module RMUX_T3_WEST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[15:15];
endmodule

module RMUX_T3_SOUTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[14:14];
endmodule

module RMUX_T3_SOUTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[14:14];
endmodule

module RMUX_T3_NORTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[13:13];
endmodule

module RMUX_T3_NORTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[13:13];
endmodule

module RMUX_T3_EAST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[12:12];
endmodule

module RMUX_T3_EAST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[12:12];
endmodule

module RMUX_T2_WEST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[11:11];
endmodule

module RMUX_T2_WEST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[11:11];
endmodule

module RMUX_T2_SOUTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[10:10];
endmodule

module RMUX_T2_SOUTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[10:10];
endmodule

module RMUX_T2_NORTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[9:9];
endmodule

module RMUX_T2_NORTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[9:9];
endmodule

module RMUX_T2_EAST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[8:8];
endmodule

module RMUX_T2_EAST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[8:8];
endmodule

module RMUX_T1_WEST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[7:7];
endmodule

module RMUX_T1_WEST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[7:7];
endmodule

module RMUX_T1_SOUTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[6:6];
endmodule

module RMUX_T1_SOUTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[6:6];
endmodule

module RMUX_T1_NORTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[5:5];
endmodule

module RMUX_T1_NORTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[5:5];
endmodule

module RMUX_T1_EAST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[4:4];
endmodule

module RMUX_T1_EAST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[4:4];
endmodule

module RMUX_T0_WEST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[3:3];
endmodule

module RMUX_T0_WEST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[3:3];
endmodule

module RMUX_T0_SOUTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[2:2];
endmodule

module RMUX_T0_SOUTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[2:2];
endmodule

module RMUX_T0_NORTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[1:1];
endmodule

module RMUX_T0_NORTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[1:1];
endmodule

module RMUX_T0_EAST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[0:0];
endmodule

module RMUX_T0_EAST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[0:0];
endmodule

module PowerDomainOR (
    input [31:0] I0,
    input [31:0] I1,
    output [31:0] O,
    input [0:0] I_not
);
wire [0:0] Invert1_inst0_out;
wire [0:0] and1_inst0_out;
wire [0:0] and1_inst1_out;
wire [0:0] and1_inst10_out;
wire [0:0] and1_inst11_out;
wire [0:0] and1_inst12_out;
wire [0:0] and1_inst13_out;
wire [0:0] and1_inst14_out;
wire [0:0] and1_inst15_out;
wire [0:0] and1_inst16_out;
wire [0:0] and1_inst17_out;
wire [0:0] and1_inst18_out;
wire [0:0] and1_inst19_out;
wire [0:0] and1_inst2_out;
wire [0:0] and1_inst20_out;
wire [0:0] and1_inst21_out;
wire [0:0] and1_inst22_out;
wire [0:0] and1_inst23_out;
wire [0:0] and1_inst24_out;
wire [0:0] and1_inst25_out;
wire [0:0] and1_inst26_out;
wire [0:0] and1_inst27_out;
wire [0:0] and1_inst28_out;
wire [0:0] and1_inst29_out;
wire [0:0] and1_inst3_out;
wire [0:0] and1_inst30_out;
wire [0:0] and1_inst31_out;
wire [0:0] and1_inst4_out;
wire [0:0] and1_inst5_out;
wire [0:0] and1_inst6_out;
wire [0:0] and1_inst7_out;
wire [0:0] and1_inst8_out;
wire [0:0] and1_inst9_out;
wire [31:0] or32_inst0_out;
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(I_not),
    .out(Invert1_inst0_out)
);
coreir_and #(
    .width(1)
) and1_inst0 (
    .in0(I0[0]),
    .in1(Invert1_inst0_out),
    .out(and1_inst0_out)
);
coreir_and #(
    .width(1)
) and1_inst1 (
    .in0(I0[1]),
    .in1(Invert1_inst0_out),
    .out(and1_inst1_out)
);
coreir_and #(
    .width(1)
) and1_inst10 (
    .in0(I0[10]),
    .in1(Invert1_inst0_out),
    .out(and1_inst10_out)
);
coreir_and #(
    .width(1)
) and1_inst11 (
    .in0(I0[11]),
    .in1(Invert1_inst0_out),
    .out(and1_inst11_out)
);
coreir_and #(
    .width(1)
) and1_inst12 (
    .in0(I0[12]),
    .in1(Invert1_inst0_out),
    .out(and1_inst12_out)
);
coreir_and #(
    .width(1)
) and1_inst13 (
    .in0(I0[13]),
    .in1(Invert1_inst0_out),
    .out(and1_inst13_out)
);
coreir_and #(
    .width(1)
) and1_inst14 (
    .in0(I0[14]),
    .in1(Invert1_inst0_out),
    .out(and1_inst14_out)
);
coreir_and #(
    .width(1)
) and1_inst15 (
    .in0(I0[15]),
    .in1(Invert1_inst0_out),
    .out(and1_inst15_out)
);
coreir_and #(
    .width(1)
) and1_inst16 (
    .in0(I0[16]),
    .in1(Invert1_inst0_out),
    .out(and1_inst16_out)
);
coreir_and #(
    .width(1)
) and1_inst17 (
    .in0(I0[17]),
    .in1(Invert1_inst0_out),
    .out(and1_inst17_out)
);
coreir_and #(
    .width(1)
) and1_inst18 (
    .in0(I0[18]),
    .in1(Invert1_inst0_out),
    .out(and1_inst18_out)
);
coreir_and #(
    .width(1)
) and1_inst19 (
    .in0(I0[19]),
    .in1(Invert1_inst0_out),
    .out(and1_inst19_out)
);
coreir_and #(
    .width(1)
) and1_inst2 (
    .in0(I0[2]),
    .in1(Invert1_inst0_out),
    .out(and1_inst2_out)
);
coreir_and #(
    .width(1)
) and1_inst20 (
    .in0(I0[20]),
    .in1(Invert1_inst0_out),
    .out(and1_inst20_out)
);
coreir_and #(
    .width(1)
) and1_inst21 (
    .in0(I0[21]),
    .in1(Invert1_inst0_out),
    .out(and1_inst21_out)
);
coreir_and #(
    .width(1)
) and1_inst22 (
    .in0(I0[22]),
    .in1(Invert1_inst0_out),
    .out(and1_inst22_out)
);
coreir_and #(
    .width(1)
) and1_inst23 (
    .in0(I0[23]),
    .in1(Invert1_inst0_out),
    .out(and1_inst23_out)
);
coreir_and #(
    .width(1)
) and1_inst24 (
    .in0(I0[24]),
    .in1(Invert1_inst0_out),
    .out(and1_inst24_out)
);
coreir_and #(
    .width(1)
) and1_inst25 (
    .in0(I0[25]),
    .in1(Invert1_inst0_out),
    .out(and1_inst25_out)
);
coreir_and #(
    .width(1)
) and1_inst26 (
    .in0(I0[26]),
    .in1(Invert1_inst0_out),
    .out(and1_inst26_out)
);
coreir_and #(
    .width(1)
) and1_inst27 (
    .in0(I0[27]),
    .in1(Invert1_inst0_out),
    .out(and1_inst27_out)
);
coreir_and #(
    .width(1)
) and1_inst28 (
    .in0(I0[28]),
    .in1(Invert1_inst0_out),
    .out(and1_inst28_out)
);
coreir_and #(
    .width(1)
) and1_inst29 (
    .in0(I0[29]),
    .in1(Invert1_inst0_out),
    .out(and1_inst29_out)
);
coreir_and #(
    .width(1)
) and1_inst3 (
    .in0(I0[3]),
    .in1(Invert1_inst0_out),
    .out(and1_inst3_out)
);
coreir_and #(
    .width(1)
) and1_inst30 (
    .in0(I0[30]),
    .in1(Invert1_inst0_out),
    .out(and1_inst30_out)
);
coreir_and #(
    .width(1)
) and1_inst31 (
    .in0(I0[31]),
    .in1(Invert1_inst0_out),
    .out(and1_inst31_out)
);
coreir_and #(
    .width(1)
) and1_inst4 (
    .in0(I0[4]),
    .in1(Invert1_inst0_out),
    .out(and1_inst4_out)
);
coreir_and #(
    .width(1)
) and1_inst5 (
    .in0(I0[5]),
    .in1(Invert1_inst0_out),
    .out(and1_inst5_out)
);
coreir_and #(
    .width(1)
) and1_inst6 (
    .in0(I0[6]),
    .in1(Invert1_inst0_out),
    .out(and1_inst6_out)
);
coreir_and #(
    .width(1)
) and1_inst7 (
    .in0(I0[7]),
    .in1(Invert1_inst0_out),
    .out(and1_inst7_out)
);
coreir_and #(
    .width(1)
) and1_inst8 (
    .in0(I0[8]),
    .in1(Invert1_inst0_out),
    .out(and1_inst8_out)
);
coreir_and #(
    .width(1)
) and1_inst9 (
    .in0(I0[9]),
    .in1(Invert1_inst0_out),
    .out(and1_inst9_out)
);
wire [31:0] or32_inst0_in0;
assign or32_inst0_in0 = {and1_inst31_out[0],and1_inst30_out[0],and1_inst29_out[0],and1_inst28_out[0],and1_inst27_out[0],and1_inst26_out[0],and1_inst25_out[0],and1_inst24_out[0],and1_inst23_out[0],and1_inst22_out[0],and1_inst21_out[0],and1_inst20_out[0],and1_inst19_out[0],and1_inst18_out[0],and1_inst17_out[0],and1_inst16_out[0],and1_inst15_out[0],and1_inst14_out[0],and1_inst13_out[0],and1_inst12_out[0],and1_inst11_out[0],and1_inst10_out[0],and1_inst9_out[0],and1_inst8_out[0],and1_inst7_out[0],and1_inst6_out[0],and1_inst5_out[0],and1_inst4_out[0],and1_inst3_out[0],and1_inst2_out[0],and1_inst1_out[0],and1_inst0_out[0]};
coreir_or #(
    .width(32)
) or32_inst0 (
    .in0(or32_inst0_in0),
    .in1(I1),
    .out(or32_inst0_out)
);
assign O = or32_inst0_out;
endmodule

module Or4x32 (
    input [31:0] I0,
    input [31:0] I1,
    input [31:0] I2,
    input [31:0] I3,
    output [31:0] O
);
wire orr_inst0_out;
wire orr_inst1_out;
wire orr_inst10_out;
wire orr_inst11_out;
wire orr_inst12_out;
wire orr_inst13_out;
wire orr_inst14_out;
wire orr_inst15_out;
wire orr_inst16_out;
wire orr_inst17_out;
wire orr_inst18_out;
wire orr_inst19_out;
wire orr_inst2_out;
wire orr_inst20_out;
wire orr_inst21_out;
wire orr_inst22_out;
wire orr_inst23_out;
wire orr_inst24_out;
wire orr_inst25_out;
wire orr_inst26_out;
wire orr_inst27_out;
wire orr_inst28_out;
wire orr_inst29_out;
wire orr_inst3_out;
wire orr_inst30_out;
wire orr_inst31_out;
wire orr_inst4_out;
wire orr_inst5_out;
wire orr_inst6_out;
wire orr_inst7_out;
wire orr_inst8_out;
wire orr_inst9_out;
wire [3:0] orr_inst0_in;
assign orr_inst0_in = {I3[0],I2[0],I1[0],I0[0]};
coreir_orr #(
    .width(4)
) orr_inst0 (
    .in(orr_inst0_in),
    .out(orr_inst0_out)
);
wire [3:0] orr_inst1_in;
assign orr_inst1_in = {I3[1],I2[1],I1[1],I0[1]};
coreir_orr #(
    .width(4)
) orr_inst1 (
    .in(orr_inst1_in),
    .out(orr_inst1_out)
);
wire [3:0] orr_inst10_in;
assign orr_inst10_in = {I3[10],I2[10],I1[10],I0[10]};
coreir_orr #(
    .width(4)
) orr_inst10 (
    .in(orr_inst10_in),
    .out(orr_inst10_out)
);
wire [3:0] orr_inst11_in;
assign orr_inst11_in = {I3[11],I2[11],I1[11],I0[11]};
coreir_orr #(
    .width(4)
) orr_inst11 (
    .in(orr_inst11_in),
    .out(orr_inst11_out)
);
wire [3:0] orr_inst12_in;
assign orr_inst12_in = {I3[12],I2[12],I1[12],I0[12]};
coreir_orr #(
    .width(4)
) orr_inst12 (
    .in(orr_inst12_in),
    .out(orr_inst12_out)
);
wire [3:0] orr_inst13_in;
assign orr_inst13_in = {I3[13],I2[13],I1[13],I0[13]};
coreir_orr #(
    .width(4)
) orr_inst13 (
    .in(orr_inst13_in),
    .out(orr_inst13_out)
);
wire [3:0] orr_inst14_in;
assign orr_inst14_in = {I3[14],I2[14],I1[14],I0[14]};
coreir_orr #(
    .width(4)
) orr_inst14 (
    .in(orr_inst14_in),
    .out(orr_inst14_out)
);
wire [3:0] orr_inst15_in;
assign orr_inst15_in = {I3[15],I2[15],I1[15],I0[15]};
coreir_orr #(
    .width(4)
) orr_inst15 (
    .in(orr_inst15_in),
    .out(orr_inst15_out)
);
wire [3:0] orr_inst16_in;
assign orr_inst16_in = {I3[16],I2[16],I1[16],I0[16]};
coreir_orr #(
    .width(4)
) orr_inst16 (
    .in(orr_inst16_in),
    .out(orr_inst16_out)
);
wire [3:0] orr_inst17_in;
assign orr_inst17_in = {I3[17],I2[17],I1[17],I0[17]};
coreir_orr #(
    .width(4)
) orr_inst17 (
    .in(orr_inst17_in),
    .out(orr_inst17_out)
);
wire [3:0] orr_inst18_in;
assign orr_inst18_in = {I3[18],I2[18],I1[18],I0[18]};
coreir_orr #(
    .width(4)
) orr_inst18 (
    .in(orr_inst18_in),
    .out(orr_inst18_out)
);
wire [3:0] orr_inst19_in;
assign orr_inst19_in = {I3[19],I2[19],I1[19],I0[19]};
coreir_orr #(
    .width(4)
) orr_inst19 (
    .in(orr_inst19_in),
    .out(orr_inst19_out)
);
wire [3:0] orr_inst2_in;
assign orr_inst2_in = {I3[2],I2[2],I1[2],I0[2]};
coreir_orr #(
    .width(4)
) orr_inst2 (
    .in(orr_inst2_in),
    .out(orr_inst2_out)
);
wire [3:0] orr_inst20_in;
assign orr_inst20_in = {I3[20],I2[20],I1[20],I0[20]};
coreir_orr #(
    .width(4)
) orr_inst20 (
    .in(orr_inst20_in),
    .out(orr_inst20_out)
);
wire [3:0] orr_inst21_in;
assign orr_inst21_in = {I3[21],I2[21],I1[21],I0[21]};
coreir_orr #(
    .width(4)
) orr_inst21 (
    .in(orr_inst21_in),
    .out(orr_inst21_out)
);
wire [3:0] orr_inst22_in;
assign orr_inst22_in = {I3[22],I2[22],I1[22],I0[22]};
coreir_orr #(
    .width(4)
) orr_inst22 (
    .in(orr_inst22_in),
    .out(orr_inst22_out)
);
wire [3:0] orr_inst23_in;
assign orr_inst23_in = {I3[23],I2[23],I1[23],I0[23]};
coreir_orr #(
    .width(4)
) orr_inst23 (
    .in(orr_inst23_in),
    .out(orr_inst23_out)
);
wire [3:0] orr_inst24_in;
assign orr_inst24_in = {I3[24],I2[24],I1[24],I0[24]};
coreir_orr #(
    .width(4)
) orr_inst24 (
    .in(orr_inst24_in),
    .out(orr_inst24_out)
);
wire [3:0] orr_inst25_in;
assign orr_inst25_in = {I3[25],I2[25],I1[25],I0[25]};
coreir_orr #(
    .width(4)
) orr_inst25 (
    .in(orr_inst25_in),
    .out(orr_inst25_out)
);
wire [3:0] orr_inst26_in;
assign orr_inst26_in = {I3[26],I2[26],I1[26],I0[26]};
coreir_orr #(
    .width(4)
) orr_inst26 (
    .in(orr_inst26_in),
    .out(orr_inst26_out)
);
wire [3:0] orr_inst27_in;
assign orr_inst27_in = {I3[27],I2[27],I1[27],I0[27]};
coreir_orr #(
    .width(4)
) orr_inst27 (
    .in(orr_inst27_in),
    .out(orr_inst27_out)
);
wire [3:0] orr_inst28_in;
assign orr_inst28_in = {I3[28],I2[28],I1[28],I0[28]};
coreir_orr #(
    .width(4)
) orr_inst28 (
    .in(orr_inst28_in),
    .out(orr_inst28_out)
);
wire [3:0] orr_inst29_in;
assign orr_inst29_in = {I3[29],I2[29],I1[29],I0[29]};
coreir_orr #(
    .width(4)
) orr_inst29 (
    .in(orr_inst29_in),
    .out(orr_inst29_out)
);
wire [3:0] orr_inst3_in;
assign orr_inst3_in = {I3[3],I2[3],I1[3],I0[3]};
coreir_orr #(
    .width(4)
) orr_inst3 (
    .in(orr_inst3_in),
    .out(orr_inst3_out)
);
wire [3:0] orr_inst30_in;
assign orr_inst30_in = {I3[30],I2[30],I1[30],I0[30]};
coreir_orr #(
    .width(4)
) orr_inst30 (
    .in(orr_inst30_in),
    .out(orr_inst30_out)
);
wire [3:0] orr_inst31_in;
assign orr_inst31_in = {I3[31],I2[31],I1[31],I0[31]};
coreir_orr #(
    .width(4)
) orr_inst31 (
    .in(orr_inst31_in),
    .out(orr_inst31_out)
);
wire [3:0] orr_inst4_in;
assign orr_inst4_in = {I3[4],I2[4],I1[4],I0[4]};
coreir_orr #(
    .width(4)
) orr_inst4 (
    .in(orr_inst4_in),
    .out(orr_inst4_out)
);
wire [3:0] orr_inst5_in;
assign orr_inst5_in = {I3[5],I2[5],I1[5],I0[5]};
coreir_orr #(
    .width(4)
) orr_inst5 (
    .in(orr_inst5_in),
    .out(orr_inst5_out)
);
wire [3:0] orr_inst6_in;
assign orr_inst6_in = {I3[6],I2[6],I1[6],I0[6]};
coreir_orr #(
    .width(4)
) orr_inst6 (
    .in(orr_inst6_in),
    .out(orr_inst6_out)
);
wire [3:0] orr_inst7_in;
assign orr_inst7_in = {I3[7],I2[7],I1[7],I0[7]};
coreir_orr #(
    .width(4)
) orr_inst7 (
    .in(orr_inst7_in),
    .out(orr_inst7_out)
);
wire [3:0] orr_inst8_in;
assign orr_inst8_in = {I3[8],I2[8],I1[8],I0[8]};
coreir_orr #(
    .width(4)
) orr_inst8 (
    .in(orr_inst8_in),
    .out(orr_inst8_out)
);
wire [3:0] orr_inst9_in;
assign orr_inst9_in = {I3[9],I2[9],I1[9],I0[9]};
coreir_orr #(
    .width(4)
) orr_inst9 (
    .in(orr_inst9_in),
    .out(orr_inst9_out)
);
assign O = {orr_inst31_out,orr_inst30_out,orr_inst29_out,orr_inst28_out,orr_inst27_out,orr_inst26_out,orr_inst25_out,orr_inst24_out,orr_inst23_out,orr_inst22_out,orr_inst21_out,orr_inst20_out,orr_inst19_out,orr_inst18_out,orr_inst17_out,orr_inst16_out,orr_inst15_out,orr_inst14_out,orr_inst13_out,orr_inst12_out,orr_inst11_out,orr_inst10_out,orr_inst9_out,orr_inst8_out,orr_inst7_out,orr_inst6_out,orr_inst5_out,orr_inst4_out,orr_inst3_out,orr_inst2_out,orr_inst1_out,orr_inst0_out};
endmodule

module Or3x8 (
    input [7:0] I0,
    input [7:0] I1,
    input [7:0] I2,
    output [7:0] O
);
wire orr_inst0_out;
wire orr_inst1_out;
wire orr_inst2_out;
wire orr_inst3_out;
wire orr_inst4_out;
wire orr_inst5_out;
wire orr_inst6_out;
wire orr_inst7_out;
wire [2:0] orr_inst0_in;
assign orr_inst0_in = {I2[0],I1[0],I0[0]};
coreir_orr #(
    .width(3)
) orr_inst0 (
    .in(orr_inst0_in),
    .out(orr_inst0_out)
);
wire [2:0] orr_inst1_in;
assign orr_inst1_in = {I2[1],I1[1],I0[1]};
coreir_orr #(
    .width(3)
) orr_inst1 (
    .in(orr_inst1_in),
    .out(orr_inst1_out)
);
wire [2:0] orr_inst2_in;
assign orr_inst2_in = {I2[2],I1[2],I0[2]};
coreir_orr #(
    .width(3)
) orr_inst2 (
    .in(orr_inst2_in),
    .out(orr_inst2_out)
);
wire [2:0] orr_inst3_in;
assign orr_inst3_in = {I2[3],I1[3],I0[3]};
coreir_orr #(
    .width(3)
) orr_inst3 (
    .in(orr_inst3_in),
    .out(orr_inst3_out)
);
wire [2:0] orr_inst4_in;
assign orr_inst4_in = {I2[4],I1[4],I0[4]};
coreir_orr #(
    .width(3)
) orr_inst4 (
    .in(orr_inst4_in),
    .out(orr_inst4_out)
);
wire [2:0] orr_inst5_in;
assign orr_inst5_in = {I2[5],I1[5],I0[5]};
coreir_orr #(
    .width(3)
) orr_inst5 (
    .in(orr_inst5_in),
    .out(orr_inst5_out)
);
wire [2:0] orr_inst6_in;
assign orr_inst6_in = {I2[6],I1[6],I0[6]};
coreir_orr #(
    .width(3)
) orr_inst6 (
    .in(orr_inst6_in),
    .out(orr_inst6_out)
);
wire [2:0] orr_inst7_in;
assign orr_inst7_in = {I2[7],I1[7],I0[7]};
coreir_orr #(
    .width(3)
) orr_inst7 (
    .in(orr_inst7_in),
    .out(orr_inst7_out)
);
assign O = {orr_inst7_out,orr_inst6_out,orr_inst5_out,orr_inst4_out,orr_inst3_out,orr_inst2_out,orr_inst1_out,orr_inst0_out};
endmodule

module Or3x32 (
    input [31:0] I0,
    input [31:0] I1,
    input [31:0] I2,
    output [31:0] O
);
wire orr_inst0_out;
wire orr_inst1_out;
wire orr_inst10_out;
wire orr_inst11_out;
wire orr_inst12_out;
wire orr_inst13_out;
wire orr_inst14_out;
wire orr_inst15_out;
wire orr_inst16_out;
wire orr_inst17_out;
wire orr_inst18_out;
wire orr_inst19_out;
wire orr_inst2_out;
wire orr_inst20_out;
wire orr_inst21_out;
wire orr_inst22_out;
wire orr_inst23_out;
wire orr_inst24_out;
wire orr_inst25_out;
wire orr_inst26_out;
wire orr_inst27_out;
wire orr_inst28_out;
wire orr_inst29_out;
wire orr_inst3_out;
wire orr_inst30_out;
wire orr_inst31_out;
wire orr_inst4_out;
wire orr_inst5_out;
wire orr_inst6_out;
wire orr_inst7_out;
wire orr_inst8_out;
wire orr_inst9_out;
wire [2:0] orr_inst0_in;
assign orr_inst0_in = {I2[0],I1[0],I0[0]};
coreir_orr #(
    .width(3)
) orr_inst0 (
    .in(orr_inst0_in),
    .out(orr_inst0_out)
);
wire [2:0] orr_inst1_in;
assign orr_inst1_in = {I2[1],I1[1],I0[1]};
coreir_orr #(
    .width(3)
) orr_inst1 (
    .in(orr_inst1_in),
    .out(orr_inst1_out)
);
wire [2:0] orr_inst10_in;
assign orr_inst10_in = {I2[10],I1[10],I0[10]};
coreir_orr #(
    .width(3)
) orr_inst10 (
    .in(orr_inst10_in),
    .out(orr_inst10_out)
);
wire [2:0] orr_inst11_in;
assign orr_inst11_in = {I2[11],I1[11],I0[11]};
coreir_orr #(
    .width(3)
) orr_inst11 (
    .in(orr_inst11_in),
    .out(orr_inst11_out)
);
wire [2:0] orr_inst12_in;
assign orr_inst12_in = {I2[12],I1[12],I0[12]};
coreir_orr #(
    .width(3)
) orr_inst12 (
    .in(orr_inst12_in),
    .out(orr_inst12_out)
);
wire [2:0] orr_inst13_in;
assign orr_inst13_in = {I2[13],I1[13],I0[13]};
coreir_orr #(
    .width(3)
) orr_inst13 (
    .in(orr_inst13_in),
    .out(orr_inst13_out)
);
wire [2:0] orr_inst14_in;
assign orr_inst14_in = {I2[14],I1[14],I0[14]};
coreir_orr #(
    .width(3)
) orr_inst14 (
    .in(orr_inst14_in),
    .out(orr_inst14_out)
);
wire [2:0] orr_inst15_in;
assign orr_inst15_in = {I2[15],I1[15],I0[15]};
coreir_orr #(
    .width(3)
) orr_inst15 (
    .in(orr_inst15_in),
    .out(orr_inst15_out)
);
wire [2:0] orr_inst16_in;
assign orr_inst16_in = {I2[16],I1[16],I0[16]};
coreir_orr #(
    .width(3)
) orr_inst16 (
    .in(orr_inst16_in),
    .out(orr_inst16_out)
);
wire [2:0] orr_inst17_in;
assign orr_inst17_in = {I2[17],I1[17],I0[17]};
coreir_orr #(
    .width(3)
) orr_inst17 (
    .in(orr_inst17_in),
    .out(orr_inst17_out)
);
wire [2:0] orr_inst18_in;
assign orr_inst18_in = {I2[18],I1[18],I0[18]};
coreir_orr #(
    .width(3)
) orr_inst18 (
    .in(orr_inst18_in),
    .out(orr_inst18_out)
);
wire [2:0] orr_inst19_in;
assign orr_inst19_in = {I2[19],I1[19],I0[19]};
coreir_orr #(
    .width(3)
) orr_inst19 (
    .in(orr_inst19_in),
    .out(orr_inst19_out)
);
wire [2:0] orr_inst2_in;
assign orr_inst2_in = {I2[2],I1[2],I0[2]};
coreir_orr #(
    .width(3)
) orr_inst2 (
    .in(orr_inst2_in),
    .out(orr_inst2_out)
);
wire [2:0] orr_inst20_in;
assign orr_inst20_in = {I2[20],I1[20],I0[20]};
coreir_orr #(
    .width(3)
) orr_inst20 (
    .in(orr_inst20_in),
    .out(orr_inst20_out)
);
wire [2:0] orr_inst21_in;
assign orr_inst21_in = {I2[21],I1[21],I0[21]};
coreir_orr #(
    .width(3)
) orr_inst21 (
    .in(orr_inst21_in),
    .out(orr_inst21_out)
);
wire [2:0] orr_inst22_in;
assign orr_inst22_in = {I2[22],I1[22],I0[22]};
coreir_orr #(
    .width(3)
) orr_inst22 (
    .in(orr_inst22_in),
    .out(orr_inst22_out)
);
wire [2:0] orr_inst23_in;
assign orr_inst23_in = {I2[23],I1[23],I0[23]};
coreir_orr #(
    .width(3)
) orr_inst23 (
    .in(orr_inst23_in),
    .out(orr_inst23_out)
);
wire [2:0] orr_inst24_in;
assign orr_inst24_in = {I2[24],I1[24],I0[24]};
coreir_orr #(
    .width(3)
) orr_inst24 (
    .in(orr_inst24_in),
    .out(orr_inst24_out)
);
wire [2:0] orr_inst25_in;
assign orr_inst25_in = {I2[25],I1[25],I0[25]};
coreir_orr #(
    .width(3)
) orr_inst25 (
    .in(orr_inst25_in),
    .out(orr_inst25_out)
);
wire [2:0] orr_inst26_in;
assign orr_inst26_in = {I2[26],I1[26],I0[26]};
coreir_orr #(
    .width(3)
) orr_inst26 (
    .in(orr_inst26_in),
    .out(orr_inst26_out)
);
wire [2:0] orr_inst27_in;
assign orr_inst27_in = {I2[27],I1[27],I0[27]};
coreir_orr #(
    .width(3)
) orr_inst27 (
    .in(orr_inst27_in),
    .out(orr_inst27_out)
);
wire [2:0] orr_inst28_in;
assign orr_inst28_in = {I2[28],I1[28],I0[28]};
coreir_orr #(
    .width(3)
) orr_inst28 (
    .in(orr_inst28_in),
    .out(orr_inst28_out)
);
wire [2:0] orr_inst29_in;
assign orr_inst29_in = {I2[29],I1[29],I0[29]};
coreir_orr #(
    .width(3)
) orr_inst29 (
    .in(orr_inst29_in),
    .out(orr_inst29_out)
);
wire [2:0] orr_inst3_in;
assign orr_inst3_in = {I2[3],I1[3],I0[3]};
coreir_orr #(
    .width(3)
) orr_inst3 (
    .in(orr_inst3_in),
    .out(orr_inst3_out)
);
wire [2:0] orr_inst30_in;
assign orr_inst30_in = {I2[30],I1[30],I0[30]};
coreir_orr #(
    .width(3)
) orr_inst30 (
    .in(orr_inst30_in),
    .out(orr_inst30_out)
);
wire [2:0] orr_inst31_in;
assign orr_inst31_in = {I2[31],I1[31],I0[31]};
coreir_orr #(
    .width(3)
) orr_inst31 (
    .in(orr_inst31_in),
    .out(orr_inst31_out)
);
wire [2:0] orr_inst4_in;
assign orr_inst4_in = {I2[4],I1[4],I0[4]};
coreir_orr #(
    .width(3)
) orr_inst4 (
    .in(orr_inst4_in),
    .out(orr_inst4_out)
);
wire [2:0] orr_inst5_in;
assign orr_inst5_in = {I2[5],I1[5],I0[5]};
coreir_orr #(
    .width(3)
) orr_inst5 (
    .in(orr_inst5_in),
    .out(orr_inst5_out)
);
wire [2:0] orr_inst6_in;
assign orr_inst6_in = {I2[6],I1[6],I0[6]};
coreir_orr #(
    .width(3)
) orr_inst6 (
    .in(orr_inst6_in),
    .out(orr_inst6_out)
);
wire [2:0] orr_inst7_in;
assign orr_inst7_in = {I2[7],I1[7],I0[7]};
coreir_orr #(
    .width(3)
) orr_inst7 (
    .in(orr_inst7_in),
    .out(orr_inst7_out)
);
wire [2:0] orr_inst8_in;
assign orr_inst8_in = {I2[8],I1[8],I0[8]};
coreir_orr #(
    .width(3)
) orr_inst8 (
    .in(orr_inst8_in),
    .out(orr_inst8_out)
);
wire [2:0] orr_inst9_in;
assign orr_inst9_in = {I2[9],I1[9],I0[9]};
coreir_orr #(
    .width(3)
) orr_inst9 (
    .in(orr_inst9_in),
    .out(orr_inst9_out)
);
assign O = {orr_inst31_out,orr_inst30_out,orr_inst29_out,orr_inst28_out,orr_inst27_out,orr_inst26_out,orr_inst25_out,orr_inst24_out,orr_inst23_out,orr_inst22_out,orr_inst21_out,orr_inst20_out,orr_inst19_out,orr_inst18_out,orr_inst17_out,orr_inst16_out,orr_inst15_out,orr_inst14_out,orr_inst13_out,orr_inst12_out,orr_inst11_out,orr_inst10_out,orr_inst9_out,orr_inst8_out,orr_inst7_out,orr_inst6_out,orr_inst5_out,orr_inst4_out,orr_inst3_out,orr_inst2_out,orr_inst1_out,orr_inst0_out};
endmodule

module MuxWrapper_1_16 (
    input [15:0] I,
    output [15:0] O
);
assign O = I;
endmodule

module MuxWrapper_1_1 (
    input [0:0] I,
    output [0:0] O
);
assign O = I;
endmodule

module MuxWrapperAOI_1_1_Regular (
    input [0:0] I,
    output [0:0] O
);
assign O = I;
endmodule

module MuxWrapperAOI_1_1_Const (
    input [0:0] I,
    output [0:0] O
);
assign O = I;
endmodule

module MuxWrapperAOI_1_16_Regular (
    input [15:0] I,
    output [15:0] O
);
assign O = I;
endmodule

module MuxWrapperAOI_1_16_Const (
    input [15:0] I,
    output [15:0] O
);
assign O = I;
endmodule

module Tile_io_core (
    input [15:0] tile_id,
    input [0:0] glb2io_1,
    input [0:0] f2io_1,
    output [0:0] io2glb_1,
    output [0:0] io2f_1,
    input [15:0] glb2io_16,
    input [15:0] f2io_16,
    output [15:0] io2glb_16,
    output [15:0] io2f_16,
    output [8:0] hi,
    output [7:0] lo
);
wire [0:0] CB_f2io_1$CB_f2io_1_O;
wire [15:0] CB_f2io_16$CB_f2io_16_O;
wire [7:0] const_0_8_out;
wire [8:0] const_511_9_out;
wire [15:0] io_core_inst0_io2glb_16;
wire [0:0] io_core_inst0_io2glb_1;
wire [15:0] io_core_inst0_io2f_16;
wire [0:0] io_core_inst0_io2f_1;
MuxWrapperAOI_1_1_Const CB_f2io_1$CB_f2io_1 (
    .I(f2io_1),
    .O(CB_f2io_1$CB_f2io_1_O)
);
MuxWrapperAOI_1_16_Const CB_f2io_16$CB_f2io_16 (
    .I(f2io_16),
    .O(CB_f2io_16$CB_f2io_16_O)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
coreir_const #(
    .value(9'h1ff),
    .width(9)
) const_511_9 (
    .out(const_511_9_out)
);
io_core io_core_inst0 (
    .glb2io_16(glb2io_16),
    .glb2io_1(glb2io_1),
    .io2glb_16(io_core_inst0_io2glb_16),
    .io2glb_1(io_core_inst0_io2glb_1),
    .f2io_16(CB_f2io_16$CB_f2io_16_O),
    .f2io_1(CB_f2io_1$CB_f2io_1_O),
    .io2f_16(io_core_inst0_io2f_16),
    .io2f_1(io_core_inst0_io2f_1)
);
assign io2glb_1 = io_core_inst0_io2glb_1;
assign io2f_1 = io_core_inst0_io2f_1;
assign io2glb_16 = io_core_inst0_io2glb_16;
assign io2f_16 = io_core_inst0_io2f_16;
assign hi = const_511_9_out;
assign lo = const_0_8_out;
endmodule

module MuxWrapperAOIImpl_7_1 (
    input [0:0] I_0,
    input [0:0] I_1,
    input [0:0] I_2,
    input [0:0] I_3,
    input [0:0] I_4,
    input [0:0] I_5,
    input [0:0] I_6,
    output [0:0] O,
    input [2:0] S
);
wire [0:0] mux_aoi_7_1_inst0_O;
mux_aoi_7_1 mux_aoi_7_1_inst0 (
    .I0(I_0),
    .I1(I_1),
    .I2(I_2),
    .I3(I_3),
    .I4(I_4),
    .I5(I_5),
    .I6(I_6),
    .S(S),
    .O(mux_aoi_7_1_inst0_O)
);
assign O = mux_aoi_7_1_inst0_O;
endmodule

module MuxWrapperAOIImpl_5_16 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    output [15:0] O,
    input [2:0] S
);
wire [15:0] mux_aoi_5_16_inst0_O;
mux_aoi_5_16 mux_aoi_5_16_inst0 (
    .I0(I_0),
    .I1(I_1),
    .I2(I_2),
    .I3(I_3),
    .I4(I_4),
    .S(S),
    .O(mux_aoi_5_16_inst0_O)
);
assign O = mux_aoi_5_16_inst0_O;
endmodule

module MuxWrapperAOIImpl_5_1 (
    input [0:0] I_0,
    input [0:0] I_1,
    input [0:0] I_2,
    input [0:0] I_3,
    input [0:0] I_4,
    output [0:0] O,
    input [2:0] S
);
wire [0:0] mux_aoi_5_1_inst0_O;
mux_aoi_5_1 mux_aoi_5_1_inst0 (
    .I0(I_0),
    .I1(I_1),
    .I2(I_2),
    .I3(I_3),
    .I4(I_4),
    .S(S),
    .O(mux_aoi_5_1_inst0_O)
);
assign O = mux_aoi_5_1_inst0_O;
endmodule

module MuxWrapperAOIImpl_2_16 (
    input [15:0] I_0,
    input [15:0] I_1,
    output [15:0] O,
    input [0:0] S
);
wire [15:0] mux_aoi_2_16_inst0_O;
mux_aoi_2_16 mux_aoi_2_16_inst0 (
    .I0(I_0),
    .I1(I_1),
    .S(S[0]),
    .O(mux_aoi_2_16_inst0_O)
);
assign O = mux_aoi_2_16_inst0_O;
endmodule

module MuxWrapperAOIImpl_2_1 (
    input [0:0] I_0,
    input [0:0] I_1,
    output [0:0] O,
    input [0:0] S
);
wire [0:0] mux_aoi_2_1_inst0_O;
mux_aoi_2_1 mux_aoi_2_1_inst0 (
    .I0(I_0),
    .I1(I_1),
    .S(S[0]),
    .O(mux_aoi_2_1_inst0_O)
);
assign O = mux_aoi_2_1_inst0_O;
endmodule

module MuxWrapperAOIImpl_20_16 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input [4:0] S
);
wire [15:0] mux_aoi_const_20_16_inst0_O;
mux_aoi_const_20_16 mux_aoi_const_20_16_inst0 (
    .I0(I_0),
    .I1(I_1),
    .I2(I_2),
    .I3(I_3),
    .I4(I_4),
    .I5(I_5),
    .I6(I_6),
    .I7(I_7),
    .I8(I_8),
    .I9(I_9),
    .I10(I_10),
    .I11(I_11),
    .I12(I_12),
    .I13(I_13),
    .I14(I_14),
    .I15(I_15),
    .I16(I_16),
    .I17(I_17),
    .I18(I_18),
    .I19(I_19),
    .S(S),
    .O(mux_aoi_const_20_16_inst0_O)
);
assign O = mux_aoi_const_20_16_inst0_O;
endmodule

module MuxWrapperAOIImpl_20_1 (
    input [0:0] I_0,
    input [0:0] I_1,
    input [0:0] I_10,
    input [0:0] I_11,
    input [0:0] I_12,
    input [0:0] I_13,
    input [0:0] I_14,
    input [0:0] I_15,
    input [0:0] I_16,
    input [0:0] I_17,
    input [0:0] I_18,
    input [0:0] I_19,
    input [0:0] I_2,
    input [0:0] I_3,
    input [0:0] I_4,
    input [0:0] I_5,
    input [0:0] I_6,
    input [0:0] I_7,
    input [0:0] I_8,
    input [0:0] I_9,
    output [0:0] O,
    input [4:0] S
);
wire [0:0] mux_aoi_const_20_1_inst0_O;
mux_aoi_const_20_1 mux_aoi_const_20_1_inst0 (
    .I0(I_0),
    .I1(I_1),
    .I2(I_2),
    .I3(I_3),
    .I4(I_4),
    .I5(I_5),
    .I6(I_6),
    .I7(I_7),
    .I8(I_8),
    .I9(I_9),
    .I10(I_10),
    .I11(I_11),
    .I12(I_12),
    .I13(I_13),
    .I14(I_14),
    .I15(I_15),
    .I16(I_16),
    .I17(I_17),
    .I18(I_18),
    .I19(I_19),
    .S(S),
    .O(mux_aoi_const_20_1_inst0_O)
);
assign O = mux_aoi_const_20_1_inst0_O;
endmodule

module MuxWithDefaultWrapper_15_32_8_0 (
    input [0:0] EN,
    input [31:0] I_0,
    input [31:0] I_1,
    input [31:0] I_10,
    input [31:0] I_11,
    input [31:0] I_12,
    input [31:0] I_13,
    input [31:0] I_14,
    input [31:0] I_2,
    input [31:0] I_3,
    input [31:0] I_4,
    input [31:0] I_5,
    input [31:0] I_6,
    input [31:0] I_7,
    input [31:0] I_8,
    input [31:0] I_9,
    output [31:0] O,
    input [7:0] S
);
wire [31:0] MuxWrapper_15_32_inst0$Mux15xBits32_inst0$coreir_commonlib_mux15x32_inst0_out;
wire [31:0] MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
wire [31:0] const_0_32_out;
wire [7:0] const_15_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_ult_inst0_out;
wire [3:0] MuxWrapper_15_32_inst0$Mux15xBits32_inst0$coreir_commonlib_mux15x32_inst0_in_sel;
assign MuxWrapper_15_32_inst0$Mux15xBits32_inst0$coreir_commonlib_mux15x32_inst0_in_sel = {S[3],S[2],S[1],S[0]};
commonlib_muxn__N15__width32 MuxWrapper_15_32_inst0$Mux15xBits32_inst0$coreir_commonlib_mux15x32_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(MuxWrapper_15_32_inst0$Mux15xBits32_inst0$coreir_commonlib_mux15x32_inst0_in_sel),
    .out(MuxWrapper_15_32_inst0$Mux15xBits32_inst0$coreir_commonlib_mux15x32_inst0_out)
);
coreir_mux #(
    .width(32)
) MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join (
    .in0(const_0_32_out),
    .in1(MuxWrapper_15_32_inst0$Mux15xBits32_inst0$coreir_commonlib_mux15x32_inst0_out),
    .sel(magma_Bit_and_inst0_out),
    .out(MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out)
);
coreir_const #(
    .value(32'h00000000),
    .width(32)
) const_0_32 (
    .out(const_0_32_out)
);
coreir_const #(
    .value(8'h0f),
    .width(8)
) const_15_8 (
    .out(const_15_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_ult_inst0_out),
    .in1(EN[0]),
    .out(magma_Bit_and_inst0_out)
);
coreir_ult #(
    .width(8)
) magma_Bits_8_ult_inst0 (
    .in0(S),
    .in1(const_15_8_out),
    .out(magma_Bits_8_ult_inst0_out)
);
assign O = MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
endmodule

module MuxWithDefaultWrapper_13_32_8_0 (
    input [0:0] EN,
    input [31:0] I_0,
    input [31:0] I_1,
    input [31:0] I_10,
    input [31:0] I_11,
    input [31:0] I_12,
    input [31:0] I_2,
    input [31:0] I_3,
    input [31:0] I_4,
    input [31:0] I_5,
    input [31:0] I_6,
    input [31:0] I_7,
    input [31:0] I_8,
    input [31:0] I_9,
    output [31:0] O,
    input [7:0] S
);
wire [31:0] MuxWrapper_13_32_inst0$Mux13xBits32_inst0$coreir_commonlib_mux13x32_inst0_out;
wire [31:0] MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
wire [31:0] const_0_32_out;
wire [7:0] const_13_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_ult_inst0_out;
wire [3:0] MuxWrapper_13_32_inst0$Mux13xBits32_inst0$coreir_commonlib_mux13x32_inst0_in_sel;
assign MuxWrapper_13_32_inst0$Mux13xBits32_inst0$coreir_commonlib_mux13x32_inst0_in_sel = {S[3],S[2],S[1],S[0]};
commonlib_muxn__N13__width32 MuxWrapper_13_32_inst0$Mux13xBits32_inst0$coreir_commonlib_mux13x32_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(MuxWrapper_13_32_inst0$Mux13xBits32_inst0$coreir_commonlib_mux13x32_inst0_in_sel),
    .out(MuxWrapper_13_32_inst0$Mux13xBits32_inst0$coreir_commonlib_mux13x32_inst0_out)
);
coreir_mux #(
    .width(32)
) MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join (
    .in0(const_0_32_out),
    .in1(MuxWrapper_13_32_inst0$Mux13xBits32_inst0$coreir_commonlib_mux13x32_inst0_out),
    .sel(magma_Bit_and_inst0_out),
    .out(MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out)
);
coreir_const #(
    .value(32'h00000000),
    .width(32)
) const_0_32 (
    .out(const_0_32_out)
);
coreir_const #(
    .value(8'h0d),
    .width(8)
) const_13_8 (
    .out(const_13_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_ult_inst0_out),
    .in1(EN[0]),
    .out(magma_Bit_and_inst0_out)
);
coreir_ult #(
    .width(8)
) magma_Bits_8_ult_inst0 (
    .in0(S),
    .in1(const_13_8_out),
    .out(magma_Bits_8_ult_inst0_out)
);
assign O = MuxWrapper_2_32_inst0$Mux2xBits32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
endmodule

module MUL (
    input [1:0] instr,
    input [0:0] signed_,
    input [15:0] a,
    input [15:0] b,
    output [15:0] O,
    input CLK,
    input ASYNCRESET
);
wire [15:0] Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] const_0_16_out;
wire [1:0] const_0_2_out;
wire [1:0] const_1_2_out;
wire [1:0] const_2_2_out;
wire magma_Bits_2_eq_inst0_out;
wire magma_Bits_2_eq_inst1_out;
wire magma_Bits_2_eq_inst2_out;
wire [31:0] magma_UInt_32_mul_inst0_out;
coreir_mux #(
    .width(16)
) Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(a),
    .in1(const_0_16_out),
    .sel(magma_Bits_2_eq_inst0_out),
    .out(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join (
    .in0(b),
    .in1(const_0_16_out),
    .sel(magma_Bits_2_eq_inst0_out),
    .out(Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_in1 = {magma_UInt_32_mul_inst0_out[23],magma_UInt_32_mul_inst0_out[22],magma_UInt_32_mul_inst0_out[21],magma_UInt_32_mul_inst0_out[20],magma_UInt_32_mul_inst0_out[19],magma_UInt_32_mul_inst0_out[18],magma_UInt_32_mul_inst0_out[17],magma_UInt_32_mul_inst0_out[16],magma_UInt_32_mul_inst0_out[15],magma_UInt_32_mul_inst0_out[14],magma_UInt_32_mul_inst0_out[13],magma_UInt_32_mul_inst0_out[12],magma_UInt_32_mul_inst0_out[11],magma_UInt_32_mul_inst0_out[10],magma_UInt_32_mul_inst0_out[9],magma_UInt_32_mul_inst0_out[8]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join (
    .in0(const_0_16_out),
    .in1(Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_2_eq_inst2_out),
    .out(Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_in1 = {magma_UInt_32_mul_inst0_out[15],magma_UInt_32_mul_inst0_out[14],magma_UInt_32_mul_inst0_out[13],magma_UInt_32_mul_inst0_out[12],magma_UInt_32_mul_inst0_out[11],magma_UInt_32_mul_inst0_out[10],magma_UInt_32_mul_inst0_out[9],magma_UInt_32_mul_inst0_out[8],magma_UInt_32_mul_inst0_out[7],magma_UInt_32_mul_inst0_out[6],magma_UInt_32_mul_inst0_out[5],magma_UInt_32_mul_inst0_out[4],magma_UInt_32_mul_inst0_out[3],magma_UInt_32_mul_inst0_out[2],magma_UInt_32_mul_inst0_out[1],magma_UInt_32_mul_inst0_out[0]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_2_eq_inst1_out),
    .out(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
coreir_const #(
    .value(2'h0),
    .width(2)
) const_0_2 (
    .out(const_0_2_out)
);
coreir_const #(
    .value(2'h1),
    .width(2)
) const_1_2 (
    .out(const_1_2_out)
);
coreir_const #(
    .value(2'h2),
    .width(2)
) const_2_2 (
    .out(const_2_2_out)
);
coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst0 (
    .in0(instr),
    .in1(const_1_2_out),
    .out(magma_Bits_2_eq_inst0_out)
);
coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst1 (
    .in0(instr),
    .in1(const_0_2_out),
    .out(magma_Bits_2_eq_inst1_out)
);
coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst2 (
    .in0(instr),
    .in1(const_2_2_out),
    .out(magma_Bits_2_eq_inst2_out)
);
wire [31:0] magma_UInt_32_mul_inst0_in0;
assign magma_UInt_32_mul_inst0_in0 = {Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out};
wire [31:0] magma_UInt_32_mul_inst0_in1;
assign magma_UInt_32_mul_inst0_in1 = {Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15],Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out};
coreir_mul #(
    .width(32)
) magma_UInt_32_mul_inst0 (
    .in0(magma_UInt_32_mul_inst0_in0),
    .in1(magma_UInt_32_mul_inst0_in1),
    .out(magma_UInt_32_mul_inst0_out)
);
assign O = Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out;
endmodule

module Chain (
  input logic [1:0] accessor_output,
  input logic [1:0] [15:0] chain_data_in,
  input logic chain_en,
  input logic clk_en,
  input logic [1:0] [15:0] curr_tile_data_out,
  input logic flush,
  output logic [1:0] [15:0] data_out_tile
);

always_comb begin
  if (accessor_output[0]) begin
    data_out_tile[0] = curr_tile_data_out[0];
  end
  else if (chain_en) begin
    data_out_tile[0] = chain_data_in[0];
  end
  else data_out_tile[0] = 16'h0;
  if (accessor_output[1]) begin
    data_out_tile[1] = curr_tile_data_out[1];
  end
  else if (chain_en) begin
    data_out_tile[1] = chain_data_in[1];
  end
  else data_out_tile[1] = 16'h0;
end
endmodule   // Chain

module IN12LP_S1DB_W00512B032M04S2_H_2_wide_1_deep (
  input logic [8:0] A,
  input logic CEN,
  input logic CLK,
  input logic [63:0] D,
  input logic MA_SAWL0,
  input logic MA_SAWL1,
  input logic MA_STABAS0,
  input logic MA_STABAS1,
  input logic MA_VD0,
  input logic MA_VD1,
  input logic MA_WL0,
  input logic MA_WL1,
  input logic MA_WRAS0,
  input logic MA_WRAS1,
  input logic MA_WRT,
  input logic RDWEN,
  input logic T_LOGIC,
  input logic T_Q_RST,
  input logic clk_en,
  input logic flush,
  output logic [63:0] Q
);

logic [31:0] IN12LP_S1DB_W00512B032M04S2_H_0_0_D;
logic [31:0] IN12LP_S1DB_W00512B032M04S2_H_0_0_Q;
logic [31:0] IN12LP_S1DB_W00512B032M04S2_H_1_0_D;
logic [31:0] IN12LP_S1DB_W00512B032M04S2_H_1_0_Q;
assign {IN12LP_S1DB_W00512B032M04S2_H_0_0_D, IN12LP_S1DB_W00512B032M04S2_H_1_0_D} = D;
assign Q = {IN12LP_S1DB_W00512B032M04S2_H_0_0_Q, IN12LP_S1DB_W00512B032M04S2_H_1_0_Q};
IN12LP_S1DB_W00512B032M04S2_H IN12LP_S1DB_W00512B032M04S2_H_0_0 (
  .A(A),
  .CEN(CEN),
  .CLK(CLK),
  .D(IN12LP_S1DB_W00512B032M04S2_H_0_0_D),
  .MA_SAWL0(MA_SAWL0),
  .MA_SAWL1(MA_SAWL1),
  .MA_STABAS0(MA_STABAS0),
  .MA_STABAS1(MA_STABAS1),
  .MA_VD0(MA_VD0),
  .MA_VD1(MA_VD1),
  .MA_WL0(MA_WL0),
  .MA_WL1(MA_WL1),
  .MA_WRAS0(MA_WRAS0),
  .MA_WRAS1(MA_WRAS1),
  .MA_WRT(MA_WRT),
  .RDWEN(RDWEN),
  .T_LOGIC(T_LOGIC),
  .T_Q_RST(T_Q_RST),
  .Q(IN12LP_S1DB_W00512B032M04S2_H_0_0_Q)
);

IN12LP_S1DB_W00512B032M04S2_H IN12LP_S1DB_W00512B032M04S2_H_1_0 (
  .A(A),
  .CEN(CEN),
  .CLK(CLK),
  .D(IN12LP_S1DB_W00512B032M04S2_H_1_0_D),
  .MA_SAWL0(MA_SAWL0),
  .MA_SAWL1(MA_SAWL1),
  .MA_STABAS0(MA_STABAS0),
  .MA_STABAS1(MA_STABAS1),
  .MA_VD0(MA_VD0),
  .MA_VD1(MA_VD1),
  .MA_WL0(MA_WL0),
  .MA_WL1(MA_WL1),
  .MA_WRAS0(MA_WRAS0),
  .MA_WRAS1(MA_WRAS1),
  .MA_WRT(MA_WRT),
  .RDWEN(RDWEN),
  .T_LOGIC(T_LOGIC),
  .T_Q_RST(T_Q_RST),
  .Q(IN12LP_S1DB_W00512B032M04S2_H_1_0_Q)
);

endmodule   // IN12LP_S1DB_W00512B032M04S2_H_2_wide_1_deep

module LakeTop (
  input logic clk,
  input logic clk_en,
  input logic [7:0] config_addr_in,
  input logic [31:0] config_data_in,
  input logic [1:0] config_en,
  input logic config_read,
  input logic config_write,
  input logic flush,
  input logic [0:0] [15:0] input_width_16_num_0,
  input logic [0:0] [15:0] input_width_16_num_1,
  input logic [0:0] [15:0] input_width_16_num_2,
  input logic [0:0] [15:0] input_width_16_num_3,
  input logic input_width_1_num_0,
  input logic input_width_1_num_1,
  input logic [3:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality,
  input logic [5:0] [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges,
  input logic mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable,
  input logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides,
  input logic [15:0] mem_ctrl_strg_fifo_flat_strg_fifo_inst_fifo_depth,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides,
  input logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides,
  input logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality,
  input logic [5:0] [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality,
  input logic [5:0] [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges,
  input logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides,
  input logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality,
  input logic [5:0] [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality,
  input logic [5:0] [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges,
  input logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr,
  input logic [5:0] [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr,
  input logic [5:0] [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr,
  input logic [5:0] [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr,
  input logic [5:0] [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality,
  input logic [5:0] [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality,
  input logic [5:0] [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges,
  input logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides,
  input logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality,
  input logic [5:0] [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality,
  input logic [5:0] [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides,
  input logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides,
  input logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides,
  input logic [1:0] mode,
  input logic rst_n,
  input logic tile_en,
  output logic [1:0] [31:0] config_data_out,
  output logic [0:0] [15:0] output_width_16_num_0,
  output logic [0:0] [15:0] output_width_16_num_1,
  output logic output_width_1_num_0,
  output logic output_width_1_num_1,
  output logic output_width_1_num_2,
  output logic output_width_1_num_3
);

logic [15:0] config_data_in_shrt;
logic [1:0][15:0] config_data_out_shrt;
logic [8:0] config_seq_addr_out;
logic config_seq_clk;
logic config_seq_clk_en;
logic [0:0][3:0][15:0] config_seq_rd_data_stg;
logic config_seq_ren_out;
logic config_seq_wen_out;
logic [3:0][15:0] config_seq_wr_data;
logic gclk;
logic mem_ctrl_stencil_valid_flat_clk;
logic mem_ctrl_stencil_valid_flat_stencil_valid_f_;
logic [0:0][8:0] mem_ctrl_strg_fifo_flat_addr_out_lifted;
logic mem_ctrl_strg_fifo_flat_clk;
logic [0:0][3:0][15:0] mem_ctrl_strg_fifo_flat_data_from_strg_lifted;
logic [0:0][15:0] mem_ctrl_strg_fifo_flat_data_out_f_;
logic [0:0][3:0][15:0] mem_ctrl_strg_fifo_flat_data_to_strg_lifted;
logic mem_ctrl_strg_fifo_flat_empty_f_;
logic mem_ctrl_strg_fifo_flat_full_f_;
logic mem_ctrl_strg_fifo_flat_ren_to_strg_lifted;
logic mem_ctrl_strg_fifo_flat_valid_out_f_;
logic mem_ctrl_strg_fifo_flat_wen_to_strg_lifted;
logic [0:0][8:0] mem_ctrl_strg_ram_flat_addr_out_lifted;
logic mem_ctrl_strg_ram_flat_clk;
logic [0:0][3:0][15:0] mem_ctrl_strg_ram_flat_data_from_strg_lifted;
logic [0:0][15:0] mem_ctrl_strg_ram_flat_data_out_f_;
logic [0:0][3:0][15:0] mem_ctrl_strg_ram_flat_data_to_strg_lifted;
logic mem_ctrl_strg_ram_flat_ready_f_;
logic mem_ctrl_strg_ram_flat_ren_to_strg_lifted;
logic mem_ctrl_strg_ram_flat_valid_out_f_;
logic mem_ctrl_strg_ram_flat_wen_to_strg_lifted;
logic mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_0;
logic mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_1;
logic [8:0] mem_ctrl_strg_ub_vec_flat_addr_out_lifted;
logic mem_ctrl_strg_ub_vec_flat_clk;
logic [3:0][15:0] mem_ctrl_strg_ub_vec_flat_data_from_strg_lifted;
logic [0:0][15:0] mem_ctrl_strg_ub_vec_flat_data_out_f_0;
logic [0:0][15:0] mem_ctrl_strg_ub_vec_flat_data_out_f_1;
logic [3:0][15:0] mem_ctrl_strg_ub_vec_flat_data_to_strg_lifted;
logic mem_ctrl_strg_ub_vec_flat_ren_to_strg_lifted;
logic mem_ctrl_strg_ub_vec_flat_wen_to_strg_lifted;
logic memory_0_clk;
logic memory_0_clk_en;
logic [63:0] memory_0_data_in_p0;
logic [63:0] memory_0_data_out_p0;
logic [8:0] memory_0_read_addr_p0;
logic memory_0_read_enable_p0;
logic [8:0] memory_0_write_addr_p0;
logic memory_0_write_enable_p0;
assign gclk = clk & tile_en;
assign mem_ctrl_strg_ub_vec_flat_clk = gclk & (mode == 2'h0);
assign mem_ctrl_strg_fifo_flat_clk = gclk & (mode == 2'h1);
assign mem_ctrl_strg_ram_flat_clk = gclk & (mode == 2'h2);
assign mem_ctrl_stencil_valid_flat_clk = gclk;
always_comb begin
  output_width_16_num_0 = 16'h0;
  if (mode == 2'h0) begin
    output_width_16_num_0 = mem_ctrl_strg_ub_vec_flat_data_out_f_0;
  end
  else if (mode == 2'h1) begin
    output_width_16_num_0 = mem_ctrl_strg_fifo_flat_data_out_f_;
  end
  else if (mode == 2'h2) begin
    output_width_16_num_0 = mem_ctrl_strg_ram_flat_data_out_f_;
  end
end
always_comb begin
  output_width_16_num_1 = 16'h0;
  output_width_16_num_1 = mem_ctrl_strg_ub_vec_flat_data_out_f_1;
end
always_comb begin
  output_width_1_num_0 = 1'h0;
  if (mode == 2'h0) begin
    output_width_1_num_0 = mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_0;
  end
  else if (mode == 2'h1) begin
    output_width_1_num_0 = mem_ctrl_strg_fifo_flat_empty_f_;
  end
  else if (mode == 2'h2) begin
    output_width_1_num_0 = mem_ctrl_strg_ram_flat_ready_f_;
  end
end
always_comb begin
  output_width_1_num_1 = 1'h0;
  if (mode == 2'h0) begin
    output_width_1_num_1 = mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_1;
  end
  else if (mode == 2'h1) begin
    output_width_1_num_1 = mem_ctrl_strg_fifo_flat_full_f_;
  end
  else if (mode == 2'h2) begin
    output_width_1_num_1 = mem_ctrl_strg_ram_flat_valid_out_f_;
  end
end
always_comb begin
  output_width_1_num_2 = 1'h0;
  output_width_1_num_2 = mem_ctrl_strg_fifo_flat_valid_out_f_;
end
always_comb begin
  output_width_1_num_3 = 1'h0;
  output_width_1_num_3 = mem_ctrl_stencil_valid_flat_stencil_valid_f_;
end
assign memory_0_clk = gclk;
always_comb begin
  memory_0_data_in_p0 = 64'h0;
  memory_0_write_addr_p0 = 9'h0;
  memory_0_write_enable_p0 = 1'h0;
  memory_0_read_addr_p0 = 9'h0;
  memory_0_read_enable_p0 = 1'h0;
  if (|config_en) begin
    memory_0_data_in_p0 = config_seq_wr_data;
    memory_0_write_addr_p0 = config_seq_addr_out;
    memory_0_write_enable_p0 = config_seq_wen_out;
    memory_0_read_addr_p0 = config_seq_addr_out;
    memory_0_read_enable_p0 = config_seq_ren_out;
  end
  else if (mode == 2'h0) begin
    memory_0_data_in_p0 = mem_ctrl_strg_ub_vec_flat_data_to_strg_lifted;
    memory_0_write_addr_p0 = mem_ctrl_strg_ub_vec_flat_addr_out_lifted;
    memory_0_write_enable_p0 = mem_ctrl_strg_ub_vec_flat_wen_to_strg_lifted;
    memory_0_read_addr_p0 = mem_ctrl_strg_ub_vec_flat_addr_out_lifted;
    memory_0_read_enable_p0 = mem_ctrl_strg_ub_vec_flat_ren_to_strg_lifted;
  end
  else if (mode == 2'h1) begin
    memory_0_data_in_p0 = mem_ctrl_strg_fifo_flat_data_to_strg_lifted;
    memory_0_write_addr_p0 = mem_ctrl_strg_fifo_flat_addr_out_lifted;
    memory_0_write_enable_p0 = mem_ctrl_strg_fifo_flat_wen_to_strg_lifted;
    memory_0_read_addr_p0 = mem_ctrl_strg_fifo_flat_addr_out_lifted;
    memory_0_read_enable_p0 = mem_ctrl_strg_fifo_flat_ren_to_strg_lifted;
  end
  else if (mode == 2'h2) begin
    memory_0_data_in_p0 = mem_ctrl_strg_ram_flat_data_to_strg_lifted;
    memory_0_write_addr_p0 = mem_ctrl_strg_ram_flat_addr_out_lifted;
    memory_0_write_enable_p0 = mem_ctrl_strg_ram_flat_wen_to_strg_lifted;
    memory_0_read_addr_p0 = mem_ctrl_strg_ram_flat_addr_out_lifted;
    memory_0_read_enable_p0 = mem_ctrl_strg_ram_flat_ren_to_strg_lifted;
  end
end
always_comb begin
  mem_ctrl_strg_ub_vec_flat_data_from_strg_lifted = memory_0_data_out_p0;
  mem_ctrl_strg_fifo_flat_data_from_strg_lifted = memory_0_data_out_p0;
  mem_ctrl_strg_ram_flat_data_from_strg_lifted = memory_0_data_out_p0;
  config_seq_rd_data_stg = memory_0_data_out_p0;
end
assign config_data_in_shrt = config_data_in[15:0];
assign config_data_out[0] = 32'(config_data_out_shrt[0]);
assign config_data_out[1] = 32'(config_data_out_shrt[1]);
assign config_seq_clk = gclk;
assign config_seq_clk_en = clk_en | (|config_en);
assign memory_0_clk_en = clk_en | (|config_en);
strg_ub_vec_flat mem_ctrl_strg_ub_vec_flat (
  .chain_data_in_f_0(input_width_16_num_0),
  .chain_data_in_f_1(input_width_16_num_1),
  .clk(mem_ctrl_strg_ub_vec_flat_clk),
  .clk_en(clk_en),
  .data_from_strg_lifted(mem_ctrl_strg_ub_vec_flat_data_from_strg_lifted),
  .data_in_f_0(input_width_16_num_2),
  .data_in_f_1(input_width_16_num_3),
  .flush(flush),
  .rst_n(rst_n),
  .strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr),
  .strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides),
  .strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr),
  .strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides),
  .strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr),
  .strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides),
  .strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr),
  .strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides),
  .strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable),
  .strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr),
  .strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides),
  .strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable),
  .strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr),
  .strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides),
  .strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality),
  .strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges),
  .strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality),
  .strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges),
  .strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable),
  .strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr),
  .strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides),
  .strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable),
  .strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr),
  .strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides),
  .strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality),
  .strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges),
  .strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality),
  .strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges),
  .strg_ub_vec_inst_chain_chain_en(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en),
  .strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr),
  .strg_ub_vec_inst_sram_only_input_addr_gen_0_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides),
  .strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr),
  .strg_ub_vec_inst_sram_only_input_addr_gen_1_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides),
  .strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr),
  .strg_ub_vec_inst_sram_only_output_addr_gen_0_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides),
  .strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr),
  .strg_ub_vec_inst_sram_only_output_addr_gen_1_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides),
  .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality),
  .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges),
  .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality),
  .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides),
  .strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality),
  .strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges),
  .strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality),
  .strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges),
  .strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr),
  .strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides),
  .strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr),
  .strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides),
  .strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr),
  .strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides),
  .strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr),
  .strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides),
  .accessor_output_f_b_0(mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_0),
  .accessor_output_f_b_1(mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_1),
  .addr_out_lifted(mem_ctrl_strg_ub_vec_flat_addr_out_lifted),
  .data_out_f_0(mem_ctrl_strg_ub_vec_flat_data_out_f_0),
  .data_out_f_1(mem_ctrl_strg_ub_vec_flat_data_out_f_1),
  .data_to_strg_lifted(mem_ctrl_strg_ub_vec_flat_data_to_strg_lifted),
  .ren_to_strg_lifted(mem_ctrl_strg_ub_vec_flat_ren_to_strg_lifted),
  .wen_to_strg_lifted(mem_ctrl_strg_ub_vec_flat_wen_to_strg_lifted)
);

strg_fifo_flat mem_ctrl_strg_fifo_flat (
  .clk(mem_ctrl_strg_fifo_flat_clk),
  .clk_en(clk_en),
  .data_from_strg_lifted(mem_ctrl_strg_fifo_flat_data_from_strg_lifted),
  .data_in_f_(input_width_16_num_0),
  .flush(flush),
  .pop_f_(input_width_1_num_0),
  .push_f_(input_width_1_num_1),
  .rst_n(rst_n),
  .strg_fifo_inst_fifo_depth(mem_ctrl_strg_fifo_flat_strg_fifo_inst_fifo_depth),
  .addr_out_lifted(mem_ctrl_strg_fifo_flat_addr_out_lifted),
  .data_out_f_(mem_ctrl_strg_fifo_flat_data_out_f_),
  .data_to_strg_lifted(mem_ctrl_strg_fifo_flat_data_to_strg_lifted),
  .empty_f_(mem_ctrl_strg_fifo_flat_empty_f_),
  .full_f_(mem_ctrl_strg_fifo_flat_full_f_),
  .ren_to_strg_lifted(mem_ctrl_strg_fifo_flat_ren_to_strg_lifted),
  .valid_out_f_(mem_ctrl_strg_fifo_flat_valid_out_f_),
  .wen_to_strg_lifted(mem_ctrl_strg_fifo_flat_wen_to_strg_lifted)
);

strg_ram_flat mem_ctrl_strg_ram_flat (
  .clk(mem_ctrl_strg_ram_flat_clk),
  .clk_en(clk_en),
  .data_from_strg_lifted(mem_ctrl_strg_ram_flat_data_from_strg_lifted),
  .data_in_f_(input_width_16_num_0),
  .flush(flush),
  .rd_addr_in_f_(input_width_16_num_1),
  .ren_f_(input_width_1_num_0),
  .rst_n(rst_n),
  .wen_f_(input_width_1_num_1),
  .wr_addr_in_f_(input_width_16_num_2),
  .addr_out_lifted(mem_ctrl_strg_ram_flat_addr_out_lifted),
  .data_out_f_(mem_ctrl_strg_ram_flat_data_out_f_),
  .data_to_strg_lifted(mem_ctrl_strg_ram_flat_data_to_strg_lifted),
  .ready_f_(mem_ctrl_strg_ram_flat_ready_f_),
  .ren_to_strg_lifted(mem_ctrl_strg_ram_flat_ren_to_strg_lifted),
  .valid_out_f_(mem_ctrl_strg_ram_flat_valid_out_f_),
  .wen_to_strg_lifted(mem_ctrl_strg_ram_flat_wen_to_strg_lifted)
);

stencil_valid_flat mem_ctrl_stencil_valid_flat (
  .clk(mem_ctrl_stencil_valid_flat_clk),
  .clk_en(clk_en),
  .flush(flush),
  .rst_n(rst_n),
  .stencil_valid_inst_loops_stencil_valid_dimensionality(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality),
  .stencil_valid_inst_loops_stencil_valid_ranges(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges),
  .stencil_valid_inst_stencil_valid_sched_gen_enable(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable),
  .stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr),
  .stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides),
  .stencil_valid_f_(mem_ctrl_stencil_valid_flat_stencil_valid_f_)
);

sram_sp__0 memory_0 (
  .clk(memory_0_clk),
  .clk_en(memory_0_clk_en),
  .data_in_p0(memory_0_data_in_p0),
  .flush(flush),
  .read_addr_p0(memory_0_read_addr_p0),
  .read_enable_p0(memory_0_read_enable_p0),
  .write_addr_p0(memory_0_write_addr_p0),
  .write_enable_p0(memory_0_write_enable_p0),
  .data_out_p0(memory_0_data_out_p0)
);

storage_config_seq_unq0 config_seq (
  .clk(config_seq_clk),
  .clk_en(config_seq_clk_en),
  .config_addr_in(config_addr_in),
  .config_data_in(config_data_in_shrt),
  .config_en(config_en),
  .config_rd(config_read),
  .config_wr(config_write),
  .flush(flush),
  .rd_data_stg(config_seq_rd_data_stg),
  .rst_n(rst_n),
  .addr_out(config_seq_addr_out),
  .rd_data_out(config_data_out_shrt),
  .ren_out(config_seq_ren_out),
  .wen_out(config_seq_wen_out),
  .wr_data(config_seq_wr_data)
);

endmodule   // LakeTop

module LakeTop_W (
  input logic clk,
  input logic clk_en,
  input logic [7:0] config_addr_in,
  input logic [31:0] config_data_in,
  input logic [1:0] config_en,
  input logic config_read,
  input logic config_write,
  input logic flush,
  input logic [0:0] [15:0] input_width_16_num_0,
  input logic [0:0] [15:0] input_width_16_num_1,
  input logic [0:0] [15:0] input_width_16_num_2,
  input logic [0:0] [15:0] input_width_16_num_3,
  input logic input_width_1_num_0,
  input logic input_width_1_num_1,
  input logic [3:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality,
  input logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0,
  input logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1,
  input logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2,
  input logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3,
  input logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4,
  input logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5,
  input logic mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable,
  input logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr,
  input logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0,
  input logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1,
  input logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2,
  input logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3,
  input logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4,
  input logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5,
  input logic [15:0] mem_ctrl_strg_fifo_flat_strg_fifo_inst_fifo_depth,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5,
  input logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5,
  input logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5,
  input logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5,
  input logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5,
  input logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4,
  input logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5,
  input logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5,
  input logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5,
  input logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5,
  input logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4,
  input logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4,
  input logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5,
  input logic [1:0] mode,
  input logic rst_n,
  input logic tile_en,
  output logic [31:0] config_data_out_0,
  output logic [31:0] config_data_out_1,
  output logic [0:0] [15:0] output_width_16_num_0,
  output logic [0:0] [15:0] output_width_16_num_1,
  output logic output_width_1_num_0,
  output logic output_width_1_num_1,
  output logic output_width_1_num_2,
  output logic output_width_1_num_3
);

logic [1:0][31:0] LakeTop_config_data_out;
logic [5:0][15:0] LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges;
logic [5:0][15:0] LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides;
logic [5:0][3:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides;
logic [5:0][3:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides;
logic [5:0][3:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides;
logic [5:0][3:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides;
logic [5:0][15:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides;
logic [5:0][15:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides;
logic [5:0][15:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges;
logic [5:0][15:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges;
logic [5:0][15:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides;
logic [5:0][15:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides;
logic [5:0][15:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges;
logic [5:0][15:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges;
logic [5:0][8:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides;
logic [5:0][8:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides;
logic [5:0][8:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides;
logic [5:0][8:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides;
logic [5:0][15:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges;
logic [5:0][15:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges;
logic [5:0][15:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides;
logic [5:0][15:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides;
logic [5:0][15:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges;
logic [5:0][15:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges;
logic [5:0][3:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides;
logic [5:0][3:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides;
logic [5:0][15:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides;
logic [5:0][15:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides;
logic [5:0][3:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides;
logic [5:0][3:0] LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides;
assign config_data_out_0 = LakeTop_config_data_out[0];
assign config_data_out_1 = LakeTop_config_data_out[1];
assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges[0] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0;
assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges[1] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1;
assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges[2] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2;
assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges[3] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3;
assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges[4] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4;
assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges[5] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5;
assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides[0] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0;
assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides[1] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1;
assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides[2] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2;
assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides[3] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3;
assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides[4] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4;
assign LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides[5] = mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides[0] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides[1] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides[2] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides[3] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides[4] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4;
assign LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides[5] = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5;
LakeTop LakeTop (
  .clk(clk),
  .clk_en(clk_en),
  .config_addr_in(config_addr_in),
  .config_data_in(config_data_in),
  .config_en(config_en),
  .config_read(config_read),
  .config_write(config_write),
  .flush(flush),
  .input_width_16_num_0(input_width_16_num_0),
  .input_width_16_num_1(input_width_16_num_1),
  .input_width_16_num_2(input_width_16_num_2),
  .input_width_16_num_3(input_width_16_num_3),
  .input_width_1_num_0(input_width_1_num_0),
  .input_width_1_num_1(input_width_1_num_1),
  .mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality),
  .mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges(LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges),
  .mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable),
  .mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr),
  .mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides(LakeTop_mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides),
  .mem_ctrl_strg_fifo_flat_strg_fifo_inst_fifo_depth(mem_ctrl_strg_fifo_flat_strg_fifo_inst_fifo_depth),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr),
  .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides(LakeTop_mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides),
  .mode(mode),
  .rst_n(rst_n),
  .tile_en(tile_en),
  .config_data_out(LakeTop_config_data_out),
  .output_width_16_num_0(output_width_16_num_0),
  .output_width_16_num_1(output_width_16_num_1),
  .output_width_1_num_0(output_width_1_num_0),
  .output_width_1_num_1(output_width_1_num_1),
  .output_width_1_num_2(output_width_1_num_2),
  .output_width_1_num_3(output_width_1_num_3)
);

endmodule   // LakeTop_W

module addr_gen_6_16 (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [2:0] mux_sel,
  input logic restart,
  input logic rst_n,
  input logic [15:0] starting_addr,
  input logic step,
  input logic [5:0] [15:0] strides,
  output logic [15:0] addr_out
);

logic [15:0] calc_addr;
logic [15:0] current_addr;
logic [15:0] strt_addr;
assign strt_addr = starting_addr;
assign addr_out = calc_addr;
assign calc_addr = strt_addr + current_addr;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    current_addr <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      current_addr <= 16'h0;
    end
    else if (step) begin
      if (restart) begin
        current_addr <= 16'h0;
      end
      else current_addr <= current_addr + strides[mux_sel];
    end
  end
end
endmodule   // addr_gen_6_16

module addr_gen_6_4 (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [2:0] mux_sel,
  input logic restart,
  input logic rst_n,
  input logic [3:0] starting_addr,
  input logic step,
  input logic [5:0] [3:0] strides,
  output logic [3:0] addr_out
);

logic [3:0] calc_addr;
logic [3:0] current_addr;
logic [3:0] strt_addr;
assign strt_addr = starting_addr;
assign addr_out = calc_addr;
assign calc_addr = strt_addr + current_addr;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    current_addr <= 4'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      current_addr <= 4'h0;
    end
    else if (step) begin
      if (restart) begin
        current_addr <= 4'h0;
      end
      else current_addr <= current_addr + strides[mux_sel];
    end
  end
end
endmodule   // addr_gen_6_4

module addr_gen_6_9 (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [2:0] mux_sel,
  input logic restart,
  input logic rst_n,
  input logic [8:0] starting_addr,
  input logic step,
  input logic [5:0] [8:0] strides,
  output logic [8:0] addr_out
);

logic [8:0] calc_addr;
logic [8:0] current_addr;
logic [8:0] strt_addr;
assign strt_addr = starting_addr;
assign addr_out = calc_addr;
assign calc_addr = strt_addr + current_addr;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    current_addr <= 9'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      current_addr <= 9'h0;
    end
    else if (step) begin
      if (restart) begin
        current_addr <= 9'h0;
      end
      else current_addr <= current_addr + strides[mux_sel];
    end
  end
end
endmodule   // addr_gen_6_9

module for_loop_6_16 #(
  parameter CONFIG_WIDTH = 5'h10,
  parameter ITERATOR_SUPPORT = 4'h6
)
(
  input logic clk,
  input logic clk_en,
  input logic [3:0] dimensionality,
  input logic flush,
  input logic [5:0] [15:0] ranges,
  input logic rst_n,
  input logic step,
  output logic [2:0] mux_sel_out,
  output logic restart
);

logic [5:0] clear;
logic [5:0][15:0] dim_counter;
logic done;
logic [5:0] inc;
logic [15:0] inced_cnt;
logic [5:0] max_value;
logic maxed_value;
logic [2:0] mux_sel;
assign mux_sel_out = mux_sel;
assign inced_cnt = dim_counter[mux_sel] + 16'h1;
assign maxed_value = (dim_counter[mux_sel] == ranges[mux_sel]) & inc[mux_sel];
always_comb begin
  mux_sel = 3'h0;
  done = 1'h0;
  if (~done) begin
    if ((~max_value[0]) & (dimensionality > 4'h0)) begin
      mux_sel = 3'h0;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[1]) & (dimensionality > 4'h1)) begin
      mux_sel = 3'h1;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[2]) & (dimensionality > 4'h2)) begin
      mux_sel = 3'h2;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[3]) & (dimensionality > 4'h3)) begin
      mux_sel = 3'h3;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[4]) & (dimensionality > 4'h4)) begin
      mux_sel = 3'h4;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[5]) & (dimensionality > 4'h5)) begin
      mux_sel = 3'h5;
      done = 1'h1;
    end
  end
end
always_comb begin
  clear[0] = 1'h0;
  if (((mux_sel > 3'h0) | (~done)) & step) begin
    clear[0] = 1'h1;
  end
end
always_comb begin
  inc[0] = 1'h0;
  if ((5'h0 == 5'h0) & step & (dimensionality > 4'h0)) begin
    inc[0] = 1'h1;
  end
  else if ((mux_sel == 3'h0) & step & (dimensionality > 4'h0)) begin
    inc[0] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[0] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[0] <= 16'h0;
    end
    else if (clear[0]) begin
      dim_counter[0] <= 16'h0;
    end
    else if (inc[0]) begin
      dim_counter[0] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[0] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[0] <= 1'h0;
    end
    else if (clear[0]) begin
      max_value[0] <= 1'h0;
    end
    else if (inc[0]) begin
      max_value[0] <= maxed_value;
    end
  end
end
always_comb begin
  clear[1] = 1'h0;
  if (((mux_sel > 3'h1) | (~done)) & step) begin
    clear[1] = 1'h1;
  end
end
always_comb begin
  inc[1] = 1'h0;
  if ((5'h1 == 5'h0) & step & (dimensionality > 4'h1)) begin
    inc[1] = 1'h1;
  end
  else if ((mux_sel == 3'h1) & step & (dimensionality > 4'h1)) begin
    inc[1] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[1] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[1] <= 16'h0;
    end
    else if (clear[1]) begin
      dim_counter[1] <= 16'h0;
    end
    else if (inc[1]) begin
      dim_counter[1] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[1] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[1] <= 1'h0;
    end
    else if (clear[1]) begin
      max_value[1] <= 1'h0;
    end
    else if (inc[1]) begin
      max_value[1] <= maxed_value;
    end
  end
end
always_comb begin
  clear[2] = 1'h0;
  if (((mux_sel > 3'h2) | (~done)) & step) begin
    clear[2] = 1'h1;
  end
end
always_comb begin
  inc[2] = 1'h0;
  if ((5'h2 == 5'h0) & step & (dimensionality > 4'h2)) begin
    inc[2] = 1'h1;
  end
  else if ((mux_sel == 3'h2) & step & (dimensionality > 4'h2)) begin
    inc[2] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[2] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[2] <= 16'h0;
    end
    else if (clear[2]) begin
      dim_counter[2] <= 16'h0;
    end
    else if (inc[2]) begin
      dim_counter[2] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[2] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[2] <= 1'h0;
    end
    else if (clear[2]) begin
      max_value[2] <= 1'h0;
    end
    else if (inc[2]) begin
      max_value[2] <= maxed_value;
    end
  end
end
always_comb begin
  clear[3] = 1'h0;
  if (((mux_sel > 3'h3) | (~done)) & step) begin
    clear[3] = 1'h1;
  end
end
always_comb begin
  inc[3] = 1'h0;
  if ((5'h3 == 5'h0) & step & (dimensionality > 4'h3)) begin
    inc[3] = 1'h1;
  end
  else if ((mux_sel == 3'h3) & step & (dimensionality > 4'h3)) begin
    inc[3] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[3] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[3] <= 16'h0;
    end
    else if (clear[3]) begin
      dim_counter[3] <= 16'h0;
    end
    else if (inc[3]) begin
      dim_counter[3] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[3] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[3] <= 1'h0;
    end
    else if (clear[3]) begin
      max_value[3] <= 1'h0;
    end
    else if (inc[3]) begin
      max_value[3] <= maxed_value;
    end
  end
end
always_comb begin
  clear[4] = 1'h0;
  if (((mux_sel > 3'h4) | (~done)) & step) begin
    clear[4] = 1'h1;
  end
end
always_comb begin
  inc[4] = 1'h0;
  if ((5'h4 == 5'h0) & step & (dimensionality > 4'h4)) begin
    inc[4] = 1'h1;
  end
  else if ((mux_sel == 3'h4) & step & (dimensionality > 4'h4)) begin
    inc[4] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[4] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[4] <= 16'h0;
    end
    else if (clear[4]) begin
      dim_counter[4] <= 16'h0;
    end
    else if (inc[4]) begin
      dim_counter[4] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[4] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[4] <= 1'h0;
    end
    else if (clear[4]) begin
      max_value[4] <= 1'h0;
    end
    else if (inc[4]) begin
      max_value[4] <= maxed_value;
    end
  end
end
always_comb begin
  clear[5] = 1'h0;
  if (((mux_sel > 3'h5) | (~done)) & step) begin
    clear[5] = 1'h1;
  end
end
always_comb begin
  inc[5] = 1'h0;
  if ((5'h5 == 5'h0) & step & (dimensionality > 4'h5)) begin
    inc[5] = 1'h1;
  end
  else if ((mux_sel == 3'h5) & step & (dimensionality > 4'h5)) begin
    inc[5] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[5] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[5] <= 16'h0;
    end
    else if (clear[5]) begin
      dim_counter[5] <= 16'h0;
    end
    else if (inc[5]) begin
      dim_counter[5] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[5] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[5] <= 1'h0;
    end
    else if (clear[5]) begin
      max_value[5] <= 1'h0;
    end
    else if (inc[5]) begin
      max_value[5] <= maxed_value;
    end
  end
end
assign restart = step & (~done);
endmodule   // for_loop_6_16

module reg_fifo_d_4_w_1 #(
  parameter data_width = 16'h10
)
(
  input logic clk,
  input logic clk_en,
  input logic [0:0] [data_width-1:0] data_in,
  input logic flush,
  input logic [2:0] num_load,
  input logic [3:0][0:0] [data_width-1:0] parallel_in,
  input logic parallel_load,
  input logic parallel_read,
  input logic pop,
  input logic push,
  input logic rst_n,
  output logic [0:0] [data_width-1:0] data_out,
  output logic empty,
  output logic full,
  output logic [3:0][0:0] [data_width-1:0] parallel_out,
  output logic [1:0] rd_ptr_out,
  output logic valid
);

logic [2:0] num_items;
logic passthru;
logic [1:0] rd_ptr;
logic read;
logic [3:0][0:0][data_width-1:0] reg_array;
logic [1:0] wr_ptr;
logic write;
assign rd_ptr_out = rd_ptr;
assign full = num_items == 3'h4;
assign empty = num_items == 3'h0;
assign read = pop & (~passthru) & (~empty);
assign passthru = pop & push & empty;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_items <= 3'h0;
  end
  else if (flush) begin
    num_items <= 3'h0;
  end
  else if (clk_en) begin
    if (parallel_load) begin
      if (num_load == 3'h0) begin
        num_items <= 3'(push);
      end
      else num_items <= num_load;
    end
    else if (parallel_read) begin
      if (push) begin
        num_items <= 3'h1;
      end
      else num_items <= 3'h0;
    end
    else if (write & (~read)) begin
      num_items <= num_items + 3'h1;
    end
    else if ((~write) & read) begin
      num_items <= num_items - 3'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    reg_array <= 64'h0;
  end
  else if (flush) begin
    reg_array <= 64'h0;
  end
  else if (clk_en) begin
    if (parallel_load) begin
      reg_array <= parallel_in;
    end
    else if (write) begin
      if (parallel_read) begin
        reg_array[0] <= data_in;
      end
      else reg_array[wr_ptr] <= data_in;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    wr_ptr <= 2'h0;
  end
  else if (flush) begin
    wr_ptr <= 2'h0;
  end
  else if (clk_en) begin
    if (parallel_load) begin
      wr_ptr <= num_load[1:0];
    end
    else if (parallel_read) begin
      if (push) begin
        wr_ptr <= 2'h1;
      end
      else wr_ptr <= 2'h0;
    end
    else if (write) begin
      wr_ptr <= wr_ptr + 2'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    rd_ptr <= 2'h0;
  end
  else if (flush) begin
    rd_ptr <= 2'h0;
  end
  else if (clk_en) begin
    if (parallel_load | parallel_read) begin
      rd_ptr <= 2'h0;
    end
    else if (read) begin
      rd_ptr <= rd_ptr + 2'h1;
    end
  end
end
assign parallel_out = reg_array;
assign write = push & (~passthru) & ((~full) | pop | parallel_read);
always_comb begin
  if (passthru) begin
    data_out = data_in;
  end
  else data_out = reg_array[rd_ptr];
end
always_comb begin
  valid = pop & ((~empty) | passthru);
end
endmodule   // reg_fifo_d_4_w_1

module reg_fifo_d_4_w_1_unq0 #(
  parameter data_width = 16'h10
)
(
  input logic clk,
  input logic clk_en,
  input logic [0:0] [data_width-1:0] data_in,
  input logic flush,
  input logic [2:0] num_load,
  input logic [3:0][0:0] [data_width-1:0] parallel_in,
  input logic parallel_load,
  input logic parallel_read,
  input logic pop,
  input logic push,
  input logic rst_n,
  output logic [0:0] [data_width-1:0] data_out,
  output logic empty,
  output logic full,
  output logic [3:0][0:0] [data_width-1:0] parallel_out,
  output logic valid
);

logic [2:0] num_items;
logic passthru;
logic [1:0] rd_ptr;
logic read;
logic [3:0][0:0][data_width-1:0] reg_array;
logic [1:0] wr_ptr;
logic write;
assign full = num_items == 3'h4;
assign empty = num_items == 3'h0;
assign read = pop & (~passthru) & (~empty);
assign passthru = pop & push & empty;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_items <= 3'h0;
  end
  else if (flush) begin
    num_items <= 3'h0;
  end
  else if (clk_en) begin
    if (parallel_load) begin
      if (num_load == 3'h0) begin
        num_items <= 3'(push);
      end
      else num_items <= num_load;
    end
    else if (parallel_read) begin
      if (push) begin
        num_items <= 3'h1;
      end
      else num_items <= 3'h0;
    end
    else if (write & (~read)) begin
      num_items <= num_items + 3'h1;
    end
    else if ((~write) & read) begin
      num_items <= num_items - 3'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    reg_array <= 64'h0;
  end
  else if (flush) begin
    reg_array <= 64'h0;
  end
  else if (clk_en) begin
    if (parallel_load) begin
      reg_array <= parallel_in;
    end
    else if (write) begin
      if (parallel_read) begin
        reg_array[0] <= data_in;
      end
      else reg_array[wr_ptr] <= data_in;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    wr_ptr <= 2'h0;
  end
  else if (flush) begin
    wr_ptr <= 2'h0;
  end
  else if (clk_en) begin
    if (parallel_load) begin
      wr_ptr <= num_load[1:0];
    end
    else if (parallel_read) begin
      if (push) begin
        wr_ptr <= 2'h1;
      end
      else wr_ptr <= 2'h0;
    end
    else if (write) begin
      wr_ptr <= wr_ptr + 2'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    rd_ptr <= 2'h0;
  end
  else if (flush) begin
    rd_ptr <= 2'h0;
  end
  else if (clk_en) begin
    if (parallel_load | parallel_read) begin
      rd_ptr <= 2'h0;
    end
    else if (read) begin
      rd_ptr <= rd_ptr + 2'h1;
    end
  end
end
assign parallel_out = reg_array;
assign write = push & (~passthru) & ((~full) | pop | parallel_read);
always_comb begin
  if (passthru) begin
    data_out = data_in;
  end
  else data_out = reg_array[rd_ptr];
end
always_comb begin
  valid = pop & ((~empty) | passthru);
end
endmodule   // reg_fifo_d_4_w_1_unq0

module sched_gen_6_16 (
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic enable,
  input logic finished,
  input logic flush,
  input logic [2:0] mux_sel,
  input logic rst_n,
  input logic [15:0] sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] sched_addr_gen_strides,
  output logic valid_output
);

logic [15:0] addr_out;
logic valid_gate;
logic valid_gate_inv;
logic valid_out;
assign valid_gate = ~valid_gate_inv;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    valid_gate_inv <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      valid_gate_inv <= 1'h0;
    end
    else if (finished) begin
      valid_gate_inv <= 1'h1;
    end
  end
end
always_comb begin
  valid_out = (cycle_count == addr_out) & valid_gate & enable;
end
always_comb begin
  valid_output = valid_out;
end
addr_gen_6_16 sched_addr_gen (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(mux_sel),
  .restart(1'h0),
  .rst_n(rst_n),
  .starting_addr(sched_addr_gen_starting_addr),
  .step(valid_out),
  .strides(sched_addr_gen_strides),
  .addr_out(addr_out)
);

endmodule   // sched_gen_6_16

module sram_sp__0 (
  input logic clk,
  input logic clk_en,
  input logic [63:0] data_in_p0,
  input logic flush,
  input logic [8:0] read_addr_p0,
  input logic read_enable_p0,
  input logic [8:0] write_addr_p0,
  input logic write_enable_p0,
  output logic [63:0] data_out_p0
);

logic [8:0] mem_stub_A;
logic mem_stub_CEN;
logic mem_stub_RDWEN;
assign mem_stub_A = write_enable_p0 ? write_addr_p0: read_addr_p0;
assign mem_stub_RDWEN = ~write_enable_p0;
assign mem_stub_CEN = ~(write_enable_p0 | read_enable_p0);
IN12LP_S1DB_W00512B032M04S2_H_2_wide_1_deep mem_stub (
  .A(mem_stub_A),
  .CEN(mem_stub_CEN),
  .CLK(clk),
  .D(data_in_p0),
  .MA_SAWL0(1'h0),
  .MA_SAWL1(1'h0),
  .MA_STABAS0(1'h0),
  .MA_STABAS1(1'h0),
  .MA_VD0(1'h0),
  .MA_VD1(1'h0),
  .MA_WL0(1'h0),
  .MA_WL1(1'h0),
  .MA_WRAS0(1'h0),
  .MA_WRAS1(1'h0),
  .MA_WRT(1'h0),
  .RDWEN(mem_stub_RDWEN),
  .T_LOGIC(1'h0),
  .T_Q_RST(1'h0),
  .clk_en(clk_en),
  .flush(flush),
  .Q(data_out_p0)
);

endmodule   // sram_sp__0

module stencil_valid (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [3:0] loops_stencil_valid_dimensionality,
  input logic [5:0] [15:0] loops_stencil_valid_ranges,
  input logic rst_n,
  input logic stencil_valid_sched_gen_enable,
  input logic [15:0] stencil_valid_sched_gen_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] stencil_valid_sched_gen_sched_addr_gen_strides,
  output logic stencil_valid
);

logic [15:0] cycle_count;
logic flushed;
logic [2:0] loops_stencil_valid_mux_sel_out;
logic loops_stencil_valid_restart;
logic stencil_valid_internal;
assign stencil_valid = stencil_valid_internal & flushed;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    cycle_count <= 16'h0;
  end
  else if (clk_en) begin
    if (flushed) begin
      cycle_count <= cycle_count + 16'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    flushed <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      flushed <= 1'h1;
    end
  end
end
for_loop_6_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(4'h6))
loops_stencil_valid (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_stencil_valid_dimensionality),
  .flush(flush),
  .ranges(loops_stencil_valid_ranges),
  .rst_n(rst_n),
  .step(stencil_valid_internal),
  .mux_sel_out(loops_stencil_valid_mux_sel_out),
  .restart(loops_stencil_valid_restart)
);

sched_gen_6_16 stencil_valid_sched_gen (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(stencil_valid_sched_gen_enable),
  .finished(loops_stencil_valid_restart),
  .flush(flush),
  .mux_sel(loops_stencil_valid_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(stencil_valid_sched_gen_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(stencil_valid_sched_gen_sched_addr_gen_strides),
  .valid_output(stencil_valid_internal)
);

endmodule   // stencil_valid

module stencil_valid_flat (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic rst_n,
  input logic [3:0] stencil_valid_inst_loops_stencil_valid_dimensionality,
  input logic [5:0] [15:0] stencil_valid_inst_loops_stencil_valid_ranges,
  input logic stencil_valid_inst_stencil_valid_sched_gen_enable,
  input logic [15:0] stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides,
  output logic stencil_valid_f_
);

stencil_valid stencil_valid_inst (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .loops_stencil_valid_dimensionality(stencil_valid_inst_loops_stencil_valid_dimensionality),
  .loops_stencil_valid_ranges(stencil_valid_inst_loops_stencil_valid_ranges),
  .rst_n(rst_n),
  .stencil_valid_sched_gen_enable(stencil_valid_inst_stencil_valid_sched_gen_enable),
  .stencil_valid_sched_gen_sched_addr_gen_starting_addr(stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr),
  .stencil_valid_sched_gen_sched_addr_gen_strides(stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides),
  .stencil_valid(stencil_valid_f_)
);

endmodule   // stencil_valid_flat

module storage_config_seq_unq0 (
  input logic clk,
  input logic clk_en,
  input logic [7:0] config_addr_in,
  input logic [15:0] config_data_in,
  input logic [1:0] config_en,
  input logic config_rd,
  input logic config_wr,
  input logic flush,
  input logic [0:0][3:0] [15:0] rd_data_stg,
  input logic rst_n,
  output logic [8:0] addr_out,
  output logic [1:0] [15:0] rd_data_out,
  output logic ren_out,
  output logic wen_out,
  output logic [3:0] [15:0] wr_data
);

logic [1:0] cnt;
logic [2:0][15:0] data_wr_reg;
logic [1:0] rd_cnt;
logic [1:0] reduce_en;
logic set_to_addr;
assign reduce_en[0] = |config_en[0];
assign reduce_en[1] = |config_en[1];
always_comb begin
  set_to_addr = 1'h0;
  for (int unsigned i = 0; i < 2; i += 1) begin
      if (reduce_en[1'(i)]) begin
        set_to_addr = 1'(i);
      end
    end
end
assign addr_out = {set_to_addr, config_addr_in};

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    cnt <= 2'h0;
  end
  else if (flush) begin
    cnt <= 2'h0;
  end
  else if ((config_wr | config_rd) & (|config_en)) begin
    cnt <= cnt + 2'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    rd_cnt <= 2'h0;
  end
  else if (flush) begin
    rd_cnt <= 2'h0;
  end
  else rd_cnt <= cnt;
end
assign rd_data_out[0] = rd_data_stg[0][rd_cnt];
assign rd_data_out[1] = rd_data_stg[0][rd_cnt];

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    data_wr_reg <= 48'h0;
  end
  else if (flush) begin
    data_wr_reg <= 48'h0;
  end
  else if (config_wr & (cnt < 2'h3)) begin
    data_wr_reg[cnt] <= config_data_in;
  end
end
assign wr_data[0] = data_wr_reg[0];
assign wr_data[1] = data_wr_reg[1];
assign wr_data[2] = data_wr_reg[2];
assign wr_data[3] = config_data_in;
assign wen_out = config_wr & (cnt == 2'h3);
assign ren_out = config_rd;
endmodule   // storage_config_seq_unq0

module strg_fifo (
  input logic clk,
  input logic clk_en,
  input logic [0:0][3:0] [15:0] data_from_strg,
  input logic [15:0] data_in,
  input logic [15:0] fifo_depth,
  input logic flush,
  input logic pop,
  input logic push,
  input logic rst_n,
  output logic [0:0] [8:0] addr_out,
  output logic [15:0] data_out,
  output logic [0:0][3:0] [15:0] data_to_strg,
  output logic empty,
  output logic full,
  output logic ren_to_strg,
  output logic valid_out,
  output logic wen_to_strg
);

logic [15:0] back_data_in;
logic [15:0] back_data_out;
logic back_empty;
logic back_full;
logic [2:0] back_num_load;
logic [2:0] back_occ;
logic [3:0][0:0][15:0] back_par_in;
logic back_pl;
logic back_pop;
logic back_push;
logic [0:0][15:0] back_rf_data_in;
logic [0:0][15:0] back_rf_data_out;
logic back_rf_parallel_load;
logic back_valid;
logic curr_bank_rd;
logic curr_bank_wr;
logic [3:0][15:0] front_combined;
logic [15:0] front_data_out;
logic front_empty;
logic front_full;
logic [2:0] front_occ;
logic [3:0][0:0][15:0] front_par_out;
logic front_par_read;
logic front_pop;
logic front_push;
logic [1:0] front_rd_ptr;
logic [0:0][15:0] front_rf_data_in;
logic [0:0][15:0] front_rf_data_out;
logic front_valid;
logic fw_is_1;
logic [15:0] num_items;
logic [15:0] num_words_mem;
logic prev_bank_rd;
logic queued_write;
logic [0:0][8:0] ren_addr;
logic ren_delay;
logic [0:0][8:0] wen_addr;
logic [0:0][3:0][15:0] write_queue;
assign curr_bank_wr = 1'h0;
assign curr_bank_rd = 1'h0;
assign front_push = push & ((~full) | pop);
assign front_rf_data_in[0] = data_in;
assign front_data_out = front_rf_data_out[0];
assign fw_is_1 = 1'h0;
assign back_pop = pop & ((~empty) | push);
assign back_rf_parallel_load = back_pl & (|back_num_load);
assign back_rf_data_in[0] = back_data_in;
assign back_data_out = back_rf_data_out[0];
always_comb begin
  wen_to_strg = ((~ren_to_strg) | 1'h0) & (queued_write | ((front_occ == 3'h4) & push &
      (~front_pop) & (curr_bank_wr == 1'h0)));
end
always_comb begin
  ren_to_strg = ((back_occ == 3'h1) | fw_is_1) & (curr_bank_rd == 1'h0) & (pop | ((back_occ ==
      3'h0) & (back_num_load == 3'h0))) & ((num_words_mem > 16'h1) | ((num_words_mem
      == 16'h1) & (~back_pl)));
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    ren_delay <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      ren_delay <= 1'h0;
    end
    else ren_delay <= |ren_to_strg;
  end
end
assign back_pl = ren_delay;
assign front_combined[0] = front_par_out[front_rd_ptr + 2'h0];
assign front_combined[1] = front_par_out[front_rd_ptr + 2'h1];
assign front_combined[2] = front_par_out[front_rd_ptr + 2'h2];
assign front_combined[3] = front_par_out[front_rd_ptr + 2'h3];
assign data_to_strg[0] = queued_write ? write_queue[0]: front_combined;
assign back_data_in = front_data_out;
assign back_push = front_valid;
always_comb begin
  front_pop = ((num_words_mem == 16'h0) | ((num_words_mem == 16'h1) & back_pl)) & ((~back_pl)
      | (back_pl & (back_num_load == 3'h0))) & ((~(back_occ == 3'h4)) | pop) &
      ((~(front_occ == 3'h0)) | push);
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    write_queue[0] <= 64'h0;
    queued_write <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      write_queue[0] <= 64'h0;
      queued_write <= 1'h0;
    end
    else if (front_par_read & (~wen_to_strg) & (curr_bank_wr == 1'h0)) begin
      write_queue[0] <= front_combined;
      queued_write <= 1'h1;
    end
    else if (wen_to_strg) begin
      queued_write <= 1'h0;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_words_mem <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      num_words_mem <= 16'h0;
    end
    else if ((~back_pl) & front_par_read) begin
      num_words_mem <= num_words_mem + 16'h1;
    end
    else if (back_pl & (~front_par_read)) begin
      num_words_mem <= num_words_mem - 16'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    front_occ <= 3'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      front_occ <= 3'h0;
    end
    else if (front_par_read) begin
      if (front_push) begin
        front_occ <= 3'h1;
      end
      else front_occ <= 3'h0;
    end
    else if (front_push & (~front_pop)) begin
      front_occ <= front_occ + 3'h1;
    end
    else if ((~front_push) & front_pop) begin
      front_occ <= front_occ - 3'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    back_occ <= 3'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      back_occ <= 3'h0;
    end
    else if (back_pl) begin
      if (back_num_load == 3'h0) begin
        back_occ <= 3'(back_push);
      end
      else back_occ <= back_num_load;
    end
    else if (back_push & (~back_pop)) begin
      back_occ <= back_occ + 3'h1;
    end
    else if ((~back_push) & back_pop) begin
      back_occ <= back_occ - 3'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    prev_bank_rd <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      prev_bank_rd <= 1'h0;
    end
    else prev_bank_rd <= curr_bank_rd;
  end
end
assign back_par_in[0] = (back_num_load == 3'h4) ? data_from_strg[prev_bank_rd][0]:
    data_from_strg[prev_bank_rd][1];
assign back_par_in[1] = (back_num_load == 3'h4) ? data_from_strg[prev_bank_rd][1]:
    data_from_strg[prev_bank_rd][2];
assign back_par_in[2] = (back_num_load == 3'h4) ? data_from_strg[prev_bank_rd][2]:
    data_from_strg[prev_bank_rd][3];
assign back_par_in[3] = (back_num_load == 3'h4) ? data_from_strg[prev_bank_rd][3]: 16'h0;
always_comb begin
  front_par_read = (front_occ == 3'h4) & push & (~front_pop);
end
always_comb begin
  if (back_pl) begin
    back_num_load = pop ? 3'h3: 3'h4;
  end
  else back_num_load = 3'h0;
end
assign data_out = back_pl ? data_from_strg[prev_bank_rd][0]: back_data_out;
assign valid_out = back_pl ? pop: back_valid;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    wen_addr[0] <= 9'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      wen_addr[0] <= 9'h0;
    end
    else if (wen_to_strg) begin
      wen_addr[0] <= wen_addr[0] + 9'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    ren_addr[0] <= 9'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      ren_addr[0] <= 9'h0;
    end
    else if (ren_to_strg) begin
      ren_addr[0] <= ren_addr[0] + 9'h1;
    end
  end
end
assign addr_out[0] = wen_to_strg ? wen_addr[0]: ren_addr[0];
always_comb begin
  num_items = 16'(num_words_mem * 16'h4) + 16'(front_occ) + 16'(back_occ);
end
assign empty = num_items == 16'h0;
assign full = fifo_depth == num_items;
reg_fifo_d_4_w_1 #(
  .data_width(16'h10))
front_rf (
  .clk(clk),
  .clk_en(clk_en),
  .data_in(front_rf_data_in),
  .flush(flush),
  .num_load(3'h0),
  .parallel_in(64'h0),
  .parallel_load(1'h0),
  .parallel_read(front_par_read),
  .pop(front_pop),
  .push(front_push),
  .rst_n(rst_n),
  .data_out(front_rf_data_out),
  .empty(front_empty),
  .full(front_full),
  .parallel_out(front_par_out),
  .rd_ptr_out(front_rd_ptr),
  .valid(front_valid)
);

reg_fifo_d_4_w_1_unq0 #(
  .data_width(16'h10))
back_rf (
  .clk(clk),
  .clk_en(clk_en),
  .data_in(back_rf_data_in),
  .flush(flush),
  .num_load(back_num_load),
  .parallel_in(back_par_in),
  .parallel_load(back_rf_parallel_load),
  .parallel_read(1'h0),
  .pop(back_pop),
  .push(back_push),
  .rst_n(rst_n),
  .data_out(back_rf_data_out),
  .empty(back_empty),
  .full(back_full),
  .valid(back_valid)
);

endmodule   // strg_fifo

module strg_fifo_flat (
  input logic clk,
  input logic clk_en,
  input logic [0:0][3:0] [15:0] data_from_strg_lifted,
  input logic [0:0] [15:0] data_in_f_,
  input logic flush,
  input logic pop_f_,
  input logic push_f_,
  input logic rst_n,
  input logic [15:0] strg_fifo_inst_fifo_depth,
  output logic [0:0] [8:0] addr_out_lifted,
  output logic [0:0] [15:0] data_out_f_,
  output logic [0:0][3:0] [15:0] data_to_strg_lifted,
  output logic empty_f_,
  output logic full_f_,
  output logic ren_to_strg_lifted,
  output logic valid_out_f_,
  output logic wen_to_strg_lifted
);

logic [0:0][15:0] data_in_f__intercept;
logic [0:0][15:0] data_out_f__intercept;
logic [15:0] strg_fifo_inst_data_out;
assign data_in_f__intercept = data_in_f_;
assign data_out_f__intercept[0] = strg_fifo_inst_data_out;
assign data_out_f_ = data_out_f__intercept;
strg_fifo strg_fifo_inst (
  .clk(clk),
  .clk_en(clk_en),
  .data_from_strg(data_from_strg_lifted),
  .data_in(data_in_f__intercept[0]),
  .fifo_depth(strg_fifo_inst_fifo_depth),
  .flush(flush),
  .pop(pop_f_),
  .push(push_f_),
  .rst_n(rst_n),
  .addr_out(addr_out_lifted),
  .data_out(strg_fifo_inst_data_out),
  .data_to_strg(data_to_strg_lifted),
  .empty(empty_f_),
  .full(full_f_),
  .ren_to_strg(ren_to_strg_lifted),
  .valid_out(valid_out_f_),
  .wen_to_strg(wen_to_strg_lifted)
);

endmodule   // strg_fifo_flat

module strg_ram (
  input logic clk,
  input logic clk_en,
  input logic [0:0][3:0] [15:0] data_from_strg,
  input logic [15:0] data_in,
  input logic flush,
  input logic [15:0] rd_addr_in,
  input logic ren,
  input logic rst_n,
  input logic wen,
  input logic [15:0] wr_addr_in,
  output logic [0:0] [8:0] addr_out,
  output logic [15:0] data_out,
  output logic [0:0][3:0] [15:0] data_to_strg,
  output logic ready,
  output logic ren_to_strg,
  output logic valid_out,
  output logic wen_to_strg
);

typedef enum logic[1:0] {
  IDLE = 2'h0,
  MODIFY = 2'h1,
  READ = 2'h2,
  _DEFAULT = 2'h3
} r_w_seq_state;
logic [15:0] addr_to_write;
logic [3:0][15:0] data_combined;
logic [15:0] data_to_write;
r_w_seq_state r_w_seq_current_state;
r_w_seq_state r_w_seq_next_state;
logic [15:0] rd_addr;
logic rd_bank;
logic rd_valid;
logic read_gate;
logic [15:0] wr_addr;
logic write_gate;
assign wr_addr = wr_addr_in;
assign rd_addr = wr_addr_in;
assign rd_bank = 1'h0;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    rd_valid <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      rd_valid <= 1'h0;
    end
    else rd_valid <= ren & (~wen);
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    data_to_write <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      data_to_write <= 16'h0;
    end
    else data_to_write <= data_in;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    addr_to_write <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      addr_to_write <= 16'h0;
    end
    else addr_to_write <= wr_addr;
  end
end
assign data_to_strg[0] = data_combined;
assign ren_to_strg = (wen | ren) & read_gate;
assign wen_to_strg = write_gate;
always_comb begin
  addr_out[0] = rd_addr[10:2];
  if (wen & (~write_gate)) begin
    addr_out[0] = wr_addr[10:2];
  end
  else if (write_gate) begin
    addr_out[0] = addr_to_write[10:2];
  end
end
always_comb begin
  if (addr_to_write[1:0] == 2'h0) begin
    data_combined[0] = data_to_write;
  end
  else data_combined[0] = data_from_strg[rd_bank][0];
end
always_comb begin
  if (addr_to_write[1:0] == 2'h1) begin
    data_combined[1] = data_to_write;
  end
  else data_combined[1] = data_from_strg[rd_bank][1];
end
always_comb begin
  if (addr_to_write[1:0] == 2'h2) begin
    data_combined[2] = data_to_write;
  end
  else data_combined[2] = data_from_strg[rd_bank][2];
end
always_comb begin
  if (addr_to_write[1:0] == 2'h3) begin
    data_combined[3] = data_to_write;
  end
  else data_combined[3] = data_from_strg[rd_bank][3];
end

always_ff @(posedge clk, negedge rst_n) begin
  if (!rst_n) begin
    r_w_seq_current_state <= IDLE;
  end
  else r_w_seq_current_state <= r_w_seq_next_state;
end
always_comb begin
  r_w_seq_next_state = r_w_seq_current_state;
  unique case (r_w_seq_current_state)
    IDLE: begin
        if ((~wen) & (~ren)) begin
          r_w_seq_next_state = IDLE;
        end
        else if (wen) begin
          r_w_seq_next_state = MODIFY;
        end
        else if (ren & (~wen)) begin
          r_w_seq_next_state = READ;
        end
      end
    MODIFY: begin
        if (1'h1) begin
          r_w_seq_next_state = IDLE;
        end
      end
    READ: begin
        if ((~wen) & (~ren)) begin
          r_w_seq_next_state = IDLE;
        end
        else if (wen) begin
          r_w_seq_next_state = MODIFY;
        end
        else if (ren & (~wen)) begin
          r_w_seq_next_state = READ;
        end
      end
    _DEFAULT: begin
        if (1'h1) begin
          r_w_seq_next_state = _DEFAULT;
        end
      end
  endcase
end
always_comb begin
  unique case (r_w_seq_current_state)
    IDLE: begin :r_w_seq_IDLE_Output
        data_out = 16'h0;
        read_gate = 1'h1;
        ready = 1'h1;
        valid_out = 1'h0;
        write_gate = 1'h0;
      end :r_w_seq_IDLE_Output
    MODIFY: begin :r_w_seq_MODIFY_Output
        data_out = 16'h0;
        read_gate = 1'h0;
        ready = 1'h0;
        valid_out = 1'h0;
        write_gate = 1'h1;
      end :r_w_seq_MODIFY_Output
    READ: begin :r_w_seq_READ_Output
        data_out = data_from_strg[rd_bank][addr_to_write[1:0]];
        read_gate = 1'h1;
        ready = 1'h1;
        valid_out = 1'h1;
        write_gate = 1'h0;
      end :r_w_seq_READ_Output
    _DEFAULT: begin :r_w_seq__DEFAULT_Output
        data_out = 16'h0;
        read_gate = 1'h0;
        ready = 1'h0;
        valid_out = 1'h0;
        write_gate = 1'h0;
      end :r_w_seq__DEFAULT_Output
  endcase
end
endmodule   // strg_ram

module strg_ram_flat (
  input logic clk,
  input logic clk_en,
  input logic [0:0][3:0] [15:0] data_from_strg_lifted,
  input logic [0:0] [15:0] data_in_f_,
  input logic flush,
  input logic [0:0] [15:0] rd_addr_in_f_,
  input logic ren_f_,
  input logic rst_n,
  input logic wen_f_,
  input logic [0:0] [15:0] wr_addr_in_f_,
  output logic [0:0] [8:0] addr_out_lifted,
  output logic [0:0] [15:0] data_out_f_,
  output logic [0:0][3:0] [15:0] data_to_strg_lifted,
  output logic ready_f_,
  output logic ren_to_strg_lifted,
  output logic valid_out_f_,
  output logic wen_to_strg_lifted
);

logic [0:0][15:0] data_in_f__intercept;
logic [0:0][15:0] data_out_f__intercept;
logic [0:0][15:0] rd_addr_in_f__intercept;
logic [15:0] strg_ram_inst_data_out;
logic [0:0][15:0] wr_addr_in_f__intercept;
assign rd_addr_in_f__intercept = rd_addr_in_f_;
assign wr_addr_in_f__intercept = wr_addr_in_f_;
assign data_in_f__intercept = data_in_f_;
assign data_out_f__intercept[0] = strg_ram_inst_data_out;
assign data_out_f_ = data_out_f__intercept;
strg_ram strg_ram_inst (
  .clk(clk),
  .clk_en(clk_en),
  .data_from_strg(data_from_strg_lifted),
  .data_in(data_in_f__intercept[0]),
  .flush(flush),
  .rd_addr_in(rd_addr_in_f__intercept[0]),
  .ren(ren_f_),
  .rst_n(rst_n),
  .wen(wen_f_),
  .wr_addr_in(wr_addr_in_f__intercept[0]),
  .addr_out(addr_out_lifted),
  .data_out(strg_ram_inst_data_out),
  .data_to_strg(data_to_strg_lifted),
  .ready(ready_f_),
  .ren_to_strg(ren_to_strg_lifted),
  .valid_out(valid_out_f_),
  .wen_to_strg(wen_to_strg_lifted)
);

endmodule   // strg_ram_flat

module strg_ub_agg_only (
  input logic [1:0] agg_read,
  input logic [3:0] agg_read_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] agg_read_addr_gen_0_strides,
  input logic [3:0] agg_read_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] agg_read_addr_gen_1_strides,
  input logic [3:0] agg_write_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] agg_write_addr_gen_0_strides,
  input logic [3:0] agg_write_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] agg_write_addr_gen_1_strides,
  input logic agg_write_sched_gen_0_enable,
  input logic [15:0] agg_write_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] agg_write_sched_gen_0_sched_addr_gen_strides,
  input logic agg_write_sched_gen_1_enable,
  input logic [15:0] agg_write_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] agg_write_sched_gen_1_sched_addr_gen_strides,
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic [1:0] [15:0] data_in,
  input logic [1:0] [2:0] floop_mux_sel,
  input logic [1:0] floop_restart,
  input logic flush,
  input logic [3:0] loops_in2buf_0_dimensionality,
  input logic [5:0] [15:0] loops_in2buf_0_ranges,
  input logic [3:0] loops_in2buf_1_dimensionality,
  input logic [5:0] [15:0] loops_in2buf_1_ranges,
  input logic rst_n,
  output logic [1:0][3:0] [15:0] agg_data_out
);

logic [1:0][3:0][3:0][15:0] agg;
logic [1:0][1:0] agg_read_addr;
logic [3:0] agg_read_addr_gen_0_addr_out;
logic [3:0] agg_read_addr_gen_1_addr_out;
logic [1:0][7:0] agg_read_addr_gen_out;
logic [1:0] agg_write;
logic [1:0][3:0] agg_write_addr;
logic [3:0] agg_write_addr_gen_0_addr_out;
logic [3:0] agg_write_addr_gen_1_addr_out;
logic agg_write_sched_gen_0_valid_output;
logic agg_write_sched_gen_1_valid_output;
logic [2:0] loops_in2buf_0_mux_sel_out;
logic loops_in2buf_0_restart;
logic [2:0] loops_in2buf_1_mux_sel_out;
logic loops_in2buf_1_restart;
assign agg_write_addr[0] = agg_write_addr_gen_0_addr_out;
assign agg_write[0] = agg_write_sched_gen_0_valid_output;

always_ff @(posedge clk) begin
  if (clk_en) begin
    if (agg_write[0]) begin
      agg[0][agg_write_addr[0][3:2]][agg_write_addr[0][1:0]] <= data_in[0];
    end
  end
end
assign agg_read_addr_gen_out[0][3:0] = agg_read_addr_gen_0_addr_out;
assign agg_read_addr_gen_out[0][7:4] = 4'h0;
assign agg_read_addr[0] = agg_read_addr_gen_out[0][1:0];
always_comb begin
  agg_data_out[0] = agg[0][agg_read_addr[0]];
end
assign agg_write_addr[1] = agg_write_addr_gen_1_addr_out;
assign agg_write[1] = agg_write_sched_gen_1_valid_output;

always_ff @(posedge clk) begin
  if (clk_en) begin
    if (agg_write[1]) begin
      agg[1][agg_write_addr[1][3:2]][agg_write_addr[1][1:0]] <= data_in[1];
    end
  end
end
assign agg_read_addr_gen_out[1][3:0] = agg_read_addr_gen_1_addr_out;
assign agg_read_addr_gen_out[1][7:4] = 4'h0;
assign agg_read_addr[1] = agg_read_addr_gen_out[1][1:0];
always_comb begin
  agg_data_out[1] = agg[1][agg_read_addr[1]];
end
for_loop_6_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(4'h6))
loops_in2buf_0 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_in2buf_0_dimensionality),
  .flush(flush),
  .ranges(loops_in2buf_0_ranges),
  .rst_n(rst_n),
  .step(agg_write[0]),
  .mux_sel_out(loops_in2buf_0_mux_sel_out),
  .restart(loops_in2buf_0_restart)
);

addr_gen_6_4 agg_write_addr_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(loops_in2buf_0_mux_sel_out),
  .restart(loops_in2buf_0_restart),
  .rst_n(rst_n),
  .starting_addr(agg_write_addr_gen_0_starting_addr),
  .step(agg_write[0]),
  .strides(agg_write_addr_gen_0_strides),
  .addr_out(agg_write_addr_gen_0_addr_out)
);

sched_gen_6_16 agg_write_sched_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(agg_write_sched_gen_0_enable),
  .finished(loops_in2buf_0_restart),
  .flush(flush),
  .mux_sel(loops_in2buf_0_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(agg_write_sched_gen_0_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(agg_write_sched_gen_0_sched_addr_gen_strides),
  .valid_output(agg_write_sched_gen_0_valid_output)
);

addr_gen_6_4 agg_read_addr_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(floop_mux_sel[0]),
  .restart(floop_restart[0]),
  .rst_n(rst_n),
  .starting_addr(agg_read_addr_gen_0_starting_addr),
  .step(agg_read[0]),
  .strides(agg_read_addr_gen_0_strides),
  .addr_out(agg_read_addr_gen_0_addr_out)
);

for_loop_6_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(4'h6))
loops_in2buf_1 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_in2buf_1_dimensionality),
  .flush(flush),
  .ranges(loops_in2buf_1_ranges),
  .rst_n(rst_n),
  .step(agg_write[1]),
  .mux_sel_out(loops_in2buf_1_mux_sel_out),
  .restart(loops_in2buf_1_restart)
);

addr_gen_6_4 agg_write_addr_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(loops_in2buf_1_mux_sel_out),
  .restart(loops_in2buf_1_restart),
  .rst_n(rst_n),
  .starting_addr(agg_write_addr_gen_1_starting_addr),
  .step(agg_write[1]),
  .strides(agg_write_addr_gen_1_strides),
  .addr_out(agg_write_addr_gen_1_addr_out)
);

sched_gen_6_16 agg_write_sched_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(agg_write_sched_gen_1_enable),
  .finished(loops_in2buf_1_restart),
  .flush(flush),
  .mux_sel(loops_in2buf_1_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(agg_write_sched_gen_1_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(agg_write_sched_gen_1_sched_addr_gen_strides),
  .valid_output(agg_write_sched_gen_1_valid_output)
);

addr_gen_6_4 agg_read_addr_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(floop_mux_sel[1]),
  .restart(floop_restart[1]),
  .rst_n(rst_n),
  .starting_addr(agg_read_addr_gen_1_starting_addr),
  .step(agg_read[1]),
  .strides(agg_read_addr_gen_1_strides),
  .addr_out(agg_read_addr_gen_1_addr_out)
);

endmodule   // strg_ub_agg_only

module strg_ub_agg_sram_shared (
  input logic agg_read_sched_gen_0_enable,
  input logic [15:0] agg_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] agg_read_sched_gen_0_sched_addr_gen_strides,
  input logic agg_read_sched_gen_1_enable,
  input logic [15:0] agg_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] agg_read_sched_gen_1_sched_addr_gen_strides,
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic flush,
  input logic [3:0] loops_in2buf_autovec_write_0_dimensionality,
  input logic [5:0] [15:0] loops_in2buf_autovec_write_0_ranges,
  input logic [3:0] loops_in2buf_autovec_write_1_dimensionality,
  input logic [5:0] [15:0] loops_in2buf_autovec_write_1_ranges,
  input logic rst_n,
  output logic [1:0] agg_read_out,
  output logic [1:0] [2:0] floop_mux_sel,
  output logic [1:0] floop_restart
);

logic [1:0] agg_read;
logic agg_read_sched_gen_0_valid_output;
logic agg_read_sched_gen_1_valid_output;
logic [2:0] loops_in2buf_autovec_write_0_mux_sel_out;
logic loops_in2buf_autovec_write_0_restart;
logic [2:0] loops_in2buf_autovec_write_1_mux_sel_out;
logic loops_in2buf_autovec_write_1_restart;
assign agg_read_out = agg_read;
assign floop_mux_sel[0] = loops_in2buf_autovec_write_0_mux_sel_out;
assign floop_restart[0] = loops_in2buf_autovec_write_0_restart;
assign agg_read[0] = agg_read_sched_gen_0_valid_output;
assign floop_mux_sel[1] = loops_in2buf_autovec_write_1_mux_sel_out;
assign floop_restart[1] = loops_in2buf_autovec_write_1_restart;
assign agg_read[1] = agg_read_sched_gen_1_valid_output;
for_loop_6_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(4'h6))
loops_in2buf_autovec_write_0 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_in2buf_autovec_write_0_dimensionality),
  .flush(flush),
  .ranges(loops_in2buf_autovec_write_0_ranges),
  .rst_n(rst_n),
  .step(agg_read[0]),
  .mux_sel_out(loops_in2buf_autovec_write_0_mux_sel_out),
  .restart(loops_in2buf_autovec_write_0_restart)
);

sched_gen_6_16 agg_read_sched_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(agg_read_sched_gen_0_enable),
  .finished(loops_in2buf_autovec_write_0_restart),
  .flush(flush),
  .mux_sel(loops_in2buf_autovec_write_0_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(agg_read_sched_gen_0_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(agg_read_sched_gen_0_sched_addr_gen_strides),
  .valid_output(agg_read_sched_gen_0_valid_output)
);

for_loop_6_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(4'h6))
loops_in2buf_autovec_write_1 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_in2buf_autovec_write_1_dimensionality),
  .flush(flush),
  .ranges(loops_in2buf_autovec_write_1_ranges),
  .rst_n(rst_n),
  .step(agg_read[1]),
  .mux_sel_out(loops_in2buf_autovec_write_1_mux_sel_out),
  .restart(loops_in2buf_autovec_write_1_restart)
);

sched_gen_6_16 agg_read_sched_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(agg_read_sched_gen_1_enable),
  .finished(loops_in2buf_autovec_write_1_restart),
  .flush(flush),
  .mux_sel(loops_in2buf_autovec_write_1_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(agg_read_sched_gen_1_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(agg_read_sched_gen_1_sched_addr_gen_strides),
  .valid_output(agg_read_sched_gen_1_valid_output)
);

endmodule   // strg_ub_agg_sram_shared

module strg_ub_sram_only (
  input logic [1:0][3:0] [15:0] agg_data_out,
  input logic [1:0] agg_read,
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic [1:0] [2:0] floop_mux_sel,
  input logic [1:0] floop_restart,
  input logic flush,
  input logic [8:0] input_addr_gen_0_starting_addr,
  input logic [5:0] [8:0] input_addr_gen_0_strides,
  input logic [8:0] input_addr_gen_1_starting_addr,
  input logic [5:0] [8:0] input_addr_gen_1_strides,
  input logic [1:0] [2:0] loops_sram2tb_mux_sel,
  input logic [1:0] loops_sram2tb_restart,
  input logic [8:0] output_addr_gen_0_starting_addr,
  input logic [5:0] [8:0] output_addr_gen_0_strides,
  input logic [8:0] output_addr_gen_1_starting_addr,
  input logic [5:0] [8:0] output_addr_gen_1_strides,
  input logic rst_n,
  input logic [1:0] t_read,
  output logic [8:0] addr_to_sram,
  output logic cen_to_sram,
  output logic [3:0] [15:0] data_to_sram,
  output logic wen_to_sram
);

logic [8:0] addr;
logic [3:0][15:0] decode_ret_agg_read_agg_data_out;
logic [15:0] decode_ret_agg_read_s_write_addr;
logic [15:0] decode_ret_t_read_s_read_addr;
logic decode_sel_done_agg_read_agg_data_out;
logic decode_sel_done_agg_read_s_write_addr;
logic decode_sel_done_t_read_s_read_addr;
logic [8:0] input_addr_gen_0_addr_out;
logic [8:0] input_addr_gen_1_addr_out;
logic [8:0] output_addr_gen_0_addr_out;
logic [8:0] output_addr_gen_1_addr_out;
logic read;
logic [1:0][15:0] s_read_addr;
logic [1:0][15:0] s_write_addr;
logic [3:0][15:0] sram_write_data;
logic write;
assign s_write_addr[0][8:0] = input_addr_gen_0_addr_out;
assign s_write_addr[0][15:9] = 7'h0;
assign s_write_addr[1][8:0] = input_addr_gen_1_addr_out;
assign s_write_addr[1][15:9] = 7'h0;
assign s_read_addr[0][8:0] = output_addr_gen_0_addr_out;
assign s_read_addr[0][15:9] = 7'h0;
assign s_read_addr[1][8:0] = output_addr_gen_1_addr_out;
assign s_read_addr[1][15:9] = 7'h0;
assign data_to_sram = sram_write_data;
assign wen_to_sram = write;
always_comb begin
  decode_sel_done_agg_read_s_write_addr = 1'h0;
  decode_ret_agg_read_s_write_addr = 16'h0;
  for (int unsigned i = 0; i < 2; i += 1) begin
      if ((~decode_sel_done_agg_read_s_write_addr) & agg_read[1'(i)]) begin
        decode_ret_agg_read_s_write_addr = s_write_addr[1'(i)];
        decode_sel_done_agg_read_s_write_addr = 1'h1;
      end
    end
end
always_comb begin
  decode_sel_done_t_read_s_read_addr = 1'h0;
  decode_ret_t_read_s_read_addr = 16'h0;
  for (int unsigned i = 0; i < 2; i += 1) begin
      if ((~decode_sel_done_t_read_s_read_addr) & t_read[1'(i)]) begin
        decode_ret_t_read_s_read_addr = s_read_addr[1'(i)];
        decode_sel_done_t_read_s_read_addr = 1'h1;
      end
    end
end
assign cen_to_sram = write | read;
assign addr_to_sram = addr;
always_comb begin
  if (write) begin
    addr = decode_ret_agg_read_s_write_addr[8:0];
  end
  else addr = decode_ret_t_read_s_read_addr[8:0];
end
assign write = |agg_read;
assign read = |t_read;
always_comb begin
  decode_sel_done_agg_read_agg_data_out = 1'h0;
  decode_ret_agg_read_agg_data_out = 64'h0;
  for (int unsigned i = 0; i < 2; i += 1) begin
      if ((~decode_sel_done_agg_read_agg_data_out) & agg_read[1'(i)]) begin
        decode_ret_agg_read_agg_data_out = agg_data_out[1'(i)];
        decode_sel_done_agg_read_agg_data_out = 1'h1;
      end
    end
end
assign sram_write_data = decode_ret_agg_read_agg_data_out;
addr_gen_6_9 input_addr_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(floop_mux_sel[0]),
  .restart(floop_restart[0]),
  .rst_n(rst_n),
  .starting_addr(input_addr_gen_0_starting_addr),
  .step(agg_read[0]),
  .strides(input_addr_gen_0_strides),
  .addr_out(input_addr_gen_0_addr_out)
);

addr_gen_6_9 input_addr_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(floop_mux_sel[1]),
  .restart(floop_restart[1]),
  .rst_n(rst_n),
  .starting_addr(input_addr_gen_1_starting_addr),
  .step(agg_read[1]),
  .strides(input_addr_gen_1_strides),
  .addr_out(input_addr_gen_1_addr_out)
);

addr_gen_6_9 output_addr_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(loops_sram2tb_mux_sel[0]),
  .restart(loops_sram2tb_restart[0]),
  .rst_n(rst_n),
  .starting_addr(output_addr_gen_0_starting_addr),
  .step(t_read[0]),
  .strides(output_addr_gen_0_strides),
  .addr_out(output_addr_gen_0_addr_out)
);

addr_gen_6_9 output_addr_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(loops_sram2tb_mux_sel[1]),
  .restart(loops_sram2tb_restart[1]),
  .rst_n(rst_n),
  .starting_addr(output_addr_gen_1_starting_addr),
  .step(t_read[1]),
  .strides(output_addr_gen_1_strides),
  .addr_out(output_addr_gen_1_addr_out)
);

endmodule   // strg_ub_sram_only

module strg_ub_sram_tb_shared (
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic flush,
  input logic [3:0] loops_buf2out_autovec_read_0_dimensionality,
  input logic [5:0] [15:0] loops_buf2out_autovec_read_0_ranges,
  input logic [3:0] loops_buf2out_autovec_read_1_dimensionality,
  input logic [5:0] [15:0] loops_buf2out_autovec_read_1_ranges,
  input logic output_sched_gen_0_enable,
  input logic [15:0] output_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] output_sched_gen_0_sched_addr_gen_strides,
  input logic output_sched_gen_1_enable,
  input logic [15:0] output_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] output_sched_gen_1_sched_addr_gen_strides,
  input logic rst_n,
  output logic [1:0] [2:0] loops_sram2tb_mux_sel,
  output logic [1:0] loops_sram2tb_restart,
  output logic [1:0] t_read_out
);

logic [2:0] loops_buf2out_autovec_read_0_mux_sel_out;
logic loops_buf2out_autovec_read_0_restart;
logic [2:0] loops_buf2out_autovec_read_1_mux_sel_out;
logic loops_buf2out_autovec_read_1_restart;
logic output_sched_gen_0_valid_output;
logic output_sched_gen_1_valid_output;
logic [1:0] t_read;
assign t_read_out = t_read;
assign loops_sram2tb_mux_sel[0] = loops_buf2out_autovec_read_0_mux_sel_out;
assign loops_sram2tb_restart[0] = loops_buf2out_autovec_read_0_restart;
assign t_read[0] = output_sched_gen_0_valid_output;
assign loops_sram2tb_mux_sel[1] = loops_buf2out_autovec_read_1_mux_sel_out;
assign loops_sram2tb_restart[1] = loops_buf2out_autovec_read_1_restart;
assign t_read[1] = output_sched_gen_1_valid_output;
for_loop_6_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(4'h6))
loops_buf2out_autovec_read_0 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_buf2out_autovec_read_0_dimensionality),
  .flush(flush),
  .ranges(loops_buf2out_autovec_read_0_ranges),
  .rst_n(rst_n),
  .step(t_read[0]),
  .mux_sel_out(loops_buf2out_autovec_read_0_mux_sel_out),
  .restart(loops_buf2out_autovec_read_0_restart)
);

sched_gen_6_16 output_sched_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(output_sched_gen_0_enable),
  .finished(loops_buf2out_autovec_read_0_restart),
  .flush(flush),
  .mux_sel(loops_buf2out_autovec_read_0_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(output_sched_gen_0_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(output_sched_gen_0_sched_addr_gen_strides),
  .valid_output(output_sched_gen_0_valid_output)
);

for_loop_6_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(4'h6))
loops_buf2out_autovec_read_1 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_buf2out_autovec_read_1_dimensionality),
  .flush(flush),
  .ranges(loops_buf2out_autovec_read_1_ranges),
  .rst_n(rst_n),
  .step(t_read[1]),
  .mux_sel_out(loops_buf2out_autovec_read_1_mux_sel_out),
  .restart(loops_buf2out_autovec_read_1_restart)
);

sched_gen_6_16 output_sched_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(output_sched_gen_1_enable),
  .finished(loops_buf2out_autovec_read_1_restart),
  .flush(flush),
  .mux_sel(loops_buf2out_autovec_read_1_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(output_sched_gen_1_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(output_sched_gen_1_sched_addr_gen_strides),
  .valid_output(output_sched_gen_1_valid_output)
);

endmodule   // strg_ub_sram_tb_shared

module strg_ub_tb_only (
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic flush,
  input logic [3:0] loops_buf2out_read_0_dimensionality,
  input logic [5:0] [15:0] loops_buf2out_read_0_ranges,
  input logic [3:0] loops_buf2out_read_1_dimensionality,
  input logic [5:0] [15:0] loops_buf2out_read_1_ranges,
  input logic [1:0] [2:0] loops_sram2tb_mux_sel,
  input logic [1:0] loops_sram2tb_restart,
  input logic rst_n,
  input logic [3:0] [15:0] sram_read_data,
  input logic [1:0] t_read,
  input logic [3:0] tb_read_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] tb_read_addr_gen_0_strides,
  input logic [3:0] tb_read_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] tb_read_addr_gen_1_strides,
  input logic tb_read_sched_gen_0_enable,
  input logic [15:0] tb_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] tb_read_sched_gen_0_sched_addr_gen_strides,
  input logic tb_read_sched_gen_1_enable,
  input logic [15:0] tb_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] tb_read_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] tb_write_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] tb_write_addr_gen_0_strides,
  input logic [3:0] tb_write_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] tb_write_addr_gen_1_strides,
  output logic [1:0] accessor_output,
  output logic [1:0] [15:0] data_out
);

logic [2:0] loops_buf2out_read_0_mux_sel_out;
logic loops_buf2out_read_0_restart;
logic [2:0] loops_buf2out_read_1_mux_sel_out;
logic loops_buf2out_read_1_restart;
logic [1:0][2:0] mux_sel_d1;
logic [1:0] restart_d1;
logic [1:0] t_read_d1;
logic [1:0][1:0][3:0][15:0] tb;
logic [1:0] tb_read;
logic [1:0][2:0] tb_read_addr;
logic [3:0] tb_read_addr_gen_0_addr_out;
logic [3:0] tb_read_addr_gen_1_addr_out;
logic tb_read_sched_gen_0_valid_output;
logic tb_read_sched_gen_1_valid_output;
logic [1:0][2:0] tb_write_addr;
logic [3:0] tb_write_addr_gen_0_addr_out;
logic [3:0] tb_write_addr_gen_1_addr_out;
assign accessor_output = tb_read;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    t_read_d1[0] <= 1'h0;
    mux_sel_d1[0] <= 3'h0;
    restart_d1[0] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      t_read_d1[0] <= 1'h0;
      mux_sel_d1[0] <= 3'h0;
      restart_d1[0] <= 1'h0;
    end
    else begin
      t_read_d1[0] <= t_read[0];
      mux_sel_d1[0] <= loops_sram2tb_mux_sel[0];
      restart_d1[0] <= loops_sram2tb_restart[0];
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    t_read_d1[1] <= 1'h0;
    mux_sel_d1[1] <= 3'h0;
    restart_d1[1] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      t_read_d1[1] <= 1'h0;
      mux_sel_d1[1] <= 3'h0;
      restart_d1[1] <= 1'h0;
    end
    else begin
      t_read_d1[1] <= t_read[1];
      mux_sel_d1[1] <= loops_sram2tb_mux_sel[1];
      restart_d1[1] <= loops_sram2tb_restart[1];
    end
  end
end
assign tb_write_addr[0] = tb_write_addr_gen_0_addr_out[2:0];

always_ff @(posedge clk) begin
  if (clk_en) begin
    if (t_read_d1[0]) begin
      tb[0][tb_write_addr[0][0]] <= sram_read_data;
    end
  end
end
assign tb_read_addr[0] = tb_read_addr_gen_0_addr_out[2:0];
assign tb_read[0] = tb_read_sched_gen_0_valid_output;
always_comb begin
  data_out[0] = tb[0][tb_read_addr[0][2]][tb_read_addr[0][1:0]];
end
assign tb_write_addr[1] = tb_write_addr_gen_1_addr_out[2:0];

always_ff @(posedge clk) begin
  if (clk_en) begin
    if (t_read_d1[1]) begin
      tb[1][tb_write_addr[1][0]] <= sram_read_data;
    end
  end
end
assign tb_read_addr[1] = tb_read_addr_gen_1_addr_out[2:0];
assign tb_read[1] = tb_read_sched_gen_1_valid_output;
always_comb begin
  data_out[1] = tb[1][tb_read_addr[1][2]][tb_read_addr[1][1:0]];
end
addr_gen_6_4 tb_write_addr_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(mux_sel_d1[0]),
  .restart(restart_d1[0]),
  .rst_n(rst_n),
  .starting_addr(tb_write_addr_gen_0_starting_addr),
  .step(t_read_d1[0]),
  .strides(tb_write_addr_gen_0_strides),
  .addr_out(tb_write_addr_gen_0_addr_out)
);

for_loop_6_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(4'h6))
loops_buf2out_read_0 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_buf2out_read_0_dimensionality),
  .flush(flush),
  .ranges(loops_buf2out_read_0_ranges),
  .rst_n(rst_n),
  .step(tb_read[0]),
  .mux_sel_out(loops_buf2out_read_0_mux_sel_out),
  .restart(loops_buf2out_read_0_restart)
);

addr_gen_6_4 tb_read_addr_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(loops_buf2out_read_0_mux_sel_out),
  .restart(loops_buf2out_read_0_restart),
  .rst_n(rst_n),
  .starting_addr(tb_read_addr_gen_0_starting_addr),
  .step(tb_read[0]),
  .strides(tb_read_addr_gen_0_strides),
  .addr_out(tb_read_addr_gen_0_addr_out)
);

sched_gen_6_16 tb_read_sched_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(tb_read_sched_gen_0_enable),
  .finished(loops_buf2out_read_0_restart),
  .flush(flush),
  .mux_sel(loops_buf2out_read_0_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(tb_read_sched_gen_0_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(tb_read_sched_gen_0_sched_addr_gen_strides),
  .valid_output(tb_read_sched_gen_0_valid_output)
);

addr_gen_6_4 tb_write_addr_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(mux_sel_d1[1]),
  .restart(restart_d1[1]),
  .rst_n(rst_n),
  .starting_addr(tb_write_addr_gen_1_starting_addr),
  .step(t_read_d1[1]),
  .strides(tb_write_addr_gen_1_strides),
  .addr_out(tb_write_addr_gen_1_addr_out)
);

for_loop_6_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(4'h6))
loops_buf2out_read_1 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_buf2out_read_1_dimensionality),
  .flush(flush),
  .ranges(loops_buf2out_read_1_ranges),
  .rst_n(rst_n),
  .step(tb_read[1]),
  .mux_sel_out(loops_buf2out_read_1_mux_sel_out),
  .restart(loops_buf2out_read_1_restart)
);

addr_gen_6_4 tb_read_addr_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(loops_buf2out_read_1_mux_sel_out),
  .restart(loops_buf2out_read_1_restart),
  .rst_n(rst_n),
  .starting_addr(tb_read_addr_gen_1_starting_addr),
  .step(tb_read[1]),
  .strides(tb_read_addr_gen_1_strides),
  .addr_out(tb_read_addr_gen_1_addr_out)
);

sched_gen_6_16 tb_read_sched_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(tb_read_sched_gen_1_enable),
  .finished(loops_buf2out_read_1_restart),
  .flush(flush),
  .mux_sel(loops_buf2out_read_1_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(tb_read_sched_gen_1_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(tb_read_sched_gen_1_sched_addr_gen_strides),
  .valid_output(tb_read_sched_gen_1_valid_output)
);

endmodule   // strg_ub_tb_only

module strg_ub_vec (
  input logic [3:0] agg_only_agg_read_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] agg_only_agg_read_addr_gen_0_strides,
  input logic [3:0] agg_only_agg_read_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] agg_only_agg_read_addr_gen_1_strides,
  input logic [3:0] agg_only_agg_write_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] agg_only_agg_write_addr_gen_0_strides,
  input logic [3:0] agg_only_agg_write_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] agg_only_agg_write_addr_gen_1_strides,
  input logic agg_only_agg_write_sched_gen_0_enable,
  input logic [15:0] agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] agg_only_agg_write_sched_gen_0_sched_addr_gen_strides,
  input logic agg_only_agg_write_sched_gen_1_enable,
  input logic [15:0] agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] agg_only_agg_write_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] agg_only_loops_in2buf_0_dimensionality,
  input logic [5:0] [15:0] agg_only_loops_in2buf_0_ranges,
  input logic [3:0] agg_only_loops_in2buf_1_dimensionality,
  input logic [5:0] [15:0] agg_only_loops_in2buf_1_ranges,
  input logic agg_sram_shared_agg_read_sched_gen_0_enable,
  input logic [15:0] agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides,
  input logic agg_sram_shared_agg_read_sched_gen_1_enable,
  input logic [15:0] agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality,
  input logic [5:0] [15:0] agg_sram_shared_loops_in2buf_autovec_write_0_ranges,
  input logic [3:0] agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality,
  input logic [5:0] [15:0] agg_sram_shared_loops_in2buf_autovec_write_1_ranges,
  input logic chain_chain_en,
  input logic [1:0] [15:0] chain_data_in,
  input logic clk,
  input logic clk_en,
  input logic [3:0] [15:0] data_from_strg,
  input logic [1:0] [15:0] data_in,
  input logic flush,
  input logic rst_n,
  input logic [8:0] sram_only_input_addr_gen_0_starting_addr,
  input logic [5:0] [8:0] sram_only_input_addr_gen_0_strides,
  input logic [8:0] sram_only_input_addr_gen_1_starting_addr,
  input logic [5:0] [8:0] sram_only_input_addr_gen_1_strides,
  input logic [8:0] sram_only_output_addr_gen_0_starting_addr,
  input logic [5:0] [8:0] sram_only_output_addr_gen_0_strides,
  input logic [8:0] sram_only_output_addr_gen_1_starting_addr,
  input logic [5:0] [8:0] sram_only_output_addr_gen_1_strides,
  input logic [3:0] sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality,
  input logic [5:0] [15:0] sram_tb_shared_loops_buf2out_autovec_read_0_ranges,
  input logic [3:0] sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality,
  input logic [5:0] [15:0] sram_tb_shared_loops_buf2out_autovec_read_1_ranges,
  input logic sram_tb_shared_output_sched_gen_0_enable,
  input logic [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides,
  input logic sram_tb_shared_output_sched_gen_1_enable,
  input logic [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] tb_only_loops_buf2out_read_0_dimensionality,
  input logic [5:0] [15:0] tb_only_loops_buf2out_read_0_ranges,
  input logic [3:0] tb_only_loops_buf2out_read_1_dimensionality,
  input logic [5:0] [15:0] tb_only_loops_buf2out_read_1_ranges,
  input logic [3:0] tb_only_tb_read_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] tb_only_tb_read_addr_gen_0_strides,
  input logic [3:0] tb_only_tb_read_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] tb_only_tb_read_addr_gen_1_strides,
  input logic tb_only_tb_read_sched_gen_0_enable,
  input logic [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_strides,
  input logic tb_only_tb_read_sched_gen_1_enable,
  input logic [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] tb_only_tb_write_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] tb_only_tb_write_addr_gen_0_strides,
  input logic [3:0] tb_only_tb_write_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] tb_only_tb_write_addr_gen_1_strides,
  output logic [1:0] accessor_output,
  output logic [8:0] addr_out,
  output logic [1:0] [15:0] data_out,
  output logic [3:0] [15:0] data_to_strg,
  output logic ren_to_strg,
  output logic wen_to_strg
);

logic [1:0] accessor_output_int;
logic [1:0][3:0][15:0] agg_only_agg_data_out;
logic [1:0] agg_only_agg_read;
logic [1:0][2:0] agg_only_floop_mux_sel;
logic [1:0] agg_only_floop_restart;
logic [1:0] agg_sram_shared_agg_read_out;
logic [1:0][2:0] agg_sram_shared_floop_mux_sel;
logic [1:0] agg_sram_shared_floop_restart;
logic [15:0] cycle_count;
logic [1:0][15:0] data_out_int;
logic [1:0][2:0] sram_only_loops_sram2tb_mux_sel;
logic [1:0] sram_only_loops_sram2tb_restart;
logic [1:0] sram_only_t_read;
logic [1:0][2:0] sram_tb_shared_loops_sram2tb_mux_sel;
logic [1:0] sram_tb_shared_loops_sram2tb_restart;
logic [1:0] sram_tb_shared_t_read_out;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    cycle_count <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      cycle_count <= 16'h0;
    end
    else if (1'h1) begin
      cycle_count <= cycle_count + 16'h1;
    end
  end
end
assign agg_only_agg_read = agg_sram_shared_agg_read_out;
assign agg_only_floop_mux_sel = agg_sram_shared_floop_mux_sel;
assign agg_only_floop_restart = agg_sram_shared_floop_restart;
assign sram_only_loops_sram2tb_mux_sel = sram_tb_shared_loops_sram2tb_mux_sel;
assign sram_only_loops_sram2tb_restart = sram_tb_shared_loops_sram2tb_restart;
assign sram_only_t_read = sram_tb_shared_t_read_out;
assign ren_to_strg = |sram_tb_shared_t_read_out;
assign accessor_output = accessor_output_int;
strg_ub_agg_only agg_only (
  .agg_read(agg_only_agg_read),
  .agg_read_addr_gen_0_starting_addr(agg_only_agg_read_addr_gen_0_starting_addr),
  .agg_read_addr_gen_0_strides(agg_only_agg_read_addr_gen_0_strides),
  .agg_read_addr_gen_1_starting_addr(agg_only_agg_read_addr_gen_1_starting_addr),
  .agg_read_addr_gen_1_strides(agg_only_agg_read_addr_gen_1_strides),
  .agg_write_addr_gen_0_starting_addr(agg_only_agg_write_addr_gen_0_starting_addr),
  .agg_write_addr_gen_0_strides(agg_only_agg_write_addr_gen_0_strides),
  .agg_write_addr_gen_1_starting_addr(agg_only_agg_write_addr_gen_1_starting_addr),
  .agg_write_addr_gen_1_strides(agg_only_agg_write_addr_gen_1_strides),
  .agg_write_sched_gen_0_enable(agg_only_agg_write_sched_gen_0_enable),
  .agg_write_sched_gen_0_sched_addr_gen_starting_addr(agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr),
  .agg_write_sched_gen_0_sched_addr_gen_strides(agg_only_agg_write_sched_gen_0_sched_addr_gen_strides),
  .agg_write_sched_gen_1_enable(agg_only_agg_write_sched_gen_1_enable),
  .agg_write_sched_gen_1_sched_addr_gen_starting_addr(agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr),
  .agg_write_sched_gen_1_sched_addr_gen_strides(agg_only_agg_write_sched_gen_1_sched_addr_gen_strides),
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .data_in(data_in),
  .floop_mux_sel(agg_only_floop_mux_sel),
  .floop_restart(agg_only_floop_restart),
  .flush(flush),
  .loops_in2buf_0_dimensionality(agg_only_loops_in2buf_0_dimensionality),
  .loops_in2buf_0_ranges(agg_only_loops_in2buf_0_ranges),
  .loops_in2buf_1_dimensionality(agg_only_loops_in2buf_1_dimensionality),
  .loops_in2buf_1_ranges(agg_only_loops_in2buf_1_ranges),
  .rst_n(rst_n),
  .agg_data_out(agg_only_agg_data_out)
);

strg_ub_agg_sram_shared agg_sram_shared (
  .agg_read_sched_gen_0_enable(agg_sram_shared_agg_read_sched_gen_0_enable),
  .agg_read_sched_gen_0_sched_addr_gen_starting_addr(agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr),
  .agg_read_sched_gen_0_sched_addr_gen_strides(agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides),
  .agg_read_sched_gen_1_enable(agg_sram_shared_agg_read_sched_gen_1_enable),
  .agg_read_sched_gen_1_sched_addr_gen_starting_addr(agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr),
  .agg_read_sched_gen_1_sched_addr_gen_strides(agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides),
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .flush(flush),
  .loops_in2buf_autovec_write_0_dimensionality(agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality),
  .loops_in2buf_autovec_write_0_ranges(agg_sram_shared_loops_in2buf_autovec_write_0_ranges),
  .loops_in2buf_autovec_write_1_dimensionality(agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality),
  .loops_in2buf_autovec_write_1_ranges(agg_sram_shared_loops_in2buf_autovec_write_1_ranges),
  .rst_n(rst_n),
  .agg_read_out(agg_sram_shared_agg_read_out),
  .floop_mux_sel(agg_sram_shared_floop_mux_sel),
  .floop_restart(agg_sram_shared_floop_restart)
);

strg_ub_sram_only sram_only (
  .agg_data_out(agg_only_agg_data_out),
  .agg_read(agg_sram_shared_agg_read_out),
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .floop_mux_sel(agg_sram_shared_floop_mux_sel),
  .floop_restart(agg_sram_shared_floop_restart),
  .flush(flush),
  .input_addr_gen_0_starting_addr(sram_only_input_addr_gen_0_starting_addr),
  .input_addr_gen_0_strides(sram_only_input_addr_gen_0_strides),
  .input_addr_gen_1_starting_addr(sram_only_input_addr_gen_1_starting_addr),
  .input_addr_gen_1_strides(sram_only_input_addr_gen_1_strides),
  .loops_sram2tb_mux_sel(sram_only_loops_sram2tb_mux_sel),
  .loops_sram2tb_restart(sram_only_loops_sram2tb_restart),
  .output_addr_gen_0_starting_addr(sram_only_output_addr_gen_0_starting_addr),
  .output_addr_gen_0_strides(sram_only_output_addr_gen_0_strides),
  .output_addr_gen_1_starting_addr(sram_only_output_addr_gen_1_starting_addr),
  .output_addr_gen_1_strides(sram_only_output_addr_gen_1_strides),
  .rst_n(rst_n),
  .t_read(sram_only_t_read),
  .addr_to_sram(addr_out),
  .data_to_sram(data_to_strg),
  .wen_to_sram(wen_to_strg)
);

strg_ub_sram_tb_shared sram_tb_shared (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .flush(flush),
  .loops_buf2out_autovec_read_0_dimensionality(sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality),
  .loops_buf2out_autovec_read_0_ranges(sram_tb_shared_loops_buf2out_autovec_read_0_ranges),
  .loops_buf2out_autovec_read_1_dimensionality(sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality),
  .loops_buf2out_autovec_read_1_ranges(sram_tb_shared_loops_buf2out_autovec_read_1_ranges),
  .output_sched_gen_0_enable(sram_tb_shared_output_sched_gen_0_enable),
  .output_sched_gen_0_sched_addr_gen_starting_addr(sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr),
  .output_sched_gen_0_sched_addr_gen_strides(sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides),
  .output_sched_gen_1_enable(sram_tb_shared_output_sched_gen_1_enable),
  .output_sched_gen_1_sched_addr_gen_starting_addr(sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr),
  .output_sched_gen_1_sched_addr_gen_strides(sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides),
  .rst_n(rst_n),
  .loops_sram2tb_mux_sel(sram_tb_shared_loops_sram2tb_mux_sel),
  .loops_sram2tb_restart(sram_tb_shared_loops_sram2tb_restart),
  .t_read_out(sram_tb_shared_t_read_out)
);

strg_ub_tb_only tb_only (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .flush(flush),
  .loops_buf2out_read_0_dimensionality(tb_only_loops_buf2out_read_0_dimensionality),
  .loops_buf2out_read_0_ranges(tb_only_loops_buf2out_read_0_ranges),
  .loops_buf2out_read_1_dimensionality(tb_only_loops_buf2out_read_1_dimensionality),
  .loops_buf2out_read_1_ranges(tb_only_loops_buf2out_read_1_ranges),
  .loops_sram2tb_mux_sel(sram_tb_shared_loops_sram2tb_mux_sel),
  .loops_sram2tb_restart(sram_tb_shared_loops_sram2tb_restart),
  .rst_n(rst_n),
  .sram_read_data(data_from_strg),
  .t_read(sram_tb_shared_t_read_out),
  .tb_read_addr_gen_0_starting_addr(tb_only_tb_read_addr_gen_0_starting_addr),
  .tb_read_addr_gen_0_strides(tb_only_tb_read_addr_gen_0_strides),
  .tb_read_addr_gen_1_starting_addr(tb_only_tb_read_addr_gen_1_starting_addr),
  .tb_read_addr_gen_1_strides(tb_only_tb_read_addr_gen_1_strides),
  .tb_read_sched_gen_0_enable(tb_only_tb_read_sched_gen_0_enable),
  .tb_read_sched_gen_0_sched_addr_gen_starting_addr(tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr),
  .tb_read_sched_gen_0_sched_addr_gen_strides(tb_only_tb_read_sched_gen_0_sched_addr_gen_strides),
  .tb_read_sched_gen_1_enable(tb_only_tb_read_sched_gen_1_enable),
  .tb_read_sched_gen_1_sched_addr_gen_starting_addr(tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr),
  .tb_read_sched_gen_1_sched_addr_gen_strides(tb_only_tb_read_sched_gen_1_sched_addr_gen_strides),
  .tb_write_addr_gen_0_starting_addr(tb_only_tb_write_addr_gen_0_starting_addr),
  .tb_write_addr_gen_0_strides(tb_only_tb_write_addr_gen_0_strides),
  .tb_write_addr_gen_1_starting_addr(tb_only_tb_write_addr_gen_1_starting_addr),
  .tb_write_addr_gen_1_strides(tb_only_tb_write_addr_gen_1_strides),
  .accessor_output(accessor_output_int),
  .data_out(data_out_int)
);

Chain chain (
  .accessor_output(accessor_output_int),
  .chain_data_in(chain_data_in),
  .chain_en(chain_chain_en),
  .clk_en(clk_en),
  .curr_tile_data_out(data_out_int),
  .flush(flush),
  .data_out_tile(data_out)
);

endmodule   // strg_ub_vec

module strg_ub_vec_flat (
  input logic [0:0] [15:0] chain_data_in_f_0,
  input logic [0:0] [15:0] chain_data_in_f_1,
  input logic clk,
  input logic clk_en,
  input logic [3:0] [15:0] data_from_strg_lifted,
  input logic [0:0] [15:0] data_in_f_0,
  input logic [0:0] [15:0] data_in_f_1,
  input logic flush,
  input logic rst_n,
  input logic [3:0] strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides,
  input logic [3:0] strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides,
  input logic [3:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides,
  input logic [3:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides,
  input logic strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable,
  input logic [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides,
  input logic strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable,
  input logic [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality,
  input logic [5:0] [15:0] strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges,
  input logic [3:0] strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality,
  input logic [5:0] [15:0] strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges,
  input logic strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable,
  input logic [15:0] strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides,
  input logic strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable,
  input logic [15:0] strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality,
  input logic [5:0] [15:0] strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges,
  input logic [3:0] strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality,
  input logic [5:0] [15:0] strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges,
  input logic strg_ub_vec_inst_chain_chain_en,
  input logic [8:0] strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr,
  input logic [5:0] [8:0] strg_ub_vec_inst_sram_only_input_addr_gen_0_strides,
  input logic [8:0] strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr,
  input logic [5:0] [8:0] strg_ub_vec_inst_sram_only_input_addr_gen_1_strides,
  input logic [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr,
  input logic [5:0] [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_0_strides,
  input logic [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr,
  input logic [5:0] [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_1_strides,
  input logic [3:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality,
  input logic [5:0] [15:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges,
  input logic [3:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality,
  input logic [5:0] [15:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges,
  input logic strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable,
  input logic [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides,
  input logic strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable,
  input logic [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality,
  input logic [5:0] [15:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges,
  input logic [3:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality,
  input logic [5:0] [15:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides,
  input logic strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable,
  input logic [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides,
  input logic strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable,
  input logic [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides,
  output logic accessor_output_f_b_0,
  output logic accessor_output_f_b_1,
  output logic [8:0] addr_out_lifted,
  output logic [0:0] [15:0] data_out_f_0,
  output logic [0:0] [15:0] data_out_f_1,
  output logic [3:0] [15:0] data_to_strg_lifted,
  output logic ren_to_strg_lifted,
  output logic wen_to_strg_lifted
);

logic [1:0] strg_ub_vec_inst_accessor_output;
logic [1:0][15:0] strg_ub_vec_inst_chain_data_in;
logic [1:0][15:0] strg_ub_vec_inst_data_in;
logic [1:0][15:0] strg_ub_vec_inst_data_out;
assign strg_ub_vec_inst_chain_data_in[0] = chain_data_in_f_0;
assign strg_ub_vec_inst_chain_data_in[1] = chain_data_in_f_1;
assign strg_ub_vec_inst_data_in[0] = data_in_f_0;
assign strg_ub_vec_inst_data_in[1] = data_in_f_1;
assign accessor_output_f_b_0 = strg_ub_vec_inst_accessor_output[0];
assign accessor_output_f_b_1 = strg_ub_vec_inst_accessor_output[1];
assign data_out_f_0 = strg_ub_vec_inst_data_out[0];
assign data_out_f_1 = strg_ub_vec_inst_data_out[1];
strg_ub_vec strg_ub_vec_inst (
  .agg_only_agg_read_addr_gen_0_starting_addr(strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr),
  .agg_only_agg_read_addr_gen_0_strides(strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides),
  .agg_only_agg_read_addr_gen_1_starting_addr(strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr),
  .agg_only_agg_read_addr_gen_1_strides(strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides),
  .agg_only_agg_write_addr_gen_0_starting_addr(strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr),
  .agg_only_agg_write_addr_gen_0_strides(strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides),
  .agg_only_agg_write_addr_gen_1_starting_addr(strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr),
  .agg_only_agg_write_addr_gen_1_strides(strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides),
  .agg_only_agg_write_sched_gen_0_enable(strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable),
  .agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr),
  .agg_only_agg_write_sched_gen_0_sched_addr_gen_strides(strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides),
  .agg_only_agg_write_sched_gen_1_enable(strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable),
  .agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr),
  .agg_only_agg_write_sched_gen_1_sched_addr_gen_strides(strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides),
  .agg_only_loops_in2buf_0_dimensionality(strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality),
  .agg_only_loops_in2buf_0_ranges(strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges),
  .agg_only_loops_in2buf_1_dimensionality(strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality),
  .agg_only_loops_in2buf_1_ranges(strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges),
  .agg_sram_shared_agg_read_sched_gen_0_enable(strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable),
  .agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr),
  .agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides(strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides),
  .agg_sram_shared_agg_read_sched_gen_1_enable(strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable),
  .agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr),
  .agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides(strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides),
  .agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality(strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality),
  .agg_sram_shared_loops_in2buf_autovec_write_0_ranges(strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges),
  .agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality(strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality),
  .agg_sram_shared_loops_in2buf_autovec_write_1_ranges(strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges),
  .chain_chain_en(strg_ub_vec_inst_chain_chain_en),
  .chain_data_in(strg_ub_vec_inst_chain_data_in),
  .clk(clk),
  .clk_en(clk_en),
  .data_from_strg(data_from_strg_lifted),
  .data_in(strg_ub_vec_inst_data_in),
  .flush(flush),
  .rst_n(rst_n),
  .sram_only_input_addr_gen_0_starting_addr(strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr),
  .sram_only_input_addr_gen_0_strides(strg_ub_vec_inst_sram_only_input_addr_gen_0_strides),
  .sram_only_input_addr_gen_1_starting_addr(strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr),
  .sram_only_input_addr_gen_1_strides(strg_ub_vec_inst_sram_only_input_addr_gen_1_strides),
  .sram_only_output_addr_gen_0_starting_addr(strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr),
  .sram_only_output_addr_gen_0_strides(strg_ub_vec_inst_sram_only_output_addr_gen_0_strides),
  .sram_only_output_addr_gen_1_starting_addr(strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr),
  .sram_only_output_addr_gen_1_strides(strg_ub_vec_inst_sram_only_output_addr_gen_1_strides),
  .sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality),
  .sram_tb_shared_loops_buf2out_autovec_read_0_ranges(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges),
  .sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality),
  .sram_tb_shared_loops_buf2out_autovec_read_1_ranges(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges),
  .sram_tb_shared_output_sched_gen_0_enable(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable),
  .sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr),
  .sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides),
  .sram_tb_shared_output_sched_gen_1_enable(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable),
  .sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr),
  .sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides),
  .tb_only_loops_buf2out_read_0_dimensionality(strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality),
  .tb_only_loops_buf2out_read_0_ranges(strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges),
  .tb_only_loops_buf2out_read_1_dimensionality(strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality),
  .tb_only_loops_buf2out_read_1_ranges(strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges),
  .tb_only_tb_read_addr_gen_0_starting_addr(strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr),
  .tb_only_tb_read_addr_gen_0_strides(strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides),
  .tb_only_tb_read_addr_gen_1_starting_addr(strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr),
  .tb_only_tb_read_addr_gen_1_strides(strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides),
  .tb_only_tb_read_sched_gen_0_enable(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable),
  .tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr),
  .tb_only_tb_read_sched_gen_0_sched_addr_gen_strides(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides),
  .tb_only_tb_read_sched_gen_1_enable(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable),
  .tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr),
  .tb_only_tb_read_sched_gen_1_sched_addr_gen_strides(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides),
  .tb_only_tb_write_addr_gen_0_starting_addr(strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr),
  .tb_only_tb_write_addr_gen_0_strides(strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides),
  .tb_only_tb_write_addr_gen_1_starting_addr(strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr),
  .tb_only_tb_write_addr_gen_1_strides(strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides),
  .accessor_output(strg_ub_vec_inst_accessor_output),
  .addr_out(addr_out_lifted),
  .data_out(strg_ub_vec_inst_data_out),
  .data_to_strg(data_to_strg_lifted),
  .ren_to_strg(ren_to_strg_lifted),
  .wen_to_strg(wen_to_strg_lifted)
);

endmodule   // strg_ub_vec_flat


module LUT (
    input [7:0] lut,
    input bit0,
    input bit1,
    input bit2,
    output O,
    input CLK,
    input ASYNCRESET
);
wire bit_const_0_None_out;
wire [7:0] const_1_8_out;
wire [7:0] magma_Bits_8_and_inst0_out;
wire [7:0] magma_Bits_8_lshr_inst0_out;
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
coreir_const #(
    .value(8'h01),
    .width(8)
) const_1_8 (
    .out(const_1_8_out)
);
coreir_and #(
    .width(8)
) magma_Bits_8_and_inst0 (
    .in0(magma_Bits_8_lshr_inst0_out),
    .in1(const_1_8_out),
    .out(magma_Bits_8_and_inst0_out)
);
wire [7:0] magma_Bits_8_lshr_inst0_in1;
assign magma_Bits_8_lshr_inst0_in1 = {bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit2,bit1,bit0};
coreir_lshr #(
    .width(8)
) magma_Bits_8_lshr_inst0 (
    .in0(lut),
    .in1(magma_Bits_8_lshr_inst0_in1),
    .out(magma_Bits_8_lshr_inst0_out)
);
assign O = magma_Bits_8_and_inst0_out[0];
endmodule

module LTE (
    input [0:0] signed_,
    input [15:0] a,
    input [15:0] b,
    output [15:0] O0,
    output O1,
    output O2,
    output O3,
    output O4,
    output O5,
    input CLK,
    input ASYNCRESET
);
wire [0:0] Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [15:0] Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire bit_const_0_None_out;
wire [15:0] const_0_16_out;
wire [0:0] const_1_1_out;
wire magma_Bits_16_eq_inst0_out;
wire magma_Bits_1_eq_inst0_out;
wire magma_SInt_16_sle_inst0_out;
wire magma_UInt_16_ule_inst0_out;
coreir_mux #(
    .width(1)
) Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(magma_UInt_16_ule_inst0_out),
    .in1(magma_SInt_16_sle_inst0_out),
    .sel(magma_Bits_1_eq_inst0_out),
    .out(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(b),
    .in1(a),
    .sel(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .out(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_eq #(
    .width(16)
) magma_Bits_16_eq_inst0 (
    .in0(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(const_0_16_out),
    .out(magma_Bits_16_eq_inst0_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst0 (
    .in0(signed_),
    .in1(const_1_1_out),
    .out(magma_Bits_1_eq_inst0_out)
);
coreir_sle #(
    .width(16)
) magma_SInt_16_sle_inst0 (
    .in0(a),
    .in1(b),
    .out(magma_SInt_16_sle_inst0_out)
);
coreir_ule #(
    .width(16)
) magma_UInt_16_ule_inst0 (
    .in0(a),
    .in1(b),
    .out(magma_UInt_16_ule_inst0_out)
);
assign O0 = Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign O1 = Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign O2 = magma_Bits_16_eq_inst0_out;
assign O3 = Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15];
assign O4 = bit_const_0_None_out;
assign O5 = bit_const_0_None_out;
endmodule

module GTE (
    input [0:0] signed_,
    input [15:0] a,
    input [15:0] b,
    output [15:0] O0,
    output O1,
    output O2,
    output O3,
    output O4,
    output O5,
    input CLK,
    input ASYNCRESET
);
wire [0:0] Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [15:0] Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire bit_const_0_None_out;
wire [15:0] const_0_16_out;
wire [0:0] const_1_1_out;
wire magma_Bits_16_eq_inst0_out;
wire magma_Bits_1_eq_inst0_out;
wire magma_SInt_16_sge_inst0_out;
wire magma_UInt_16_uge_inst0_out;
coreir_mux #(
    .width(1)
) Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(magma_UInt_16_uge_inst0_out),
    .in1(magma_SInt_16_sge_inst0_out),
    .sel(magma_Bits_1_eq_inst0_out),
    .out(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(b),
    .in1(a),
    .sel(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .out(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_eq #(
    .width(16)
) magma_Bits_16_eq_inst0 (
    .in0(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(const_0_16_out),
    .out(magma_Bits_16_eq_inst0_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst0 (
    .in0(signed_),
    .in1(const_1_1_out),
    .out(magma_Bits_1_eq_inst0_out)
);
coreir_sge #(
    .width(16)
) magma_SInt_16_sge_inst0 (
    .in0(a),
    .in1(b),
    .out(magma_SInt_16_sge_inst0_out)
);
coreir_uge #(
    .width(16)
) magma_UInt_16_uge_inst0 (
    .in0(a),
    .in1(b),
    .out(magma_UInt_16_uge_inst0_out)
);
assign O0 = Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign O1 = Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign O2 = magma_Bits_16_eq_inst0_out;
assign O3 = Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15];
assign O4 = bit_const_0_None_out;
assign O5 = bit_const_0_None_out;
endmodule

module Decode98 (
    input [7:0] I,
    output O
);
wire [7:0] const_9_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h09),
    .width(8)
) const_9_8 (
    .out(const_9_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_9_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode88 (
    input [7:0] I,
    output O
);
wire [7:0] const_8_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h08),
    .width(8)
) const_8_8 (
    .out(const_8_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_8_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode78 (
    input [7:0] I,
    output O
);
wire [7:0] const_7_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h07),
    .width(8)
) const_7_8 (
    .out(const_7_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_7_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode68 (
    input [7:0] I,
    output O
);
wire [7:0] const_6_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h06),
    .width(8)
) const_6_8 (
    .out(const_6_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_6_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode58 (
    input [7:0] I,
    output O
);
wire [7:0] const_5_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h05),
    .width(8)
) const_5_8 (
    .out(const_5_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_5_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode48 (
    input [7:0] I,
    output O
);
wire [7:0] const_4_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h04),
    .width(8)
) const_4_8 (
    .out(const_4_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_4_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode38 (
    input [7:0] I,
    output O
);
wire [7:0] const_3_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h03),
    .width(8)
) const_3_8 (
    .out(const_3_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_3_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode28 (
    input [7:0] I,
    output O
);
wire [7:0] const_2_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h02),
    .width(8)
) const_2_8 (
    .out(const_2_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_2_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode18 (
    input [7:0] I,
    output O
);
wire [7:0] const_1_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h01),
    .width(8)
) const_1_8 (
    .out(const_1_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_1_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode148 (
    input [7:0] I,
    output O
);
wire [7:0] const_14_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0e),
    .width(8)
) const_14_8 (
    .out(const_14_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_14_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode138 (
    input [7:0] I,
    output O
);
wire [7:0] const_13_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0d),
    .width(8)
) const_13_8 (
    .out(const_13_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_13_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode128 (
    input [7:0] I,
    output O
);
wire [7:0] const_12_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0c),
    .width(8)
) const_12_8 (
    .out(const_12_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_12_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode118 (
    input [7:0] I,
    output O
);
wire [7:0] const_11_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0b),
    .width(8)
) const_11_8 (
    .out(const_11_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_11_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode108 (
    input [7:0] I,
    output O
);
wire [7:0] const_10_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0a),
    .width(8)
) const_10_8 (
    .out(const_10_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_10_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode08 (
    input [7:0] I,
    output O
);
wire [7:0] const_0_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_0_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module ConfigRegister_5_8_32_0 (
    input clk,
    input reset,
    output [4:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [4:0] Register_inst0_O;
wire [7:0] const_0_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq1 Register_inst0 (
    .I(config_data[4:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_0_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_9 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_9_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h09),
    .width(8)
) const_9_8 (
    .out(const_9_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_9_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_82 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_82_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h52),
    .width(8)
) const_82_8 (
    .out(const_82_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_82_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_81 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_81_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h51),
    .width(8)
) const_81_8 (
    .out(const_81_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_81_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_80 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_80_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h50),
    .width(8)
) const_80_8 (
    .out(const_80_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_80_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_8 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_8_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h08),
    .width(8)
) const_8_8 (
    .out(const_8_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_8_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_79 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_79_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h4f),
    .width(8)
) const_79_8 (
    .out(const_79_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_79_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_77 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_77_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h4d),
    .width(8)
) const_77_8 (
    .out(const_77_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_77_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_76 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_76_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h4c),
    .width(8)
) const_76_8 (
    .out(const_76_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_76_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_75 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_75_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h4b),
    .width(8)
) const_75_8 (
    .out(const_75_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_75_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_73 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_73_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h49),
    .width(8)
) const_73_8 (
    .out(const_73_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_73_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_72 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_72_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h48),
    .width(8)
) const_72_8 (
    .out(const_72_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_72_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_71 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_71_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h47),
    .width(8)
) const_71_8 (
    .out(const_71_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_71_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_70 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_70_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h46),
    .width(8)
) const_70_8 (
    .out(const_70_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_70_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_7 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_7_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h07),
    .width(8)
) const_7_8 (
    .out(const_7_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_7_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_68 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_68_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h44),
    .width(8)
) const_68_8 (
    .out(const_68_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_68_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_67 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_67_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h43),
    .width(8)
) const_67_8 (
    .out(const_67_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_67_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_66 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_66_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h42),
    .width(8)
) const_66_8 (
    .out(const_66_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_66_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_64 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_64_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h40),
    .width(8)
) const_64_8 (
    .out(const_64_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_64_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_63 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_63_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h3f),
    .width(8)
) const_63_8 (
    .out(const_63_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_63_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_62 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_62_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h3e),
    .width(8)
) const_62_8 (
    .out(const_62_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_62_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_60 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_60_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h3c),
    .width(8)
) const_60_8 (
    .out(const_60_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_60_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_6 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_6_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h06),
    .width(8)
) const_6_8 (
    .out(const_6_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_6_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_59 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_59_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h3b),
    .width(8)
) const_59_8 (
    .out(const_59_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_59_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_58 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_58_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h3a),
    .width(8)
) const_58_8 (
    .out(const_58_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_58_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_56 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_56_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h38),
    .width(8)
) const_56_8 (
    .out(const_56_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_56_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_55 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_55_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h37),
    .width(8)
) const_55_8 (
    .out(const_55_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_55_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_53 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_53_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h35),
    .width(8)
) const_53_8 (
    .out(const_53_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_53_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_52 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_52_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h34),
    .width(8)
) const_52_8 (
    .out(const_52_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_52_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_51 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_51_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h33),
    .width(8)
) const_51_8 (
    .out(const_51_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_51_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_5 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_5_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h05),
    .width(8)
) const_5_8 (
    .out(const_5_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_5_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_40 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_40_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h28),
    .width(8)
) const_40_8 (
    .out(const_40_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_40_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_4 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_4_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h04),
    .width(8)
) const_4_8 (
    .out(const_4_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_4_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_39 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_39_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h27),
    .width(8)
) const_39_8 (
    .out(const_39_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_39_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_37 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_37_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h25),
    .width(8)
) const_37_8 (
    .out(const_37_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_37_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_36 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_36_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h24),
    .width(8)
) const_36_8 (
    .out(const_36_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_36_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_35 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_35_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h23),
    .width(8)
) const_35_8 (
    .out(const_35_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_35_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_33 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_33_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h21),
    .width(8)
) const_33_8 (
    .out(const_33_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_33_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_32 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_32_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h20),
    .width(8)
) const_32_8 (
    .out(const_32_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_32_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_31 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_31_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h1f),
    .width(8)
) const_31_8 (
    .out(const_31_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_31_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_3 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_3_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h03),
    .width(8)
) const_3_8 (
    .out(const_3_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_3_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_29 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_29_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h1d),
    .width(8)
) const_29_8 (
    .out(const_29_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_29_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_28 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_28_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h1c),
    .width(8)
) const_28_8 (
    .out(const_28_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_28_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_27 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_27_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h1b),
    .width(8)
) const_27_8 (
    .out(const_27_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_27_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_25 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_25_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h19),
    .width(8)
) const_25_8 (
    .out(const_25_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_25_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_24 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_24_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h18),
    .width(8)
) const_24_8 (
    .out(const_24_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_24_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_22 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_22_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h16),
    .width(8)
) const_22_8 (
    .out(const_22_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_22_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_21 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_21_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h15),
    .width(8)
) const_21_8 (
    .out(const_21_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_21_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_20 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_20_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h14),
    .width(8)
) const_20_8 (
    .out(const_20_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_20_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_2 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_2_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h02),
    .width(8)
) const_2_8 (
    .out(const_2_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_2_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_18 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_18_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h12),
    .width(8)
) const_18_8 (
    .out(const_18_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_18_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_17 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_17_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h11),
    .width(8)
) const_17_8 (
    .out(const_17_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_17_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_16 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_16_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h10),
    .width(8)
) const_16_8 (
    .out(const_16_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_16_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_14 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_14_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0e),
    .width(8)
) const_14_8 (
    .out(const_14_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_14_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_13 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_13_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0d),
    .width(8)
) const_13_8 (
    .out(const_13_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_13_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_12 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_12_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0c),
    .width(8)
) const_12_8 (
    .out(const_12_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_12_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_10 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_10_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0a),
    .width(8)
) const_10_8 (
    .out(const_10_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_10_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_1 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_1_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h01),
    .width(8)
) const_1_8 (
    .out(const_1_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_1_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_0 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_0_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_0_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_31_8_32_50 (
    input clk,
    input reset,
    output [30:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [30:0] Register_inst0_O;
wire [7:0] const_50_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq12 Register_inst0 (
    .I(config_data[30:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h32),
    .width(8)
) const_50_8 (
    .out(const_50_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_50_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_30_8_32_1 (
    input clk,
    input reset,
    output [29:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [29:0] Register_inst0_O;
wire [7:0] const_1_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq6 Register_inst0 (
    .I(config_data[29:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h01),
    .width(8)
) const_1_8 (
    .out(const_1_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_1_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_27_8_32_83 (
    input clk,
    input reset,
    output [26:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [26:0] Register_inst0_O;
wire [7:0] const_83_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq11 Register_inst0 (
    .I(config_data[26:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h53),
    .width(8)
) const_83_8 (
    .out(const_83_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_83_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_27_8_32_49 (
    input clk,
    input reset,
    output [26:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [26:0] Register_inst0_O;
wire [7:0] const_49_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq11 Register_inst0 (
    .I(config_data[26:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h31),
    .width(8)
) const_49_8 (
    .out(const_49_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_49_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_27_8_32_48 (
    input clk,
    input reset,
    output [26:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [26:0] Register_inst0_O;
wire [7:0] const_48_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq11 Register_inst0 (
    .I(config_data[26:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h30),
    .width(8)
) const_48_8 (
    .out(const_48_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_48_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_27_8_32_47 (
    input clk,
    input reset,
    output [26:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [26:0] Register_inst0_O;
wire [7:0] const_47_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq11 Register_inst0 (
    .I(config_data[26:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h2f),
    .width(8)
) const_47_8 (
    .out(const_47_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_47_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_27_8_32_46 (
    input clk,
    input reset,
    output [26:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [26:0] Register_inst0_O;
wire [7:0] const_46_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq11 Register_inst0 (
    .I(config_data[26:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h2e),
    .width(8)
) const_46_8 (
    .out(const_46_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_46_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_27_8_32_45 (
    input clk,
    input reset,
    output [26:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [26:0] Register_inst0_O;
wire [7:0] const_45_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq11 Register_inst0 (
    .I(config_data[26:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h2d),
    .width(8)
) const_45_8 (
    .out(const_45_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_45_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_27_8_32_44 (
    input clk,
    input reset,
    output [26:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [26:0] Register_inst0_O;
wire [7:0] const_44_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq11 Register_inst0 (
    .I(config_data[26:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h2c),
    .width(8)
) const_44_8 (
    .out(const_44_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_44_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_27_8_32_43 (
    input clk,
    input reset,
    output [26:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [26:0] Register_inst0_O;
wire [7:0] const_43_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq11 Register_inst0 (
    .I(config_data[26:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h2b),
    .width(8)
) const_43_8 (
    .out(const_43_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_43_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_27_8_32_42 (
    input clk,
    input reset,
    output [26:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [26:0] Register_inst0_O;
wire [7:0] const_42_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq11 Register_inst0 (
    .I(config_data[26:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h2a),
    .width(8)
) const_42_8 (
    .out(const_42_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_42_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_26_8_32_41 (
    input clk,
    input reset,
    output [25:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [25:0] Register_inst0_O;
wire [7:0] const_41_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq10 Register_inst0 (
    .I(config_data[25:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h29),
    .width(8)
) const_41_8 (
    .out(const_41_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_41_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_25_8_32_74 (
    input clk,
    input reset,
    output [24:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [24:0] Register_inst0_O;
wire [7:0] const_74_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq8 Register_inst0 (
    .I(config_data[24:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h4a),
    .width(8)
) const_74_8 (
    .out(const_74_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_74_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_25_8_32_0 (
    input clk,
    input reset,
    output [24:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [24:0] Register_inst0_O;
wire [7:0] const_0_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq8 Register_inst0 (
    .I(config_data[24:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_0_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_24_8_32_0 (
    input clk,
    input reset,
    output [23:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [23:0] Register_inst0_O;
wire [7:0] const_0_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq2 Register_inst0 (
    .I(config_data[23:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_0_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_23_8_32_5 (
    input clk,
    input reset,
    output [22:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [22:0] Register_inst0_O;
wire [7:0] const_5_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq4 Register_inst0 (
    .I(config_data[22:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h05),
    .width(8)
) const_5_8 (
    .out(const_5_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_5_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_20_8_32_69 (
    input clk,
    input reset,
    output [19:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [19:0] Register_inst0_O;
wire [7:0] const_69_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq9 Register_inst0 (
    .I(config_data[19:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h45),
    .width(8)
) const_69_8 (
    .out(const_69_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_69_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_20_8_32_65 (
    input clk,
    input reset,
    output [19:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [19:0] Register_inst0_O;
wire [7:0] const_65_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq9 Register_inst0 (
    .I(config_data[19:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h41),
    .width(8)
) const_65_8 (
    .out(const_65_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_65_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_20_8_32_54 (
    input clk,
    input reset,
    output [19:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [19:0] Register_inst0_O;
wire [7:0] const_54_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq9 Register_inst0 (
    .I(config_data[19:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h36),
    .width(8)
) const_54_8 (
    .out(const_54_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_54_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_20_8_32_38 (
    input clk,
    input reset,
    output [19:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [19:0] Register_inst0_O;
wire [7:0] const_38_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq9 Register_inst0 (
    .I(config_data[19:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h26),
    .width(8)
) const_38_8 (
    .out(const_38_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_38_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_20_8_32_34 (
    input clk,
    input reset,
    output [19:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [19:0] Register_inst0_O;
wire [7:0] const_34_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq9 Register_inst0 (
    .I(config_data[19:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h22),
    .width(8)
) const_34_8 (
    .out(const_34_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_34_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_20_8_32_23 (
    input clk,
    input reset,
    output [19:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [19:0] Register_inst0_O;
wire [7:0] const_23_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq9 Register_inst0 (
    .I(config_data[19:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h17),
    .width(8)
) const_23_8 (
    .out(const_23_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_23_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_20_8_32_19 (
    input clk,
    input reset,
    output [19:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [19:0] Register_inst0_O;
wire [7:0] const_19_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq9 Register_inst0 (
    .I(config_data[19:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h13),
    .width(8)
) const_19_8 (
    .out(const_19_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_19_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_1_8_32_10 (
    input clk,
    input reset,
    output [0:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [0:0] Register_inst0_O;
wire [7:0] const_10_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq5 Register_inst0 (
    .I(config_data[0:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0a),
    .width(8)
) const_10_8 (
    .out(const_10_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_10_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_1_8_32_0 (
    input clk,
    input reset,
    output [0:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [0:0] Register_inst0_O;
wire [7:0] const_0_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq5 Register_inst0 (
    .I(config_data[0:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_0_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module PowerDomainConfigReg (
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [0:0] ps_en_out,
    output [31:0] read_config_data,
    input reset
);
wire ZextWrapper_1_32_inst0$bit_const_0_None_out;
wire [0:0] config_reg_0_O;
wire [0:0] ps_en_inst0_O;
corebit_const #(
    .value(1'b0)
) ZextWrapper_1_32_inst0$bit_const_0_None (
    .out(ZextWrapper_1_32_inst0$bit_const_0_None_out)
);
ConfigRegister_1_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ps_en ps_en_inst0 (
    .I(config_reg_0_O),
    .O(ps_en_inst0_O)
);
assign ps_en_out = ps_en_inst0_O;
assign read_config_data = {ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,config_reg_0_O[0]};
endmodule

module ConfigRegister_18_8_32_2 (
    input clk,
    input reset,
    output [17:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [17:0] Register_inst0_O;
wire [7:0] const_2_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq7 Register_inst0 (
    .I(config_data[17:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h02),
    .width(8)
) const_2_8 (
    .out(const_2_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_2_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module SB_ID0_5TRACKS_B1_PE (
    input [0:0] SB_T0_EAST_SB_IN_B1,
    output [0:0] SB_T0_EAST_SB_OUT_B1,
    input [0:0] SB_T0_NORTH_SB_IN_B1,
    output [0:0] SB_T0_NORTH_SB_OUT_B1,
    input [0:0] SB_T0_SOUTH_SB_IN_B1,
    output [0:0] SB_T0_SOUTH_SB_OUT_B1,
    input [0:0] SB_T0_WEST_SB_IN_B1,
    output [0:0] SB_T0_WEST_SB_OUT_B1,
    input [0:0] SB_T1_EAST_SB_IN_B1,
    output [0:0] SB_T1_EAST_SB_OUT_B1,
    input [0:0] SB_T1_NORTH_SB_IN_B1,
    output [0:0] SB_T1_NORTH_SB_OUT_B1,
    input [0:0] SB_T1_SOUTH_SB_IN_B1,
    output [0:0] SB_T1_SOUTH_SB_OUT_B1,
    input [0:0] SB_T1_WEST_SB_IN_B1,
    output [0:0] SB_T1_WEST_SB_OUT_B1,
    input [0:0] SB_T2_EAST_SB_IN_B1,
    output [0:0] SB_T2_EAST_SB_OUT_B1,
    input [0:0] SB_T2_NORTH_SB_IN_B1,
    output [0:0] SB_T2_NORTH_SB_OUT_B1,
    input [0:0] SB_T2_SOUTH_SB_IN_B1,
    output [0:0] SB_T2_SOUTH_SB_OUT_B1,
    input [0:0] SB_T2_WEST_SB_IN_B1,
    output [0:0] SB_T2_WEST_SB_OUT_B1,
    input [0:0] SB_T3_EAST_SB_IN_B1,
    output [0:0] SB_T3_EAST_SB_OUT_B1,
    input [0:0] SB_T3_NORTH_SB_IN_B1,
    output [0:0] SB_T3_NORTH_SB_OUT_B1,
    input [0:0] SB_T3_SOUTH_SB_IN_B1,
    output [0:0] SB_T3_SOUTH_SB_OUT_B1,
    input [0:0] SB_T3_WEST_SB_IN_B1,
    output [0:0] SB_T3_WEST_SB_OUT_B1,
    input [0:0] SB_T4_EAST_SB_IN_B1,
    output [0:0] SB_T4_EAST_SB_OUT_B1,
    input [0:0] SB_T4_NORTH_SB_IN_B1,
    output [0:0] SB_T4_NORTH_SB_OUT_B1,
    input [0:0] SB_T4_SOUTH_SB_IN_B1,
    output [0:0] SB_T4_SOUTH_SB_OUT_B1,
    input [0:0] SB_T4_WEST_SB_IN_B1,
    output [0:0] SB_T4_WEST_SB_OUT_B1,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    input [0:0] pe_outputs_1,
    output [31:0] read_config_data,
    input reset,
    input [0:0] stall,
    input [0:0] valid_out_pond
);
wire [0:0] Invert1_inst0_out;
wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1_O;
wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1_O;
wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1_O;
wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1_O;
wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1_O;
wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1_O;
wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1_O;
wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1_O;
wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1_O;
wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1_O;
wire [31:0] MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0_out;
wire [0:0] REG_T0_EAST_B1_O;
wire [0:0] REG_T0_NORTH_B1_O;
wire [0:0] REG_T0_SOUTH_B1_O;
wire [0:0] REG_T0_WEST_B1_O;
wire [0:0] REG_T1_EAST_B1_O;
wire [0:0] REG_T1_NORTH_B1_O;
wire [0:0] REG_T1_SOUTH_B1_O;
wire [0:0] REG_T1_WEST_B1_O;
wire [0:0] REG_T2_EAST_B1_O;
wire [0:0] REG_T2_NORTH_B1_O;
wire [0:0] REG_T2_SOUTH_B1_O;
wire [0:0] REG_T2_WEST_B1_O;
wire [0:0] REG_T3_EAST_B1_O;
wire [0:0] REG_T3_NORTH_B1_O;
wire [0:0] REG_T3_SOUTH_B1_O;
wire [0:0] REG_T3_WEST_B1_O;
wire [0:0] REG_T4_EAST_B1_O;
wire [0:0] REG_T4_NORTH_B1_O;
wire [0:0] REG_T4_SOUTH_B1_O;
wire [0:0] REG_T4_WEST_B1_O;
wire [0:0] RMUX_T0_EAST_B1_O;
wire [0:0] RMUX_T0_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T0_NORTH_B1_O;
wire [0:0] RMUX_T0_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T0_SOUTH_B1_O;
wire [0:0] RMUX_T0_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T0_WEST_B1_O;
wire [0:0] RMUX_T0_WEST_B1_sel_inst0_O;
wire [0:0] RMUX_T1_EAST_B1_O;
wire [0:0] RMUX_T1_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T1_NORTH_B1_O;
wire [0:0] RMUX_T1_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T1_SOUTH_B1_O;
wire [0:0] RMUX_T1_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T1_WEST_B1_O;
wire [0:0] RMUX_T1_WEST_B1_sel_inst0_O;
wire [0:0] RMUX_T2_EAST_B1_O;
wire [0:0] RMUX_T2_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T2_NORTH_B1_O;
wire [0:0] RMUX_T2_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T2_SOUTH_B1_O;
wire [0:0] RMUX_T2_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T2_WEST_B1_O;
wire [0:0] RMUX_T2_WEST_B1_sel_inst0_O;
wire [0:0] RMUX_T3_EAST_B1_O;
wire [0:0] RMUX_T3_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T3_NORTH_B1_O;
wire [0:0] RMUX_T3_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T3_SOUTH_B1_O;
wire [0:0] RMUX_T3_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T3_WEST_B1_O;
wire [0:0] RMUX_T3_WEST_B1_sel_inst0_O;
wire [0:0] RMUX_T4_EAST_B1_O;
wire [0:0] RMUX_T4_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T4_NORTH_B1_O;
wire [0:0] RMUX_T4_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T4_SOUTH_B1_O;
wire [0:0] RMUX_T4_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T4_WEST_B1_O;
wire [0:0] RMUX_T4_WEST_B1_sel_inst0_O;
wire [2:0] SB_T0_EAST_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T0_NORTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T0_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T0_WEST_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T1_EAST_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T1_NORTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T1_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T1_WEST_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T2_EAST_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T2_NORTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T2_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T2_WEST_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T3_EAST_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T3_NORTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T3_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T3_WEST_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T4_EAST_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T4_NORTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T4_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T4_WEST_SB_OUT_B1_sel_inst0_O;
wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1_O;
wire ZextWrapper_18_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_18_32_inst0$self_O_in;
wire ZextWrapper_30_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_30_32_inst0$self_O_in;
wire [0:0] and1_inst0_out;
wire [0:0] and1_inst1_out;
wire [0:0] and1_inst10_out;
wire [0:0] and1_inst11_out;
wire [0:0] and1_inst12_out;
wire [0:0] and1_inst13_out;
wire [0:0] and1_inst14_out;
wire [0:0] and1_inst15_out;
wire [0:0] and1_inst16_out;
wire [0:0] and1_inst17_out;
wire [0:0] and1_inst18_out;
wire [0:0] and1_inst19_out;
wire [0:0] and1_inst2_out;
wire [0:0] and1_inst3_out;
wire [0:0] and1_inst4_out;
wire [0:0] and1_inst5_out;
wire [0:0] and1_inst6_out;
wire [0:0] and1_inst7_out;
wire [0:0] and1_inst8_out;
wire [0:0] and1_inst9_out;
wire [31:0] config_reg_0_O;
wire [29:0] config_reg_1_O;
wire [17:0] config_reg_2_O;
wire [0:0] const_1_1_out;
wire coreir_eq_1_inst0_out;
wire coreir_eq_1_inst1_out;
wire coreir_eq_1_inst10_out;
wire coreir_eq_1_inst11_out;
wire coreir_eq_1_inst12_out;
wire coreir_eq_1_inst13_out;
wire coreir_eq_1_inst14_out;
wire coreir_eq_1_inst15_out;
wire coreir_eq_1_inst16_out;
wire coreir_eq_1_inst17_out;
wire coreir_eq_1_inst18_out;
wire coreir_eq_1_inst19_out;
wire coreir_eq_1_inst2_out;
wire coreir_eq_1_inst3_out;
wire coreir_eq_1_inst4_out;
wire coreir_eq_1_inst5_out;
wire coreir_eq_1_inst6_out;
wire coreir_eq_1_inst7_out;
wire coreir_eq_1_inst8_out;
wire coreir_eq_1_inst9_out;
wire [7:0] self_config_config_addr_out;
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(stall),
    .out(Invert1_inst0_out)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T0_EAST_SB_OUT_B1 (
    .I_0(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_1(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T0_EAST_SB_OUT_B1_O),
    .S(SB_T0_EAST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T0_NORTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_1(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T0_NORTH_SB_OUT_B1_O),
    .S(SB_T0_NORTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T0_SOUTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T0_SOUTH_SB_OUT_B1_O),
    .S(SB_T0_SOUTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T0_WEST_SB_OUT_B1 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T0_WEST_SB_OUT_B1_O),
    .S(SB_T0_WEST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T1_EAST_SB_OUT_B1 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_2(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T1_EAST_SB_OUT_B1_O),
    .S(SB_T1_EAST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T1_NORTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_1(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T1_NORTH_SB_OUT_B1_O),
    .S(SB_T1_NORTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T1_SOUTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_1(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T1_SOUTH_SB_OUT_B1_O),
    .S(SB_T1_SOUTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T1_WEST_SB_OUT_B1 (
    .I_0(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T1_WEST_SB_OUT_B1_O),
    .S(SB_T1_WEST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T2_EAST_SB_OUT_B1 (
    .I_0(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T2_EAST_SB_OUT_B1_O),
    .S(SB_T2_EAST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T2_NORTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_1(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T2_NORTH_SB_OUT_B1_O),
    .S(SB_T2_NORTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T2_SOUTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_1(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T2_SOUTH_SB_OUT_B1_O),
    .S(SB_T2_SOUTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T2_WEST_SB_OUT_B1 (
    .I_0(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T2_WEST_SB_OUT_B1_O),
    .S(SB_T2_WEST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T3_EAST_SB_OUT_B1 (
    .I_0(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T3_EAST_SB_OUT_B1_O),
    .S(SB_T3_EAST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T3_NORTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_1(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_2(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T3_NORTH_SB_OUT_B1_O),
    .S(SB_T3_NORTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T3_SOUTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_1(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T3_SOUTH_SB_OUT_B1_O),
    .S(SB_T3_SOUTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T3_WEST_SB_OUT_B1 (
    .I_0(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T3_WEST_SB_OUT_B1_O),
    .S(SB_T3_WEST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T4_EAST_SB_OUT_B1 (
    .I_0(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T4_EAST_SB_OUT_B1_O),
    .S(SB_T4_EAST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T4_NORTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_2(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T4_NORTH_SB_OUT_B1_O),
    .S(SB_T4_NORTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T4_SOUTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_1(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_2(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T4_SOUTH_SB_OUT_B1_O),
    .S(SB_T4_SOUTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_5_1 MUX_SB_T4_WEST_SB_OUT_B1 (
    .I_0(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_3(pe_outputs_1),
    .I_4(valid_out_pond),
    .O(MUX_SB_T4_WEST_SB_OUT_B1_O),
    .S(SB_T4_WEST_SB_OUT_B1_sel_inst0_O)
);
commonlib_muxn__N3__width32 MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0 (
    .in_data_0(config_reg_0_O),
    .in_data_1(ZextWrapper_30_32_inst0$self_O_in),
    .in_data_2(ZextWrapper_18_32_inst0$self_O_in),
    .in_sel(self_config_config_addr_out[1:0]),
    .out(MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0_out)
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_EAST_B1 (
    .I(MUX_SB_T0_EAST_SB_OUT_B1_O),
    .O(REG_T0_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst2_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_NORTH_B1 (
    .I(MUX_SB_T0_NORTH_SB_OUT_B1_O),
    .O(REG_T0_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst0_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_SOUTH_B1 (
    .I(MUX_SB_T0_SOUTH_SB_OUT_B1_O),
    .O(REG_T0_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst1_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_WEST_B1 (
    .I(MUX_SB_T0_WEST_SB_OUT_B1_O),
    .O(REG_T0_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst3_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_EAST_B1 (
    .I(MUX_SB_T1_EAST_SB_OUT_B1_O),
    .O(REG_T1_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst6_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_NORTH_B1 (
    .I(MUX_SB_T1_NORTH_SB_OUT_B1_O),
    .O(REG_T1_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst4_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_SOUTH_B1 (
    .I(MUX_SB_T1_SOUTH_SB_OUT_B1_O),
    .O(REG_T1_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst5_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_WEST_B1 (
    .I(MUX_SB_T1_WEST_SB_OUT_B1_O),
    .O(REG_T1_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst7_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_EAST_B1 (
    .I(MUX_SB_T2_EAST_SB_OUT_B1_O),
    .O(REG_T2_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst10_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_NORTH_B1 (
    .I(MUX_SB_T2_NORTH_SB_OUT_B1_O),
    .O(REG_T2_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst8_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_SOUTH_B1 (
    .I(MUX_SB_T2_SOUTH_SB_OUT_B1_O),
    .O(REG_T2_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst9_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_WEST_B1 (
    .I(MUX_SB_T2_WEST_SB_OUT_B1_O),
    .O(REG_T2_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst11_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T3_EAST_B1 (
    .I(MUX_SB_T3_EAST_SB_OUT_B1_O),
    .O(REG_T3_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst14_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T3_NORTH_B1 (
    .I(MUX_SB_T3_NORTH_SB_OUT_B1_O),
    .O(REG_T3_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst12_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T3_SOUTH_B1 (
    .I(MUX_SB_T3_SOUTH_SB_OUT_B1_O),
    .O(REG_T3_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst13_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T3_WEST_B1 (
    .I(MUX_SB_T3_WEST_SB_OUT_B1_O),
    .O(REG_T3_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst15_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T4_EAST_B1 (
    .I(MUX_SB_T4_EAST_SB_OUT_B1_O),
    .O(REG_T4_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst18_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T4_NORTH_B1 (
    .I(MUX_SB_T4_NORTH_SB_OUT_B1_O),
    .O(REG_T4_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst16_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T4_SOUTH_B1 (
    .I(MUX_SB_T4_SOUTH_SB_OUT_B1_O),
    .O(REG_T4_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst17_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T4_WEST_B1 (
    .I(MUX_SB_T4_WEST_SB_OUT_B1_O),
    .O(REG_T4_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst19_out[0])
);
MuxWrapperAOIImpl_2_1 RMUX_T0_EAST_B1 (
    .I_0(MUX_SB_T0_EAST_SB_OUT_B1_O),
    .I_1(REG_T0_EAST_B1_O),
    .O(RMUX_T0_EAST_B1_O),
    .S(RMUX_T0_EAST_B1_sel_inst0_O)
);
RMUX_T0_EAST_B1_sel RMUX_T0_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_EAST_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T0_NORTH_B1 (
    .I_0(MUX_SB_T0_NORTH_SB_OUT_B1_O),
    .I_1(REG_T0_NORTH_B1_O),
    .O(RMUX_T0_NORTH_B1_O),
    .S(RMUX_T0_NORTH_B1_sel_inst0_O)
);
RMUX_T0_NORTH_B1_sel RMUX_T0_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_NORTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T0_SOUTH_B1 (
    .I_0(MUX_SB_T0_SOUTH_SB_OUT_B1_O),
    .I_1(REG_T0_SOUTH_B1_O),
    .O(RMUX_T0_SOUTH_B1_O),
    .S(RMUX_T0_SOUTH_B1_sel_inst0_O)
);
RMUX_T0_SOUTH_B1_sel RMUX_T0_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_SOUTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T0_WEST_B1 (
    .I_0(MUX_SB_T0_WEST_SB_OUT_B1_O),
    .I_1(REG_T0_WEST_B1_O),
    .O(RMUX_T0_WEST_B1_O),
    .S(RMUX_T0_WEST_B1_sel_inst0_O)
);
RMUX_T0_WEST_B1_sel RMUX_T0_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_WEST_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T1_EAST_B1 (
    .I_0(MUX_SB_T1_EAST_SB_OUT_B1_O),
    .I_1(REG_T1_EAST_B1_O),
    .O(RMUX_T1_EAST_B1_O),
    .S(RMUX_T1_EAST_B1_sel_inst0_O)
);
RMUX_T1_EAST_B1_sel RMUX_T1_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_EAST_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T1_NORTH_B1 (
    .I_0(MUX_SB_T1_NORTH_SB_OUT_B1_O),
    .I_1(REG_T1_NORTH_B1_O),
    .O(RMUX_T1_NORTH_B1_O),
    .S(RMUX_T1_NORTH_B1_sel_inst0_O)
);
RMUX_T1_NORTH_B1_sel RMUX_T1_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_NORTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T1_SOUTH_B1 (
    .I_0(MUX_SB_T1_SOUTH_SB_OUT_B1_O),
    .I_1(REG_T1_SOUTH_B1_O),
    .O(RMUX_T1_SOUTH_B1_O),
    .S(RMUX_T1_SOUTH_B1_sel_inst0_O)
);
RMUX_T1_SOUTH_B1_sel RMUX_T1_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_SOUTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T1_WEST_B1 (
    .I_0(MUX_SB_T1_WEST_SB_OUT_B1_O),
    .I_1(REG_T1_WEST_B1_O),
    .O(RMUX_T1_WEST_B1_O),
    .S(RMUX_T1_WEST_B1_sel_inst0_O)
);
RMUX_T1_WEST_B1_sel RMUX_T1_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_WEST_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T2_EAST_B1 (
    .I_0(MUX_SB_T2_EAST_SB_OUT_B1_O),
    .I_1(REG_T2_EAST_B1_O),
    .O(RMUX_T2_EAST_B1_O),
    .S(RMUX_T2_EAST_B1_sel_inst0_O)
);
RMUX_T2_EAST_B1_sel RMUX_T2_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_EAST_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T2_NORTH_B1 (
    .I_0(MUX_SB_T2_NORTH_SB_OUT_B1_O),
    .I_1(REG_T2_NORTH_B1_O),
    .O(RMUX_T2_NORTH_B1_O),
    .S(RMUX_T2_NORTH_B1_sel_inst0_O)
);
RMUX_T2_NORTH_B1_sel RMUX_T2_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_NORTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T2_SOUTH_B1 (
    .I_0(MUX_SB_T2_SOUTH_SB_OUT_B1_O),
    .I_1(REG_T2_SOUTH_B1_O),
    .O(RMUX_T2_SOUTH_B1_O),
    .S(RMUX_T2_SOUTH_B1_sel_inst0_O)
);
RMUX_T2_SOUTH_B1_sel RMUX_T2_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_SOUTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T2_WEST_B1 (
    .I_0(MUX_SB_T2_WEST_SB_OUT_B1_O),
    .I_1(REG_T2_WEST_B1_O),
    .O(RMUX_T2_WEST_B1_O),
    .S(RMUX_T2_WEST_B1_sel_inst0_O)
);
RMUX_T2_WEST_B1_sel RMUX_T2_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_WEST_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T3_EAST_B1 (
    .I_0(MUX_SB_T3_EAST_SB_OUT_B1_O),
    .I_1(REG_T3_EAST_B1_O),
    .O(RMUX_T3_EAST_B1_O),
    .S(RMUX_T3_EAST_B1_sel_inst0_O)
);
RMUX_T3_EAST_B1_sel RMUX_T3_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_EAST_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T3_NORTH_B1 (
    .I_0(MUX_SB_T3_NORTH_SB_OUT_B1_O),
    .I_1(REG_T3_NORTH_B1_O),
    .O(RMUX_T3_NORTH_B1_O),
    .S(RMUX_T3_NORTH_B1_sel_inst0_O)
);
RMUX_T3_NORTH_B1_sel RMUX_T3_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_NORTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T3_SOUTH_B1 (
    .I_0(MUX_SB_T3_SOUTH_SB_OUT_B1_O),
    .I_1(REG_T3_SOUTH_B1_O),
    .O(RMUX_T3_SOUTH_B1_O),
    .S(RMUX_T3_SOUTH_B1_sel_inst0_O)
);
RMUX_T3_SOUTH_B1_sel RMUX_T3_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_SOUTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T3_WEST_B1 (
    .I_0(MUX_SB_T3_WEST_SB_OUT_B1_O),
    .I_1(REG_T3_WEST_B1_O),
    .O(RMUX_T3_WEST_B1_O),
    .S(RMUX_T3_WEST_B1_sel_inst0_O)
);
RMUX_T3_WEST_B1_sel RMUX_T3_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_WEST_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T4_EAST_B1 (
    .I_0(MUX_SB_T4_EAST_SB_OUT_B1_O),
    .I_1(REG_T4_EAST_B1_O),
    .O(RMUX_T4_EAST_B1_O),
    .S(RMUX_T4_EAST_B1_sel_inst0_O)
);
RMUX_T4_EAST_B1_sel RMUX_T4_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_EAST_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T4_NORTH_B1 (
    .I_0(MUX_SB_T4_NORTH_SB_OUT_B1_O),
    .I_1(REG_T4_NORTH_B1_O),
    .O(RMUX_T4_NORTH_B1_O),
    .S(RMUX_T4_NORTH_B1_sel_inst0_O)
);
RMUX_T4_NORTH_B1_sel RMUX_T4_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_NORTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T4_SOUTH_B1 (
    .I_0(MUX_SB_T4_SOUTH_SB_OUT_B1_O),
    .I_1(REG_T4_SOUTH_B1_O),
    .O(RMUX_T4_SOUTH_B1_O),
    .S(RMUX_T4_SOUTH_B1_sel_inst0_O)
);
RMUX_T4_SOUTH_B1_sel RMUX_T4_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_SOUTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T4_WEST_B1 (
    .I_0(MUX_SB_T4_WEST_SB_OUT_B1_O),
    .I_1(REG_T4_WEST_B1_O),
    .O(RMUX_T4_WEST_B1_O),
    .S(RMUX_T4_WEST_B1_sel_inst0_O)
);
RMUX_T4_WEST_B1_sel RMUX_T4_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_WEST_B1_sel_inst0_O)
);
SB_T0_EAST_SB_OUT_B1_sel SB_T0_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T0_NORTH_SB_OUT_B1_sel SB_T0_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T0_SOUTH_SB_OUT_B1_sel SB_T0_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T0_WEST_SB_OUT_B1_sel SB_T0_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_WEST_SB_OUT_B1_sel_inst0_O)
);
SB_T1_EAST_SB_OUT_B1_sel SB_T1_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T1_NORTH_SB_OUT_B1_sel SB_T1_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T1_SOUTH_SB_OUT_B1_sel SB_T1_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T1_WEST_SB_OUT_B1_sel SB_T1_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_WEST_SB_OUT_B1_sel_inst0_O)
);
SB_T2_EAST_SB_OUT_B1_sel SB_T2_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T2_NORTH_SB_OUT_B1_sel SB_T2_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T2_SOUTH_SB_OUT_B1_sel SB_T2_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T2_WEST_SB_OUT_B1_sel SB_T2_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_WEST_SB_OUT_B1_sel_inst0_O)
);
SB_T3_EAST_SB_OUT_B1_sel SB_T3_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T3_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T3_NORTH_SB_OUT_B1_sel SB_T3_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T3_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T3_SOUTH_SB_OUT_B1_sel SB_T3_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T3_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T3_WEST_SB_OUT_B1_sel SB_T3_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T3_WEST_SB_OUT_B1_sel_inst0_O)
);
SB_T4_EAST_SB_OUT_B1_sel SB_T4_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T4_NORTH_SB_OUT_B1_sel SB_T4_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T4_SOUTH_SB_OUT_B1_sel SB_T4_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T4_WEST_SB_OUT_B1_sel SB_T4_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_WEST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T0_EAST_SB_IN_B1 (
    .I(SB_T0_EAST_SB_IN_B1),
    .O(WIRE_SB_T0_EAST_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T0_NORTH_SB_IN_B1 (
    .I(SB_T0_NORTH_SB_IN_B1),
    .O(WIRE_SB_T0_NORTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T0_SOUTH_SB_IN_B1 (
    .I(SB_T0_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T0_WEST_SB_IN_B1 (
    .I(SB_T0_WEST_SB_IN_B1),
    .O(WIRE_SB_T0_WEST_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T1_EAST_SB_IN_B1 (
    .I(SB_T1_EAST_SB_IN_B1),
    .O(WIRE_SB_T1_EAST_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T1_NORTH_SB_IN_B1 (
    .I(SB_T1_NORTH_SB_IN_B1),
    .O(WIRE_SB_T1_NORTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T1_SOUTH_SB_IN_B1 (
    .I(SB_T1_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T1_WEST_SB_IN_B1 (
    .I(SB_T1_WEST_SB_IN_B1),
    .O(WIRE_SB_T1_WEST_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T2_EAST_SB_IN_B1 (
    .I(SB_T2_EAST_SB_IN_B1),
    .O(WIRE_SB_T2_EAST_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T2_NORTH_SB_IN_B1 (
    .I(SB_T2_NORTH_SB_IN_B1),
    .O(WIRE_SB_T2_NORTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T2_SOUTH_SB_IN_B1 (
    .I(SB_T2_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T2_WEST_SB_IN_B1 (
    .I(SB_T2_WEST_SB_IN_B1),
    .O(WIRE_SB_T2_WEST_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T3_EAST_SB_IN_B1 (
    .I(SB_T3_EAST_SB_IN_B1),
    .O(WIRE_SB_T3_EAST_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T3_NORTH_SB_IN_B1 (
    .I(SB_T3_NORTH_SB_IN_B1),
    .O(WIRE_SB_T3_NORTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T3_SOUTH_SB_IN_B1 (
    .I(SB_T3_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T3_WEST_SB_IN_B1 (
    .I(SB_T3_WEST_SB_IN_B1),
    .O(WIRE_SB_T3_WEST_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T4_EAST_SB_IN_B1 (
    .I(SB_T4_EAST_SB_IN_B1),
    .O(WIRE_SB_T4_EAST_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T4_NORTH_SB_IN_B1 (
    .I(SB_T4_NORTH_SB_IN_B1),
    .O(WIRE_SB_T4_NORTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T4_SOUTH_SB_IN_B1 (
    .I(SB_T4_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T4_WEST_SB_IN_B1 (
    .I(SB_T4_WEST_SB_IN_B1),
    .O(WIRE_SB_T4_WEST_SB_IN_B1_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_18_32_inst0$bit_const_0_None (
    .out(ZextWrapper_18_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_18_32_inst0$self_O_out;
assign ZextWrapper_18_32_inst0$self_O_out = {ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,config_reg_2_O};
mantle_wire__typeBitIn32 ZextWrapper_18_32_inst0$self_O (
    .in(ZextWrapper_18_32_inst0$self_O_in),
    .out(ZextWrapper_18_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_30_32_inst0$bit_const_0_None (
    .out(ZextWrapper_30_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_30_32_inst0$self_O_out;
assign ZextWrapper_30_32_inst0$self_O_out = {ZextWrapper_30_32_inst0$bit_const_0_None_out,ZextWrapper_30_32_inst0$bit_const_0_None_out,config_reg_1_O};
mantle_wire__typeBitIn32 ZextWrapper_30_32_inst0$self_O (
    .in(ZextWrapper_30_32_inst0$self_O_in),
    .out(ZextWrapper_30_32_inst0$self_O_out)
);
coreir_and #(
    .width(1)
) and1_inst0 (
    .in0(coreir_eq_1_inst0_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst0_out)
);
coreir_and #(
    .width(1)
) and1_inst1 (
    .in0(coreir_eq_1_inst1_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst1_out)
);
coreir_and #(
    .width(1)
) and1_inst10 (
    .in0(coreir_eq_1_inst10_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst10_out)
);
coreir_and #(
    .width(1)
) and1_inst11 (
    .in0(coreir_eq_1_inst11_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst11_out)
);
coreir_and #(
    .width(1)
) and1_inst12 (
    .in0(coreir_eq_1_inst12_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst12_out)
);
coreir_and #(
    .width(1)
) and1_inst13 (
    .in0(coreir_eq_1_inst13_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst13_out)
);
coreir_and #(
    .width(1)
) and1_inst14 (
    .in0(coreir_eq_1_inst14_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst14_out)
);
coreir_and #(
    .width(1)
) and1_inst15 (
    .in0(coreir_eq_1_inst15_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst15_out)
);
coreir_and #(
    .width(1)
) and1_inst16 (
    .in0(coreir_eq_1_inst16_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst16_out)
);
coreir_and #(
    .width(1)
) and1_inst17 (
    .in0(coreir_eq_1_inst17_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst17_out)
);
coreir_and #(
    .width(1)
) and1_inst18 (
    .in0(coreir_eq_1_inst18_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst18_out)
);
coreir_and #(
    .width(1)
) and1_inst19 (
    .in0(coreir_eq_1_inst19_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst19_out)
);
coreir_and #(
    .width(1)
) and1_inst2 (
    .in0(coreir_eq_1_inst2_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst2_out)
);
coreir_and #(
    .width(1)
) and1_inst3 (
    .in0(coreir_eq_1_inst3_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst3_out)
);
coreir_and #(
    .width(1)
) and1_inst4 (
    .in0(coreir_eq_1_inst4_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst4_out)
);
coreir_and #(
    .width(1)
) and1_inst5 (
    .in0(coreir_eq_1_inst5_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst5_out)
);
coreir_and #(
    .width(1)
) and1_inst6 (
    .in0(coreir_eq_1_inst6_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst6_out)
);
coreir_and #(
    .width(1)
) and1_inst7 (
    .in0(coreir_eq_1_inst7_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst7_out)
);
coreir_and #(
    .width(1)
) and1_inst8 (
    .in0(coreir_eq_1_inst8_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst8_out)
);
coreir_and #(
    .width(1)
) and1_inst9 (
    .in0(coreir_eq_1_inst9_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst9_out)
);
wire [7:0] config_reg_0_config_addr;
assign config_reg_0_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2],self_config_config_addr_out[1:0]};
ConfigRegister_32_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_reg_0_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_1_config_addr;
assign config_reg_1_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2],self_config_config_addr_out[1:0]};
ConfigRegister_30_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_reg_1_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_2_config_addr;
assign config_reg_2_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2],self_config_config_addr_out[1:0]};
ConfigRegister_18_8_32_2 config_reg_2 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_2_O),
    .config_addr(config_reg_2_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst0 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst0_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst1 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst10 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst10_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst11 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst11_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst12 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst12_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst13 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst13_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst14 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst14_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst15 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst15_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst16 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst16_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst17 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst17_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst18 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst18_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst19 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst19_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst2 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst2_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst3 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst3_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst4 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst4_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst5 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst5_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst6 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst6_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst7 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst7_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst8 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst8_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst9 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst9_out)
);
mantle_wire__typeBit8 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
assign SB_T0_EAST_SB_OUT_B1 = RMUX_T0_EAST_B1_O;
assign SB_T0_NORTH_SB_OUT_B1 = RMUX_T0_NORTH_B1_O;
assign SB_T0_SOUTH_SB_OUT_B1 = RMUX_T0_SOUTH_B1_O;
assign SB_T0_WEST_SB_OUT_B1 = RMUX_T0_WEST_B1_O;
assign SB_T1_EAST_SB_OUT_B1 = RMUX_T1_EAST_B1_O;
assign SB_T1_NORTH_SB_OUT_B1 = RMUX_T1_NORTH_B1_O;
assign SB_T1_SOUTH_SB_OUT_B1 = RMUX_T1_SOUTH_B1_O;
assign SB_T1_WEST_SB_OUT_B1 = RMUX_T1_WEST_B1_O;
assign SB_T2_EAST_SB_OUT_B1 = RMUX_T2_EAST_B1_O;
assign SB_T2_NORTH_SB_OUT_B1 = RMUX_T2_NORTH_B1_O;
assign SB_T2_SOUTH_SB_OUT_B1 = RMUX_T2_SOUTH_B1_O;
assign SB_T2_WEST_SB_OUT_B1 = RMUX_T2_WEST_B1_O;
assign SB_T3_EAST_SB_OUT_B1 = RMUX_T3_EAST_B1_O;
assign SB_T3_NORTH_SB_OUT_B1 = RMUX_T3_NORTH_B1_O;
assign SB_T3_SOUTH_SB_OUT_B1 = RMUX_T3_SOUTH_B1_O;
assign SB_T3_WEST_SB_OUT_B1 = RMUX_T3_WEST_B1_O;
assign SB_T4_EAST_SB_OUT_B1 = RMUX_T4_EAST_B1_O;
assign SB_T4_NORTH_SB_OUT_B1 = RMUX_T4_NORTH_B1_O;
assign SB_T4_SOUTH_SB_OUT_B1 = RMUX_T4_SOUTH_B1_O;
assign SB_T4_WEST_SB_OUT_B1 = RMUX_T4_WEST_B1_O;
assign read_config_data = MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0_out;
endmodule

module SB_ID0_5TRACKS_B1_MemCore (
    input [0:0] SB_T0_EAST_SB_IN_B1,
    output [0:0] SB_T0_EAST_SB_OUT_B1,
    input [0:0] SB_T0_NORTH_SB_IN_B1,
    output [0:0] SB_T0_NORTH_SB_OUT_B1,
    input [0:0] SB_T0_SOUTH_SB_IN_B1,
    output [0:0] SB_T0_SOUTH_SB_OUT_B1,
    input [0:0] SB_T0_WEST_SB_IN_B1,
    output [0:0] SB_T0_WEST_SB_OUT_B1,
    input [0:0] SB_T1_EAST_SB_IN_B1,
    output [0:0] SB_T1_EAST_SB_OUT_B1,
    input [0:0] SB_T1_NORTH_SB_IN_B1,
    output [0:0] SB_T1_NORTH_SB_OUT_B1,
    input [0:0] SB_T1_SOUTH_SB_IN_B1,
    output [0:0] SB_T1_SOUTH_SB_OUT_B1,
    input [0:0] SB_T1_WEST_SB_IN_B1,
    output [0:0] SB_T1_WEST_SB_OUT_B1,
    input [0:0] SB_T2_EAST_SB_IN_B1,
    output [0:0] SB_T2_EAST_SB_OUT_B1,
    input [0:0] SB_T2_NORTH_SB_IN_B1,
    output [0:0] SB_T2_NORTH_SB_OUT_B1,
    input [0:0] SB_T2_SOUTH_SB_IN_B1,
    output [0:0] SB_T2_SOUTH_SB_OUT_B1,
    input [0:0] SB_T2_WEST_SB_IN_B1,
    output [0:0] SB_T2_WEST_SB_OUT_B1,
    input [0:0] SB_T3_EAST_SB_IN_B1,
    output [0:0] SB_T3_EAST_SB_OUT_B1,
    input [0:0] SB_T3_NORTH_SB_IN_B1,
    output [0:0] SB_T3_NORTH_SB_OUT_B1,
    input [0:0] SB_T3_SOUTH_SB_IN_B1,
    output [0:0] SB_T3_SOUTH_SB_OUT_B1,
    input [0:0] SB_T3_WEST_SB_IN_B1,
    output [0:0] SB_T3_WEST_SB_OUT_B1,
    input [0:0] SB_T4_EAST_SB_IN_B1,
    output [0:0] SB_T4_EAST_SB_OUT_B1,
    input [0:0] SB_T4_NORTH_SB_IN_B1,
    output [0:0] SB_T4_NORTH_SB_OUT_B1,
    input [0:0] SB_T4_SOUTH_SB_IN_B1,
    output [0:0] SB_T4_SOUTH_SB_OUT_B1,
    input [0:0] SB_T4_WEST_SB_IN_B1,
    output [0:0] SB_T4_WEST_SB_OUT_B1,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    input [0:0] output_width_1_num_0,
    input [0:0] output_width_1_num_1,
    input [0:0] output_width_1_num_2,
    input [0:0] output_width_1_num_3,
    output [31:0] read_config_data,
    input reset,
    input [0:0] stall
);
wire [0:0] Invert1_inst0_out;
wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1_O;
wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1_O;
wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1_O;
wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1_O;
wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1_O;
wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1_O;
wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1_O;
wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1_O;
wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1_O;
wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1_O;
wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1_O;
wire [31:0] MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0_out;
wire [0:0] REG_T0_EAST_B1_O;
wire [0:0] REG_T0_NORTH_B1_O;
wire [0:0] REG_T0_SOUTH_B1_O;
wire [0:0] REG_T0_WEST_B1_O;
wire [0:0] REG_T1_EAST_B1_O;
wire [0:0] REG_T1_NORTH_B1_O;
wire [0:0] REG_T1_SOUTH_B1_O;
wire [0:0] REG_T1_WEST_B1_O;
wire [0:0] REG_T2_EAST_B1_O;
wire [0:0] REG_T2_NORTH_B1_O;
wire [0:0] REG_T2_SOUTH_B1_O;
wire [0:0] REG_T2_WEST_B1_O;
wire [0:0] REG_T3_EAST_B1_O;
wire [0:0] REG_T3_NORTH_B1_O;
wire [0:0] REG_T3_SOUTH_B1_O;
wire [0:0] REG_T3_WEST_B1_O;
wire [0:0] REG_T4_EAST_B1_O;
wire [0:0] REG_T4_NORTH_B1_O;
wire [0:0] REG_T4_SOUTH_B1_O;
wire [0:0] REG_T4_WEST_B1_O;
wire [0:0] RMUX_T0_EAST_B1_O;
wire [0:0] RMUX_T0_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T0_NORTH_B1_O;
wire [0:0] RMUX_T0_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T0_SOUTH_B1_O;
wire [0:0] RMUX_T0_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T0_WEST_B1_O;
wire [0:0] RMUX_T0_WEST_B1_sel_inst0_O;
wire [0:0] RMUX_T1_EAST_B1_O;
wire [0:0] RMUX_T1_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T1_NORTH_B1_O;
wire [0:0] RMUX_T1_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T1_SOUTH_B1_O;
wire [0:0] RMUX_T1_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T1_WEST_B1_O;
wire [0:0] RMUX_T1_WEST_B1_sel_inst0_O;
wire [0:0] RMUX_T2_EAST_B1_O;
wire [0:0] RMUX_T2_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T2_NORTH_B1_O;
wire [0:0] RMUX_T2_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T2_SOUTH_B1_O;
wire [0:0] RMUX_T2_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T2_WEST_B1_O;
wire [0:0] RMUX_T2_WEST_B1_sel_inst0_O;
wire [0:0] RMUX_T3_EAST_B1_O;
wire [0:0] RMUX_T3_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T3_NORTH_B1_O;
wire [0:0] RMUX_T3_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T3_SOUTH_B1_O;
wire [0:0] RMUX_T3_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T3_WEST_B1_O;
wire [0:0] RMUX_T3_WEST_B1_sel_inst0_O;
wire [0:0] RMUX_T4_EAST_B1_O;
wire [0:0] RMUX_T4_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T4_NORTH_B1_O;
wire [0:0] RMUX_T4_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T4_SOUTH_B1_O;
wire [0:0] RMUX_T4_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T4_WEST_B1_O;
wire [0:0] RMUX_T4_WEST_B1_sel_inst0_O;
wire [2:0] SB_T0_EAST_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T0_NORTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T0_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T0_WEST_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T1_EAST_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T1_NORTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T1_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T1_WEST_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T2_EAST_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T2_NORTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T2_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T2_WEST_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T3_EAST_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T3_NORTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T3_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T3_WEST_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T4_EAST_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T4_NORTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T4_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [2:0] SB_T4_WEST_SB_OUT_B1_sel_inst0_O;
wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1_O;
wire ZextWrapper_18_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_18_32_inst0$self_O_in;
wire ZextWrapper_30_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_30_32_inst0$self_O_in;
wire [0:0] and1_inst0_out;
wire [0:0] and1_inst1_out;
wire [0:0] and1_inst10_out;
wire [0:0] and1_inst11_out;
wire [0:0] and1_inst12_out;
wire [0:0] and1_inst13_out;
wire [0:0] and1_inst14_out;
wire [0:0] and1_inst15_out;
wire [0:0] and1_inst16_out;
wire [0:0] and1_inst17_out;
wire [0:0] and1_inst18_out;
wire [0:0] and1_inst19_out;
wire [0:0] and1_inst2_out;
wire [0:0] and1_inst3_out;
wire [0:0] and1_inst4_out;
wire [0:0] and1_inst5_out;
wire [0:0] and1_inst6_out;
wire [0:0] and1_inst7_out;
wire [0:0] and1_inst8_out;
wire [0:0] and1_inst9_out;
wire [31:0] config_reg_0_O;
wire [29:0] config_reg_1_O;
wire [17:0] config_reg_2_O;
wire [0:0] const_1_1_out;
wire coreir_eq_1_inst0_out;
wire coreir_eq_1_inst1_out;
wire coreir_eq_1_inst10_out;
wire coreir_eq_1_inst11_out;
wire coreir_eq_1_inst12_out;
wire coreir_eq_1_inst13_out;
wire coreir_eq_1_inst14_out;
wire coreir_eq_1_inst15_out;
wire coreir_eq_1_inst16_out;
wire coreir_eq_1_inst17_out;
wire coreir_eq_1_inst18_out;
wire coreir_eq_1_inst19_out;
wire coreir_eq_1_inst2_out;
wire coreir_eq_1_inst3_out;
wire coreir_eq_1_inst4_out;
wire coreir_eq_1_inst5_out;
wire coreir_eq_1_inst6_out;
wire coreir_eq_1_inst7_out;
wire coreir_eq_1_inst8_out;
wire coreir_eq_1_inst9_out;
wire [7:0] self_config_config_addr_out;
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(stall),
    .out(Invert1_inst0_out)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T0_EAST_SB_OUT_B1 (
    .I_0(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_1(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T0_EAST_SB_OUT_B1_O),
    .S(SB_T0_EAST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T0_NORTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_1(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T0_NORTH_SB_OUT_B1_O),
    .S(SB_T0_NORTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T0_SOUTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T0_SOUTH_SB_OUT_B1_O),
    .S(SB_T0_SOUTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T0_WEST_SB_OUT_B1 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T0_WEST_SB_OUT_B1_O),
    .S(SB_T0_WEST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T1_EAST_SB_OUT_B1 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_2(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T1_EAST_SB_OUT_B1_O),
    .S(SB_T1_EAST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T1_NORTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_1(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T1_NORTH_SB_OUT_B1_O),
    .S(SB_T1_NORTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T1_SOUTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_1(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T1_SOUTH_SB_OUT_B1_O),
    .S(SB_T1_SOUTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T1_WEST_SB_OUT_B1 (
    .I_0(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T1_WEST_SB_OUT_B1_O),
    .S(SB_T1_WEST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T2_EAST_SB_OUT_B1 (
    .I_0(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T2_EAST_SB_OUT_B1_O),
    .S(SB_T2_EAST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T2_NORTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_1(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T2_NORTH_SB_OUT_B1_O),
    .S(SB_T2_NORTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T2_SOUTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_1(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T2_SOUTH_SB_OUT_B1_O),
    .S(SB_T2_SOUTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T2_WEST_SB_OUT_B1 (
    .I_0(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T2_WEST_SB_OUT_B1_O),
    .S(SB_T2_WEST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T3_EAST_SB_OUT_B1 (
    .I_0(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T3_EAST_SB_OUT_B1_O),
    .S(SB_T3_EAST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T3_NORTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_1(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_2(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T3_NORTH_SB_OUT_B1_O),
    .S(SB_T3_NORTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T3_SOUTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_1(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T3_SOUTH_SB_OUT_B1_O),
    .S(SB_T3_SOUTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T3_WEST_SB_OUT_B1 (
    .I_0(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T3_WEST_SB_OUT_B1_O),
    .S(SB_T3_WEST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T4_EAST_SB_OUT_B1 (
    .I_0(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T4_EAST_SB_OUT_B1_O),
    .S(SB_T4_EAST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T4_NORTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_2(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T4_NORTH_SB_OUT_B1_O),
    .S(SB_T4_NORTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T4_SOUTH_SB_OUT_B1 (
    .I_0(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_1(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_2(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T4_SOUTH_SB_OUT_B1_O),
    .S(SB_T4_SOUTH_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_7_1 MUX_SB_T4_WEST_SB_OUT_B1 (
    .I_0(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_2(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_3(output_width_1_num_0),
    .I_4(output_width_1_num_1),
    .I_5(output_width_1_num_2),
    .I_6(output_width_1_num_3),
    .O(MUX_SB_T4_WEST_SB_OUT_B1_O),
    .S(SB_T4_WEST_SB_OUT_B1_sel_inst0_O)
);
commonlib_muxn__N3__width32 MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0 (
    .in_data_0(config_reg_0_O),
    .in_data_1(ZextWrapper_30_32_inst0$self_O_in),
    .in_data_2(ZextWrapper_18_32_inst0$self_O_in),
    .in_sel(self_config_config_addr_out[1:0]),
    .out(MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0_out)
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_EAST_B1 (
    .I(MUX_SB_T0_EAST_SB_OUT_B1_O),
    .O(REG_T0_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst2_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_NORTH_B1 (
    .I(MUX_SB_T0_NORTH_SB_OUT_B1_O),
    .O(REG_T0_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst0_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_SOUTH_B1 (
    .I(MUX_SB_T0_SOUTH_SB_OUT_B1_O),
    .O(REG_T0_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst1_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_WEST_B1 (
    .I(MUX_SB_T0_WEST_SB_OUT_B1_O),
    .O(REG_T0_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst3_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_EAST_B1 (
    .I(MUX_SB_T1_EAST_SB_OUT_B1_O),
    .O(REG_T1_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst6_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_NORTH_B1 (
    .I(MUX_SB_T1_NORTH_SB_OUT_B1_O),
    .O(REG_T1_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst4_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_SOUTH_B1 (
    .I(MUX_SB_T1_SOUTH_SB_OUT_B1_O),
    .O(REG_T1_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst5_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_WEST_B1 (
    .I(MUX_SB_T1_WEST_SB_OUT_B1_O),
    .O(REG_T1_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst7_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_EAST_B1 (
    .I(MUX_SB_T2_EAST_SB_OUT_B1_O),
    .O(REG_T2_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst10_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_NORTH_B1 (
    .I(MUX_SB_T2_NORTH_SB_OUT_B1_O),
    .O(REG_T2_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst8_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_SOUTH_B1 (
    .I(MUX_SB_T2_SOUTH_SB_OUT_B1_O),
    .O(REG_T2_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst9_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_WEST_B1 (
    .I(MUX_SB_T2_WEST_SB_OUT_B1_O),
    .O(REG_T2_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst11_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T3_EAST_B1 (
    .I(MUX_SB_T3_EAST_SB_OUT_B1_O),
    .O(REG_T3_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst14_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T3_NORTH_B1 (
    .I(MUX_SB_T3_NORTH_SB_OUT_B1_O),
    .O(REG_T3_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst12_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T3_SOUTH_B1 (
    .I(MUX_SB_T3_SOUTH_SB_OUT_B1_O),
    .O(REG_T3_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst13_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T3_WEST_B1 (
    .I(MUX_SB_T3_WEST_SB_OUT_B1_O),
    .O(REG_T3_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst15_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T4_EAST_B1 (
    .I(MUX_SB_T4_EAST_SB_OUT_B1_O),
    .O(REG_T4_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst18_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T4_NORTH_B1 (
    .I(MUX_SB_T4_NORTH_SB_OUT_B1_O),
    .O(REG_T4_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst16_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T4_SOUTH_B1 (
    .I(MUX_SB_T4_SOUTH_SB_OUT_B1_O),
    .O(REG_T4_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst17_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T4_WEST_B1 (
    .I(MUX_SB_T4_WEST_SB_OUT_B1_O),
    .O(REG_T4_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst19_out[0])
);
MuxWrapperAOIImpl_2_1 RMUX_T0_EAST_B1 (
    .I_0(MUX_SB_T0_EAST_SB_OUT_B1_O),
    .I_1(REG_T0_EAST_B1_O),
    .O(RMUX_T0_EAST_B1_O),
    .S(RMUX_T0_EAST_B1_sel_inst0_O)
);
RMUX_T0_EAST_B1_sel RMUX_T0_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_EAST_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T0_NORTH_B1 (
    .I_0(MUX_SB_T0_NORTH_SB_OUT_B1_O),
    .I_1(REG_T0_NORTH_B1_O),
    .O(RMUX_T0_NORTH_B1_O),
    .S(RMUX_T0_NORTH_B1_sel_inst0_O)
);
RMUX_T0_NORTH_B1_sel RMUX_T0_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_NORTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T0_SOUTH_B1 (
    .I_0(MUX_SB_T0_SOUTH_SB_OUT_B1_O),
    .I_1(REG_T0_SOUTH_B1_O),
    .O(RMUX_T0_SOUTH_B1_O),
    .S(RMUX_T0_SOUTH_B1_sel_inst0_O)
);
RMUX_T0_SOUTH_B1_sel RMUX_T0_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_SOUTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T0_WEST_B1 (
    .I_0(MUX_SB_T0_WEST_SB_OUT_B1_O),
    .I_1(REG_T0_WEST_B1_O),
    .O(RMUX_T0_WEST_B1_O),
    .S(RMUX_T0_WEST_B1_sel_inst0_O)
);
RMUX_T0_WEST_B1_sel RMUX_T0_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_WEST_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T1_EAST_B1 (
    .I_0(MUX_SB_T1_EAST_SB_OUT_B1_O),
    .I_1(REG_T1_EAST_B1_O),
    .O(RMUX_T1_EAST_B1_O),
    .S(RMUX_T1_EAST_B1_sel_inst0_O)
);
RMUX_T1_EAST_B1_sel RMUX_T1_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_EAST_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T1_NORTH_B1 (
    .I_0(MUX_SB_T1_NORTH_SB_OUT_B1_O),
    .I_1(REG_T1_NORTH_B1_O),
    .O(RMUX_T1_NORTH_B1_O),
    .S(RMUX_T1_NORTH_B1_sel_inst0_O)
);
RMUX_T1_NORTH_B1_sel RMUX_T1_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_NORTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T1_SOUTH_B1 (
    .I_0(MUX_SB_T1_SOUTH_SB_OUT_B1_O),
    .I_1(REG_T1_SOUTH_B1_O),
    .O(RMUX_T1_SOUTH_B1_O),
    .S(RMUX_T1_SOUTH_B1_sel_inst0_O)
);
RMUX_T1_SOUTH_B1_sel RMUX_T1_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_SOUTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T1_WEST_B1 (
    .I_0(MUX_SB_T1_WEST_SB_OUT_B1_O),
    .I_1(REG_T1_WEST_B1_O),
    .O(RMUX_T1_WEST_B1_O),
    .S(RMUX_T1_WEST_B1_sel_inst0_O)
);
RMUX_T1_WEST_B1_sel RMUX_T1_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_WEST_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T2_EAST_B1 (
    .I_0(MUX_SB_T2_EAST_SB_OUT_B1_O),
    .I_1(REG_T2_EAST_B1_O),
    .O(RMUX_T2_EAST_B1_O),
    .S(RMUX_T2_EAST_B1_sel_inst0_O)
);
RMUX_T2_EAST_B1_sel RMUX_T2_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_EAST_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T2_NORTH_B1 (
    .I_0(MUX_SB_T2_NORTH_SB_OUT_B1_O),
    .I_1(REG_T2_NORTH_B1_O),
    .O(RMUX_T2_NORTH_B1_O),
    .S(RMUX_T2_NORTH_B1_sel_inst0_O)
);
RMUX_T2_NORTH_B1_sel RMUX_T2_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_NORTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T2_SOUTH_B1 (
    .I_0(MUX_SB_T2_SOUTH_SB_OUT_B1_O),
    .I_1(REG_T2_SOUTH_B1_O),
    .O(RMUX_T2_SOUTH_B1_O),
    .S(RMUX_T2_SOUTH_B1_sel_inst0_O)
);
RMUX_T2_SOUTH_B1_sel RMUX_T2_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_SOUTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T2_WEST_B1 (
    .I_0(MUX_SB_T2_WEST_SB_OUT_B1_O),
    .I_1(REG_T2_WEST_B1_O),
    .O(RMUX_T2_WEST_B1_O),
    .S(RMUX_T2_WEST_B1_sel_inst0_O)
);
RMUX_T2_WEST_B1_sel RMUX_T2_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_WEST_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T3_EAST_B1 (
    .I_0(MUX_SB_T3_EAST_SB_OUT_B1_O),
    .I_1(REG_T3_EAST_B1_O),
    .O(RMUX_T3_EAST_B1_O),
    .S(RMUX_T3_EAST_B1_sel_inst0_O)
);
RMUX_T3_EAST_B1_sel RMUX_T3_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_EAST_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T3_NORTH_B1 (
    .I_0(MUX_SB_T3_NORTH_SB_OUT_B1_O),
    .I_1(REG_T3_NORTH_B1_O),
    .O(RMUX_T3_NORTH_B1_O),
    .S(RMUX_T3_NORTH_B1_sel_inst0_O)
);
RMUX_T3_NORTH_B1_sel RMUX_T3_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_NORTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T3_SOUTH_B1 (
    .I_0(MUX_SB_T3_SOUTH_SB_OUT_B1_O),
    .I_1(REG_T3_SOUTH_B1_O),
    .O(RMUX_T3_SOUTH_B1_O),
    .S(RMUX_T3_SOUTH_B1_sel_inst0_O)
);
RMUX_T3_SOUTH_B1_sel RMUX_T3_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_SOUTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T3_WEST_B1 (
    .I_0(MUX_SB_T3_WEST_SB_OUT_B1_O),
    .I_1(REG_T3_WEST_B1_O),
    .O(RMUX_T3_WEST_B1_O),
    .S(RMUX_T3_WEST_B1_sel_inst0_O)
);
RMUX_T3_WEST_B1_sel RMUX_T3_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_WEST_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T4_EAST_B1 (
    .I_0(MUX_SB_T4_EAST_SB_OUT_B1_O),
    .I_1(REG_T4_EAST_B1_O),
    .O(RMUX_T4_EAST_B1_O),
    .S(RMUX_T4_EAST_B1_sel_inst0_O)
);
RMUX_T4_EAST_B1_sel RMUX_T4_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_EAST_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T4_NORTH_B1 (
    .I_0(MUX_SB_T4_NORTH_SB_OUT_B1_O),
    .I_1(REG_T4_NORTH_B1_O),
    .O(RMUX_T4_NORTH_B1_O),
    .S(RMUX_T4_NORTH_B1_sel_inst0_O)
);
RMUX_T4_NORTH_B1_sel RMUX_T4_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_NORTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T4_SOUTH_B1 (
    .I_0(MUX_SB_T4_SOUTH_SB_OUT_B1_O),
    .I_1(REG_T4_SOUTH_B1_O),
    .O(RMUX_T4_SOUTH_B1_O),
    .S(RMUX_T4_SOUTH_B1_sel_inst0_O)
);
RMUX_T4_SOUTH_B1_sel RMUX_T4_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_SOUTH_B1_sel_inst0_O)
);
MuxWrapperAOIImpl_2_1 RMUX_T4_WEST_B1 (
    .I_0(MUX_SB_T4_WEST_SB_OUT_B1_O),
    .I_1(REG_T4_WEST_B1_O),
    .O(RMUX_T4_WEST_B1_O),
    .S(RMUX_T4_WEST_B1_sel_inst0_O)
);
RMUX_T4_WEST_B1_sel RMUX_T4_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_WEST_B1_sel_inst0_O)
);
SB_T0_EAST_SB_OUT_B1_sel SB_T0_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T0_NORTH_SB_OUT_B1_sel SB_T0_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T0_SOUTH_SB_OUT_B1_sel SB_T0_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T0_WEST_SB_OUT_B1_sel SB_T0_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_WEST_SB_OUT_B1_sel_inst0_O)
);
SB_T1_EAST_SB_OUT_B1_sel SB_T1_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T1_NORTH_SB_OUT_B1_sel SB_T1_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T1_SOUTH_SB_OUT_B1_sel SB_T1_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T1_WEST_SB_OUT_B1_sel SB_T1_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_WEST_SB_OUT_B1_sel_inst0_O)
);
SB_T2_EAST_SB_OUT_B1_sel SB_T2_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T2_NORTH_SB_OUT_B1_sel SB_T2_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T2_SOUTH_SB_OUT_B1_sel SB_T2_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T2_WEST_SB_OUT_B1_sel SB_T2_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_WEST_SB_OUT_B1_sel_inst0_O)
);
SB_T3_EAST_SB_OUT_B1_sel SB_T3_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T3_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T3_NORTH_SB_OUT_B1_sel SB_T3_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T3_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T3_SOUTH_SB_OUT_B1_sel SB_T3_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T3_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T3_WEST_SB_OUT_B1_sel SB_T3_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T3_WEST_SB_OUT_B1_sel_inst0_O)
);
SB_T4_EAST_SB_OUT_B1_sel SB_T4_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T4_NORTH_SB_OUT_B1_sel SB_T4_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T4_SOUTH_SB_OUT_B1_sel SB_T4_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T4_WEST_SB_OUT_B1_sel SB_T4_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_WEST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T0_EAST_SB_IN_B1 (
    .I(SB_T0_EAST_SB_IN_B1),
    .O(WIRE_SB_T0_EAST_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T0_NORTH_SB_IN_B1 (
    .I(SB_T0_NORTH_SB_IN_B1),
    .O(WIRE_SB_T0_NORTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T0_SOUTH_SB_IN_B1 (
    .I(SB_T0_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T0_WEST_SB_IN_B1 (
    .I(SB_T0_WEST_SB_IN_B1),
    .O(WIRE_SB_T0_WEST_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T1_EAST_SB_IN_B1 (
    .I(SB_T1_EAST_SB_IN_B1),
    .O(WIRE_SB_T1_EAST_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T1_NORTH_SB_IN_B1 (
    .I(SB_T1_NORTH_SB_IN_B1),
    .O(WIRE_SB_T1_NORTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T1_SOUTH_SB_IN_B1 (
    .I(SB_T1_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T1_WEST_SB_IN_B1 (
    .I(SB_T1_WEST_SB_IN_B1),
    .O(WIRE_SB_T1_WEST_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T2_EAST_SB_IN_B1 (
    .I(SB_T2_EAST_SB_IN_B1),
    .O(WIRE_SB_T2_EAST_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T2_NORTH_SB_IN_B1 (
    .I(SB_T2_NORTH_SB_IN_B1),
    .O(WIRE_SB_T2_NORTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T2_SOUTH_SB_IN_B1 (
    .I(SB_T2_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T2_WEST_SB_IN_B1 (
    .I(SB_T2_WEST_SB_IN_B1),
    .O(WIRE_SB_T2_WEST_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T3_EAST_SB_IN_B1 (
    .I(SB_T3_EAST_SB_IN_B1),
    .O(WIRE_SB_T3_EAST_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T3_NORTH_SB_IN_B1 (
    .I(SB_T3_NORTH_SB_IN_B1),
    .O(WIRE_SB_T3_NORTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T3_SOUTH_SB_IN_B1 (
    .I(SB_T3_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T3_WEST_SB_IN_B1 (
    .I(SB_T3_WEST_SB_IN_B1),
    .O(WIRE_SB_T3_WEST_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T4_EAST_SB_IN_B1 (
    .I(SB_T4_EAST_SB_IN_B1),
    .O(WIRE_SB_T4_EAST_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T4_NORTH_SB_IN_B1 (
    .I(SB_T4_NORTH_SB_IN_B1),
    .O(WIRE_SB_T4_NORTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T4_SOUTH_SB_IN_B1 (
    .I(SB_T4_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B1_O)
);
MuxWrapperAOI_1_1_Regular WIRE_SB_T4_WEST_SB_IN_B1 (
    .I(SB_T4_WEST_SB_IN_B1),
    .O(WIRE_SB_T4_WEST_SB_IN_B1_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_18_32_inst0$bit_const_0_None (
    .out(ZextWrapper_18_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_18_32_inst0$self_O_out;
assign ZextWrapper_18_32_inst0$self_O_out = {ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,config_reg_2_O};
mantle_wire__typeBitIn32 ZextWrapper_18_32_inst0$self_O (
    .in(ZextWrapper_18_32_inst0$self_O_in),
    .out(ZextWrapper_18_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_30_32_inst0$bit_const_0_None (
    .out(ZextWrapper_30_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_30_32_inst0$self_O_out;
assign ZextWrapper_30_32_inst0$self_O_out = {ZextWrapper_30_32_inst0$bit_const_0_None_out,ZextWrapper_30_32_inst0$bit_const_0_None_out,config_reg_1_O};
mantle_wire__typeBitIn32 ZextWrapper_30_32_inst0$self_O (
    .in(ZextWrapper_30_32_inst0$self_O_in),
    .out(ZextWrapper_30_32_inst0$self_O_out)
);
coreir_and #(
    .width(1)
) and1_inst0 (
    .in0(coreir_eq_1_inst0_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst0_out)
);
coreir_and #(
    .width(1)
) and1_inst1 (
    .in0(coreir_eq_1_inst1_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst1_out)
);
coreir_and #(
    .width(1)
) and1_inst10 (
    .in0(coreir_eq_1_inst10_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst10_out)
);
coreir_and #(
    .width(1)
) and1_inst11 (
    .in0(coreir_eq_1_inst11_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst11_out)
);
coreir_and #(
    .width(1)
) and1_inst12 (
    .in0(coreir_eq_1_inst12_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst12_out)
);
coreir_and #(
    .width(1)
) and1_inst13 (
    .in0(coreir_eq_1_inst13_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst13_out)
);
coreir_and #(
    .width(1)
) and1_inst14 (
    .in0(coreir_eq_1_inst14_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst14_out)
);
coreir_and #(
    .width(1)
) and1_inst15 (
    .in0(coreir_eq_1_inst15_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst15_out)
);
coreir_and #(
    .width(1)
) and1_inst16 (
    .in0(coreir_eq_1_inst16_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst16_out)
);
coreir_and #(
    .width(1)
) and1_inst17 (
    .in0(coreir_eq_1_inst17_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst17_out)
);
coreir_and #(
    .width(1)
) and1_inst18 (
    .in0(coreir_eq_1_inst18_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst18_out)
);
coreir_and #(
    .width(1)
) and1_inst19 (
    .in0(coreir_eq_1_inst19_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst19_out)
);
coreir_and #(
    .width(1)
) and1_inst2 (
    .in0(coreir_eq_1_inst2_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst2_out)
);
coreir_and #(
    .width(1)
) and1_inst3 (
    .in0(coreir_eq_1_inst3_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst3_out)
);
coreir_and #(
    .width(1)
) and1_inst4 (
    .in0(coreir_eq_1_inst4_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst4_out)
);
coreir_and #(
    .width(1)
) and1_inst5 (
    .in0(coreir_eq_1_inst5_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst5_out)
);
coreir_and #(
    .width(1)
) and1_inst6 (
    .in0(coreir_eq_1_inst6_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst6_out)
);
coreir_and #(
    .width(1)
) and1_inst7 (
    .in0(coreir_eq_1_inst7_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst7_out)
);
coreir_and #(
    .width(1)
) and1_inst8 (
    .in0(coreir_eq_1_inst8_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst8_out)
);
coreir_and #(
    .width(1)
) and1_inst9 (
    .in0(coreir_eq_1_inst9_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst9_out)
);
wire [7:0] config_reg_0_config_addr;
assign config_reg_0_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2],self_config_config_addr_out[1:0]};
ConfigRegister_32_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_reg_0_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_1_config_addr;
assign config_reg_1_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2],self_config_config_addr_out[1:0]};
ConfigRegister_30_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_reg_1_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_2_config_addr;
assign config_reg_2_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2],self_config_config_addr_out[1:0]};
ConfigRegister_18_8_32_2 config_reg_2 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_2_O),
    .config_addr(config_reg_2_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst0 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst0_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst1 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst10 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst10_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst11 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst11_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst12 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst12_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst13 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst13_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst14 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst14_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst15 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst15_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst16 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst16_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst17 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst17_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst18 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst18_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst19 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst19_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst2 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst2_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst3 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst3_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst4 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst4_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst5 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst5_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst6 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst6_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst7 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst7_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst8 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst8_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst9 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst9_out)
);
mantle_wire__typeBit8 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
assign SB_T0_EAST_SB_OUT_B1 = RMUX_T0_EAST_B1_O;
assign SB_T0_NORTH_SB_OUT_B1 = RMUX_T0_NORTH_B1_O;
assign SB_T0_SOUTH_SB_OUT_B1 = RMUX_T0_SOUTH_B1_O;
assign SB_T0_WEST_SB_OUT_B1 = RMUX_T0_WEST_B1_O;
assign SB_T1_EAST_SB_OUT_B1 = RMUX_T1_EAST_B1_O;
assign SB_T1_NORTH_SB_OUT_B1 = RMUX_T1_NORTH_B1_O;
assign SB_T1_SOUTH_SB_OUT_B1 = RMUX_T1_SOUTH_B1_O;
assign SB_T1_WEST_SB_OUT_B1 = RMUX_T1_WEST_B1_O;
assign SB_T2_EAST_SB_OUT_B1 = RMUX_T2_EAST_B1_O;
assign SB_T2_NORTH_SB_OUT_B1 = RMUX_T2_NORTH_B1_O;
assign SB_T2_SOUTH_SB_OUT_B1 = RMUX_T2_SOUTH_B1_O;
assign SB_T2_WEST_SB_OUT_B1 = RMUX_T2_WEST_B1_O;
assign SB_T3_EAST_SB_OUT_B1 = RMUX_T3_EAST_B1_O;
assign SB_T3_NORTH_SB_OUT_B1 = RMUX_T3_NORTH_B1_O;
assign SB_T3_SOUTH_SB_OUT_B1 = RMUX_T3_SOUTH_B1_O;
assign SB_T3_WEST_SB_OUT_B1 = RMUX_T3_WEST_B1_O;
assign SB_T4_EAST_SB_OUT_B1 = RMUX_T4_EAST_B1_O;
assign SB_T4_NORTH_SB_OUT_B1 = RMUX_T4_NORTH_B1_O;
assign SB_T4_SOUTH_SB_OUT_B1 = RMUX_T4_SOUTH_B1_O;
assign SB_T4_WEST_SB_OUT_B1 = RMUX_T4_WEST_B1_O;
assign read_config_data = MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0_out;
endmodule

module SB_ID0_5TRACKS_B16_PE (
    input [15:0] SB_T0_EAST_SB_IN_B16,
    output [15:0] SB_T0_EAST_SB_OUT_B16,
    input [15:0] SB_T0_NORTH_SB_IN_B16,
    output [15:0] SB_T0_NORTH_SB_OUT_B16,
    input [15:0] SB_T0_SOUTH_SB_IN_B16,
    output [15:0] SB_T0_SOUTH_SB_OUT_B16,
    input [15:0] SB_T0_WEST_SB_IN_B16,
    output [15:0] SB_T0_WEST_SB_OUT_B16,
    input [15:0] SB_T1_EAST_SB_IN_B16,
    output [15:0] SB_T1_EAST_SB_OUT_B16,
    input [15:0] SB_T1_NORTH_SB_IN_B16,
    output [15:0] SB_T1_NORTH_SB_OUT_B16,
    input [15:0] SB_T1_SOUTH_SB_IN_B16,
    output [15:0] SB_T1_SOUTH_SB_OUT_B16,
    input [15:0] SB_T1_WEST_SB_IN_B16,
    output [15:0] SB_T1_WEST_SB_OUT_B16,
    input [15:0] SB_T2_EAST_SB_IN_B16,
    output [15:0] SB_T2_EAST_SB_OUT_B16,
    input [15:0] SB_T2_NORTH_SB_IN_B16,
    output [15:0] SB_T2_NORTH_SB_OUT_B16,
    input [15:0] SB_T2_SOUTH_SB_IN_B16,
    output [15:0] SB_T2_SOUTH_SB_OUT_B16,
    input [15:0] SB_T2_WEST_SB_IN_B16,
    output [15:0] SB_T2_WEST_SB_OUT_B16,
    input [15:0] SB_T3_EAST_SB_IN_B16,
    output [15:0] SB_T3_EAST_SB_OUT_B16,
    input [15:0] SB_T3_NORTH_SB_IN_B16,
    output [15:0] SB_T3_NORTH_SB_OUT_B16,
    input [15:0] SB_T3_SOUTH_SB_IN_B16,
    output [15:0] SB_T3_SOUTH_SB_OUT_B16,
    input [15:0] SB_T3_WEST_SB_IN_B16,
    output [15:0] SB_T3_WEST_SB_OUT_B16,
    input [15:0] SB_T4_EAST_SB_IN_B16,
    output [15:0] SB_T4_EAST_SB_OUT_B16,
    input [15:0] SB_T4_NORTH_SB_IN_B16,
    output [15:0] SB_T4_NORTH_SB_OUT_B16,
    input [15:0] SB_T4_SOUTH_SB_IN_B16,
    output [15:0] SB_T4_SOUTH_SB_OUT_B16,
    input [15:0] SB_T4_WEST_SB_IN_B16,
    output [15:0] SB_T4_WEST_SB_OUT_B16,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    input [15:0] data_out_pond,
    input [15:0] pe_outputs_0,
    output [31:0] read_config_data,
    input reset,
    input [0:0] stall
);
wire [0:0] Invert1_inst0_out;
wire [15:0] MUX_SB_T0_EAST_SB_OUT_B16_O;
wire [15:0] MUX_SB_T0_NORTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T0_SOUTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T0_WEST_SB_OUT_B16_O;
wire [15:0] MUX_SB_T1_EAST_SB_OUT_B16_O;
wire [15:0] MUX_SB_T1_NORTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T1_SOUTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T1_WEST_SB_OUT_B16_O;
wire [15:0] MUX_SB_T2_EAST_SB_OUT_B16_O;
wire [15:0] MUX_SB_T2_NORTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T2_SOUTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T2_WEST_SB_OUT_B16_O;
wire [15:0] MUX_SB_T3_EAST_SB_OUT_B16_O;
wire [15:0] MUX_SB_T3_NORTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T3_SOUTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T3_WEST_SB_OUT_B16_O;
wire [15:0] MUX_SB_T4_EAST_SB_OUT_B16_O;
wire [15:0] MUX_SB_T4_NORTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T4_SOUTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T4_WEST_SB_OUT_B16_O;
wire [31:0] MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0_out;
wire [15:0] REG_T0_EAST_B16_O;
wire [15:0] REG_T0_NORTH_B16_O;
wire [15:0] REG_T0_SOUTH_B16_O;
wire [15:0] REG_T0_WEST_B16_O;
wire [15:0] REG_T1_EAST_B16_O;
wire [15:0] REG_T1_NORTH_B16_O;
wire [15:0] REG_T1_SOUTH_B16_O;
wire [15:0] REG_T1_WEST_B16_O;
wire [15:0] REG_T2_EAST_B16_O;
wire [15:0] REG_T2_NORTH_B16_O;
wire [15:0] REG_T2_SOUTH_B16_O;
wire [15:0] REG_T2_WEST_B16_O;
wire [15:0] REG_T3_EAST_B16_O;
wire [15:0] REG_T3_NORTH_B16_O;
wire [15:0] REG_T3_SOUTH_B16_O;
wire [15:0] REG_T3_WEST_B16_O;
wire [15:0] REG_T4_EAST_B16_O;
wire [15:0] REG_T4_NORTH_B16_O;
wire [15:0] REG_T4_SOUTH_B16_O;
wire [15:0] REG_T4_WEST_B16_O;
wire [15:0] RMUX_T0_EAST_B16_O;
wire [0:0] RMUX_T0_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T0_NORTH_B16_O;
wire [0:0] RMUX_T0_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T0_SOUTH_B16_O;
wire [0:0] RMUX_T0_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T0_WEST_B16_O;
wire [0:0] RMUX_T0_WEST_B16_sel_inst0_O;
wire [15:0] RMUX_T1_EAST_B16_O;
wire [0:0] RMUX_T1_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T1_NORTH_B16_O;
wire [0:0] RMUX_T1_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T1_SOUTH_B16_O;
wire [0:0] RMUX_T1_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T1_WEST_B16_O;
wire [0:0] RMUX_T1_WEST_B16_sel_inst0_O;
wire [15:0] RMUX_T2_EAST_B16_O;
wire [0:0] RMUX_T2_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T2_NORTH_B16_O;
wire [0:0] RMUX_T2_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T2_SOUTH_B16_O;
wire [0:0] RMUX_T2_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T2_WEST_B16_O;
wire [0:0] RMUX_T2_WEST_B16_sel_inst0_O;
wire [15:0] RMUX_T3_EAST_B16_O;
wire [0:0] RMUX_T3_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T3_NORTH_B16_O;
wire [0:0] RMUX_T3_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T3_SOUTH_B16_O;
wire [0:0] RMUX_T3_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T3_WEST_B16_O;
wire [0:0] RMUX_T3_WEST_B16_sel_inst0_O;
wire [15:0] RMUX_T4_EAST_B16_O;
wire [0:0] RMUX_T4_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T4_NORTH_B16_O;
wire [0:0] RMUX_T4_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T4_SOUTH_B16_O;
wire [0:0] RMUX_T4_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T4_WEST_B16_O;
wire [0:0] RMUX_T4_WEST_B16_sel_inst0_O;
wire [2:0] SB_T0_EAST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T0_NORTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T0_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T0_WEST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T1_EAST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T1_NORTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T1_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T1_WEST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T2_EAST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T2_NORTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T2_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T2_WEST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T3_EAST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T3_NORTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T3_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T3_WEST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T4_EAST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T4_NORTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T4_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T4_WEST_SB_OUT_B16_sel_inst0_O;
wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T3_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T3_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T3_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T3_WEST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T4_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T4_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T4_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T4_WEST_SB_IN_B16_O;
wire ZextWrapper_18_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_18_32_inst0$self_O_in;
wire ZextWrapper_30_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_30_32_inst0$self_O_in;
wire [0:0] and1_inst0_out;
wire [0:0] and1_inst1_out;
wire [0:0] and1_inst10_out;
wire [0:0] and1_inst11_out;
wire [0:0] and1_inst12_out;
wire [0:0] and1_inst13_out;
wire [0:0] and1_inst14_out;
wire [0:0] and1_inst15_out;
wire [0:0] and1_inst16_out;
wire [0:0] and1_inst17_out;
wire [0:0] and1_inst18_out;
wire [0:0] and1_inst19_out;
wire [0:0] and1_inst2_out;
wire [0:0] and1_inst3_out;
wire [0:0] and1_inst4_out;
wire [0:0] and1_inst5_out;
wire [0:0] and1_inst6_out;
wire [0:0] and1_inst7_out;
wire [0:0] and1_inst8_out;
wire [0:0] and1_inst9_out;
wire [31:0] config_reg_0_O;
wire [29:0] config_reg_1_O;
wire [17:0] config_reg_2_O;
wire [0:0] const_1_1_out;
wire coreir_eq_1_inst0_out;
wire coreir_eq_1_inst1_out;
wire coreir_eq_1_inst10_out;
wire coreir_eq_1_inst11_out;
wire coreir_eq_1_inst12_out;
wire coreir_eq_1_inst13_out;
wire coreir_eq_1_inst14_out;
wire coreir_eq_1_inst15_out;
wire coreir_eq_1_inst16_out;
wire coreir_eq_1_inst17_out;
wire coreir_eq_1_inst18_out;
wire coreir_eq_1_inst19_out;
wire coreir_eq_1_inst2_out;
wire coreir_eq_1_inst3_out;
wire coreir_eq_1_inst4_out;
wire coreir_eq_1_inst5_out;
wire coreir_eq_1_inst6_out;
wire coreir_eq_1_inst7_out;
wire coreir_eq_1_inst8_out;
wire coreir_eq_1_inst9_out;
wire [7:0] self_config_config_addr_out;
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(stall),
    .out(Invert1_inst0_out)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T0_EAST_SB_OUT_B16 (
    .I_0(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_1(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T0_EAST_SB_OUT_B16_O),
    .S(SB_T0_EAST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T0_NORTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_1(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T0_NORTH_SB_OUT_B16_O),
    .S(SB_T0_NORTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T0_SOUTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T0_SOUTH_SB_OUT_B16_O),
    .S(SB_T0_SOUTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T0_WEST_SB_OUT_B16 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T0_WEST_SB_OUT_B16_O),
    .S(SB_T0_WEST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T1_EAST_SB_OUT_B16 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T1_EAST_SB_OUT_B16_O),
    .S(SB_T1_EAST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T1_NORTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_1(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T1_NORTH_SB_OUT_B16_O),
    .S(SB_T1_NORTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T1_SOUTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_1(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T1_SOUTH_SB_OUT_B16_O),
    .S(SB_T1_SOUTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T1_WEST_SB_OUT_B16 (
    .I_0(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T1_WEST_SB_OUT_B16_O),
    .S(SB_T1_WEST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T2_EAST_SB_OUT_B16 (
    .I_0(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T2_EAST_SB_OUT_B16_O),
    .S(SB_T2_EAST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T2_NORTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_1(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T2_NORTH_SB_OUT_B16_O),
    .S(SB_T2_NORTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T2_SOUTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_1(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T2_SOUTH_SB_OUT_B16_O),
    .S(SB_T2_SOUTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T2_WEST_SB_OUT_B16 (
    .I_0(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T2_WEST_SB_OUT_B16_O),
    .S(SB_T2_WEST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T3_EAST_SB_OUT_B16 (
    .I_0(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T3_EAST_SB_OUT_B16_O),
    .S(SB_T3_EAST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T3_NORTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_1(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_2(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T3_NORTH_SB_OUT_B16_O),
    .S(SB_T3_NORTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T3_SOUTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_1(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T3_SOUTH_SB_OUT_B16_O),
    .S(SB_T3_SOUTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T3_WEST_SB_OUT_B16 (
    .I_0(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T3_WEST_SB_OUT_B16_O),
    .S(SB_T3_WEST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T4_EAST_SB_OUT_B16 (
    .I_0(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T4_EAST_SB_OUT_B16_O),
    .S(SB_T4_EAST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T4_NORTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_2(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T4_NORTH_SB_OUT_B16_O),
    .S(SB_T4_NORTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T4_SOUTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_1(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_2(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T4_SOUTH_SB_OUT_B16_O),
    .S(SB_T4_SOUTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T4_WEST_SB_OUT_B16 (
    .I_0(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_3(data_out_pond),
    .I_4(pe_outputs_0),
    .O(MUX_SB_T4_WEST_SB_OUT_B16_O),
    .S(SB_T4_WEST_SB_OUT_B16_sel_inst0_O)
);
commonlib_muxn__N3__width32 MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0 (
    .in_data_0(config_reg_0_O),
    .in_data_1(ZextWrapper_30_32_inst0$self_O_in),
    .in_data_2(ZextWrapper_18_32_inst0$self_O_in),
    .in_sel(self_config_config_addr_out[1:0]),
    .out(MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0_out)
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_EAST_B16 (
    .I(MUX_SB_T0_EAST_SB_OUT_B16_O),
    .O(REG_T0_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst2_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_NORTH_B16 (
    .I(MUX_SB_T0_NORTH_SB_OUT_B16_O),
    .O(REG_T0_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst0_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_SOUTH_B16 (
    .I(MUX_SB_T0_SOUTH_SB_OUT_B16_O),
    .O(REG_T0_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst1_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_WEST_B16 (
    .I(MUX_SB_T0_WEST_SB_OUT_B16_O),
    .O(REG_T0_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst3_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_EAST_B16 (
    .I(MUX_SB_T1_EAST_SB_OUT_B16_O),
    .O(REG_T1_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst6_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_NORTH_B16 (
    .I(MUX_SB_T1_NORTH_SB_OUT_B16_O),
    .O(REG_T1_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst4_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_SOUTH_B16 (
    .I(MUX_SB_T1_SOUTH_SB_OUT_B16_O),
    .O(REG_T1_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst5_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_WEST_B16 (
    .I(MUX_SB_T1_WEST_SB_OUT_B16_O),
    .O(REG_T1_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst7_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_EAST_B16 (
    .I(MUX_SB_T2_EAST_SB_OUT_B16_O),
    .O(REG_T2_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst10_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_NORTH_B16 (
    .I(MUX_SB_T2_NORTH_SB_OUT_B16_O),
    .O(REG_T2_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst8_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_SOUTH_B16 (
    .I(MUX_SB_T2_SOUTH_SB_OUT_B16_O),
    .O(REG_T2_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst9_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_WEST_B16 (
    .I(MUX_SB_T2_WEST_SB_OUT_B16_O),
    .O(REG_T2_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst11_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T3_EAST_B16 (
    .I(MUX_SB_T3_EAST_SB_OUT_B16_O),
    .O(REG_T3_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst14_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T3_NORTH_B16 (
    .I(MUX_SB_T3_NORTH_SB_OUT_B16_O),
    .O(REG_T3_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst12_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T3_SOUTH_B16 (
    .I(MUX_SB_T3_SOUTH_SB_OUT_B16_O),
    .O(REG_T3_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst13_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T3_WEST_B16 (
    .I(MUX_SB_T3_WEST_SB_OUT_B16_O),
    .O(REG_T3_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst15_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T4_EAST_B16 (
    .I(MUX_SB_T4_EAST_SB_OUT_B16_O),
    .O(REG_T4_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst18_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T4_NORTH_B16 (
    .I(MUX_SB_T4_NORTH_SB_OUT_B16_O),
    .O(REG_T4_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst16_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T4_SOUTH_B16 (
    .I(MUX_SB_T4_SOUTH_SB_OUT_B16_O),
    .O(REG_T4_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst17_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T4_WEST_B16 (
    .I(MUX_SB_T4_WEST_SB_OUT_B16_O),
    .O(REG_T4_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst19_out[0])
);
MuxWrapperAOIImpl_2_16 RMUX_T0_EAST_B16 (
    .I_0(MUX_SB_T0_EAST_SB_OUT_B16_O),
    .I_1(REG_T0_EAST_B16_O),
    .O(RMUX_T0_EAST_B16_O),
    .S(RMUX_T0_EAST_B16_sel_inst0_O)
);
RMUX_T0_EAST_B16_sel RMUX_T0_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_EAST_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T0_NORTH_B16 (
    .I_0(MUX_SB_T0_NORTH_SB_OUT_B16_O),
    .I_1(REG_T0_NORTH_B16_O),
    .O(RMUX_T0_NORTH_B16_O),
    .S(RMUX_T0_NORTH_B16_sel_inst0_O)
);
RMUX_T0_NORTH_B16_sel RMUX_T0_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_NORTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T0_SOUTH_B16 (
    .I_0(MUX_SB_T0_SOUTH_SB_OUT_B16_O),
    .I_1(REG_T0_SOUTH_B16_O),
    .O(RMUX_T0_SOUTH_B16_O),
    .S(RMUX_T0_SOUTH_B16_sel_inst0_O)
);
RMUX_T0_SOUTH_B16_sel RMUX_T0_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_SOUTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T0_WEST_B16 (
    .I_0(MUX_SB_T0_WEST_SB_OUT_B16_O),
    .I_1(REG_T0_WEST_B16_O),
    .O(RMUX_T0_WEST_B16_O),
    .S(RMUX_T0_WEST_B16_sel_inst0_O)
);
RMUX_T0_WEST_B16_sel RMUX_T0_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_WEST_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T1_EAST_B16 (
    .I_0(MUX_SB_T1_EAST_SB_OUT_B16_O),
    .I_1(REG_T1_EAST_B16_O),
    .O(RMUX_T1_EAST_B16_O),
    .S(RMUX_T1_EAST_B16_sel_inst0_O)
);
RMUX_T1_EAST_B16_sel RMUX_T1_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_EAST_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T1_NORTH_B16 (
    .I_0(MUX_SB_T1_NORTH_SB_OUT_B16_O),
    .I_1(REG_T1_NORTH_B16_O),
    .O(RMUX_T1_NORTH_B16_O),
    .S(RMUX_T1_NORTH_B16_sel_inst0_O)
);
RMUX_T1_NORTH_B16_sel RMUX_T1_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_NORTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T1_SOUTH_B16 (
    .I_0(MUX_SB_T1_SOUTH_SB_OUT_B16_O),
    .I_1(REG_T1_SOUTH_B16_O),
    .O(RMUX_T1_SOUTH_B16_O),
    .S(RMUX_T1_SOUTH_B16_sel_inst0_O)
);
RMUX_T1_SOUTH_B16_sel RMUX_T1_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_SOUTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T1_WEST_B16 (
    .I_0(MUX_SB_T1_WEST_SB_OUT_B16_O),
    .I_1(REG_T1_WEST_B16_O),
    .O(RMUX_T1_WEST_B16_O),
    .S(RMUX_T1_WEST_B16_sel_inst0_O)
);
RMUX_T1_WEST_B16_sel RMUX_T1_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_WEST_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T2_EAST_B16 (
    .I_0(MUX_SB_T2_EAST_SB_OUT_B16_O),
    .I_1(REG_T2_EAST_B16_O),
    .O(RMUX_T2_EAST_B16_O),
    .S(RMUX_T2_EAST_B16_sel_inst0_O)
);
RMUX_T2_EAST_B16_sel RMUX_T2_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_EAST_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T2_NORTH_B16 (
    .I_0(MUX_SB_T2_NORTH_SB_OUT_B16_O),
    .I_1(REG_T2_NORTH_B16_O),
    .O(RMUX_T2_NORTH_B16_O),
    .S(RMUX_T2_NORTH_B16_sel_inst0_O)
);
RMUX_T2_NORTH_B16_sel RMUX_T2_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_NORTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T2_SOUTH_B16 (
    .I_0(MUX_SB_T2_SOUTH_SB_OUT_B16_O),
    .I_1(REG_T2_SOUTH_B16_O),
    .O(RMUX_T2_SOUTH_B16_O),
    .S(RMUX_T2_SOUTH_B16_sel_inst0_O)
);
RMUX_T2_SOUTH_B16_sel RMUX_T2_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_SOUTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T2_WEST_B16 (
    .I_0(MUX_SB_T2_WEST_SB_OUT_B16_O),
    .I_1(REG_T2_WEST_B16_O),
    .O(RMUX_T2_WEST_B16_O),
    .S(RMUX_T2_WEST_B16_sel_inst0_O)
);
RMUX_T2_WEST_B16_sel RMUX_T2_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_WEST_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T3_EAST_B16 (
    .I_0(MUX_SB_T3_EAST_SB_OUT_B16_O),
    .I_1(REG_T3_EAST_B16_O),
    .O(RMUX_T3_EAST_B16_O),
    .S(RMUX_T3_EAST_B16_sel_inst0_O)
);
RMUX_T3_EAST_B16_sel RMUX_T3_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_EAST_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T3_NORTH_B16 (
    .I_0(MUX_SB_T3_NORTH_SB_OUT_B16_O),
    .I_1(REG_T3_NORTH_B16_O),
    .O(RMUX_T3_NORTH_B16_O),
    .S(RMUX_T3_NORTH_B16_sel_inst0_O)
);
RMUX_T3_NORTH_B16_sel RMUX_T3_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_NORTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T3_SOUTH_B16 (
    .I_0(MUX_SB_T3_SOUTH_SB_OUT_B16_O),
    .I_1(REG_T3_SOUTH_B16_O),
    .O(RMUX_T3_SOUTH_B16_O),
    .S(RMUX_T3_SOUTH_B16_sel_inst0_O)
);
RMUX_T3_SOUTH_B16_sel RMUX_T3_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_SOUTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T3_WEST_B16 (
    .I_0(MUX_SB_T3_WEST_SB_OUT_B16_O),
    .I_1(REG_T3_WEST_B16_O),
    .O(RMUX_T3_WEST_B16_O),
    .S(RMUX_T3_WEST_B16_sel_inst0_O)
);
RMUX_T3_WEST_B16_sel RMUX_T3_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_WEST_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T4_EAST_B16 (
    .I_0(MUX_SB_T4_EAST_SB_OUT_B16_O),
    .I_1(REG_T4_EAST_B16_O),
    .O(RMUX_T4_EAST_B16_O),
    .S(RMUX_T4_EAST_B16_sel_inst0_O)
);
RMUX_T4_EAST_B16_sel RMUX_T4_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_EAST_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T4_NORTH_B16 (
    .I_0(MUX_SB_T4_NORTH_SB_OUT_B16_O),
    .I_1(REG_T4_NORTH_B16_O),
    .O(RMUX_T4_NORTH_B16_O),
    .S(RMUX_T4_NORTH_B16_sel_inst0_O)
);
RMUX_T4_NORTH_B16_sel RMUX_T4_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_NORTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T4_SOUTH_B16 (
    .I_0(MUX_SB_T4_SOUTH_SB_OUT_B16_O),
    .I_1(REG_T4_SOUTH_B16_O),
    .O(RMUX_T4_SOUTH_B16_O),
    .S(RMUX_T4_SOUTH_B16_sel_inst0_O)
);
RMUX_T4_SOUTH_B16_sel RMUX_T4_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_SOUTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T4_WEST_B16 (
    .I_0(MUX_SB_T4_WEST_SB_OUT_B16_O),
    .I_1(REG_T4_WEST_B16_O),
    .O(RMUX_T4_WEST_B16_O),
    .S(RMUX_T4_WEST_B16_sel_inst0_O)
);
RMUX_T4_WEST_B16_sel RMUX_T4_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_WEST_B16_sel_inst0_O)
);
SB_T0_EAST_SB_OUT_B16_sel SB_T0_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T0_NORTH_SB_OUT_B16_sel SB_T0_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T0_SOUTH_SB_OUT_B16_sel SB_T0_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T0_WEST_SB_OUT_B16_sel SB_T0_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_WEST_SB_OUT_B16_sel_inst0_O)
);
SB_T1_EAST_SB_OUT_B16_sel SB_T1_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T1_NORTH_SB_OUT_B16_sel SB_T1_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T1_SOUTH_SB_OUT_B16_sel SB_T1_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T1_WEST_SB_OUT_B16_sel SB_T1_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_WEST_SB_OUT_B16_sel_inst0_O)
);
SB_T2_EAST_SB_OUT_B16_sel SB_T2_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T2_NORTH_SB_OUT_B16_sel SB_T2_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T2_SOUTH_SB_OUT_B16_sel SB_T2_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T2_WEST_SB_OUT_B16_sel SB_T2_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_WEST_SB_OUT_B16_sel_inst0_O)
);
SB_T3_EAST_SB_OUT_B16_sel SB_T3_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T3_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T3_NORTH_SB_OUT_B16_sel SB_T3_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T3_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T3_SOUTH_SB_OUT_B16_sel SB_T3_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T3_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T3_WEST_SB_OUT_B16_sel SB_T3_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T3_WEST_SB_OUT_B16_sel_inst0_O)
);
SB_T4_EAST_SB_OUT_B16_sel SB_T4_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T4_NORTH_SB_OUT_B16_sel SB_T4_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T4_SOUTH_SB_OUT_B16_sel SB_T4_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T4_WEST_SB_OUT_B16_sel SB_T4_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_WEST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T0_EAST_SB_IN_B16 (
    .I(SB_T0_EAST_SB_IN_B16),
    .O(WIRE_SB_T0_EAST_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T0_NORTH_SB_IN_B16 (
    .I(SB_T0_NORTH_SB_IN_B16),
    .O(WIRE_SB_T0_NORTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T0_SOUTH_SB_IN_B16 (
    .I(SB_T0_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T0_WEST_SB_IN_B16 (
    .I(SB_T0_WEST_SB_IN_B16),
    .O(WIRE_SB_T0_WEST_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T1_EAST_SB_IN_B16 (
    .I(SB_T1_EAST_SB_IN_B16),
    .O(WIRE_SB_T1_EAST_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T1_NORTH_SB_IN_B16 (
    .I(SB_T1_NORTH_SB_IN_B16),
    .O(WIRE_SB_T1_NORTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T1_SOUTH_SB_IN_B16 (
    .I(SB_T1_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T1_WEST_SB_IN_B16 (
    .I(SB_T1_WEST_SB_IN_B16),
    .O(WIRE_SB_T1_WEST_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T2_EAST_SB_IN_B16 (
    .I(SB_T2_EAST_SB_IN_B16),
    .O(WIRE_SB_T2_EAST_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T2_NORTH_SB_IN_B16 (
    .I(SB_T2_NORTH_SB_IN_B16),
    .O(WIRE_SB_T2_NORTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T2_SOUTH_SB_IN_B16 (
    .I(SB_T2_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T2_WEST_SB_IN_B16 (
    .I(SB_T2_WEST_SB_IN_B16),
    .O(WIRE_SB_T2_WEST_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T3_EAST_SB_IN_B16 (
    .I(SB_T3_EAST_SB_IN_B16),
    .O(WIRE_SB_T3_EAST_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T3_NORTH_SB_IN_B16 (
    .I(SB_T3_NORTH_SB_IN_B16),
    .O(WIRE_SB_T3_NORTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T3_SOUTH_SB_IN_B16 (
    .I(SB_T3_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T3_WEST_SB_IN_B16 (
    .I(SB_T3_WEST_SB_IN_B16),
    .O(WIRE_SB_T3_WEST_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T4_EAST_SB_IN_B16 (
    .I(SB_T4_EAST_SB_IN_B16),
    .O(WIRE_SB_T4_EAST_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T4_NORTH_SB_IN_B16 (
    .I(SB_T4_NORTH_SB_IN_B16),
    .O(WIRE_SB_T4_NORTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T4_SOUTH_SB_IN_B16 (
    .I(SB_T4_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T4_WEST_SB_IN_B16 (
    .I(SB_T4_WEST_SB_IN_B16),
    .O(WIRE_SB_T4_WEST_SB_IN_B16_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_18_32_inst0$bit_const_0_None (
    .out(ZextWrapper_18_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_18_32_inst0$self_O_out;
assign ZextWrapper_18_32_inst0$self_O_out = {ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,config_reg_2_O};
mantle_wire__typeBitIn32 ZextWrapper_18_32_inst0$self_O (
    .in(ZextWrapper_18_32_inst0$self_O_in),
    .out(ZextWrapper_18_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_30_32_inst0$bit_const_0_None (
    .out(ZextWrapper_30_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_30_32_inst0$self_O_out;
assign ZextWrapper_30_32_inst0$self_O_out = {ZextWrapper_30_32_inst0$bit_const_0_None_out,ZextWrapper_30_32_inst0$bit_const_0_None_out,config_reg_1_O};
mantle_wire__typeBitIn32 ZextWrapper_30_32_inst0$self_O (
    .in(ZextWrapper_30_32_inst0$self_O_in),
    .out(ZextWrapper_30_32_inst0$self_O_out)
);
coreir_and #(
    .width(1)
) and1_inst0 (
    .in0(coreir_eq_1_inst0_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst0_out)
);
coreir_and #(
    .width(1)
) and1_inst1 (
    .in0(coreir_eq_1_inst1_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst1_out)
);
coreir_and #(
    .width(1)
) and1_inst10 (
    .in0(coreir_eq_1_inst10_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst10_out)
);
coreir_and #(
    .width(1)
) and1_inst11 (
    .in0(coreir_eq_1_inst11_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst11_out)
);
coreir_and #(
    .width(1)
) and1_inst12 (
    .in0(coreir_eq_1_inst12_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst12_out)
);
coreir_and #(
    .width(1)
) and1_inst13 (
    .in0(coreir_eq_1_inst13_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst13_out)
);
coreir_and #(
    .width(1)
) and1_inst14 (
    .in0(coreir_eq_1_inst14_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst14_out)
);
coreir_and #(
    .width(1)
) and1_inst15 (
    .in0(coreir_eq_1_inst15_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst15_out)
);
coreir_and #(
    .width(1)
) and1_inst16 (
    .in0(coreir_eq_1_inst16_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst16_out)
);
coreir_and #(
    .width(1)
) and1_inst17 (
    .in0(coreir_eq_1_inst17_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst17_out)
);
coreir_and #(
    .width(1)
) and1_inst18 (
    .in0(coreir_eq_1_inst18_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst18_out)
);
coreir_and #(
    .width(1)
) and1_inst19 (
    .in0(coreir_eq_1_inst19_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst19_out)
);
coreir_and #(
    .width(1)
) and1_inst2 (
    .in0(coreir_eq_1_inst2_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst2_out)
);
coreir_and #(
    .width(1)
) and1_inst3 (
    .in0(coreir_eq_1_inst3_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst3_out)
);
coreir_and #(
    .width(1)
) and1_inst4 (
    .in0(coreir_eq_1_inst4_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst4_out)
);
coreir_and #(
    .width(1)
) and1_inst5 (
    .in0(coreir_eq_1_inst5_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst5_out)
);
coreir_and #(
    .width(1)
) and1_inst6 (
    .in0(coreir_eq_1_inst6_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst6_out)
);
coreir_and #(
    .width(1)
) and1_inst7 (
    .in0(coreir_eq_1_inst7_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst7_out)
);
coreir_and #(
    .width(1)
) and1_inst8 (
    .in0(coreir_eq_1_inst8_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst8_out)
);
coreir_and #(
    .width(1)
) and1_inst9 (
    .in0(coreir_eq_1_inst9_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst9_out)
);
wire [7:0] config_reg_0_config_addr;
assign config_reg_0_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2],self_config_config_addr_out[1:0]};
ConfigRegister_32_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_reg_0_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_1_config_addr;
assign config_reg_1_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2],self_config_config_addr_out[1:0]};
ConfigRegister_30_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_reg_1_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_2_config_addr;
assign config_reg_2_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2],self_config_config_addr_out[1:0]};
ConfigRegister_18_8_32_2 config_reg_2 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_2_O),
    .config_addr(config_reg_2_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst0 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst0_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst1 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst10 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst10_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst11 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst11_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst12 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst12_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst13 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst13_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst14 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst14_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst15 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst15_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst16 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst16_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst17 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst17_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst18 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst18_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst19 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst19_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst2 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst2_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst3 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst3_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst4 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst4_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst5 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst5_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst6 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst6_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst7 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst7_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst8 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst8_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst9 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst9_out)
);
mantle_wire__typeBit8 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
assign SB_T0_EAST_SB_OUT_B16 = RMUX_T0_EAST_B16_O;
assign SB_T0_NORTH_SB_OUT_B16 = RMUX_T0_NORTH_B16_O;
assign SB_T0_SOUTH_SB_OUT_B16 = RMUX_T0_SOUTH_B16_O;
assign SB_T0_WEST_SB_OUT_B16 = RMUX_T0_WEST_B16_O;
assign SB_T1_EAST_SB_OUT_B16 = RMUX_T1_EAST_B16_O;
assign SB_T1_NORTH_SB_OUT_B16 = RMUX_T1_NORTH_B16_O;
assign SB_T1_SOUTH_SB_OUT_B16 = RMUX_T1_SOUTH_B16_O;
assign SB_T1_WEST_SB_OUT_B16 = RMUX_T1_WEST_B16_O;
assign SB_T2_EAST_SB_OUT_B16 = RMUX_T2_EAST_B16_O;
assign SB_T2_NORTH_SB_OUT_B16 = RMUX_T2_NORTH_B16_O;
assign SB_T2_SOUTH_SB_OUT_B16 = RMUX_T2_SOUTH_B16_O;
assign SB_T2_WEST_SB_OUT_B16 = RMUX_T2_WEST_B16_O;
assign SB_T3_EAST_SB_OUT_B16 = RMUX_T3_EAST_B16_O;
assign SB_T3_NORTH_SB_OUT_B16 = RMUX_T3_NORTH_B16_O;
assign SB_T3_SOUTH_SB_OUT_B16 = RMUX_T3_SOUTH_B16_O;
assign SB_T3_WEST_SB_OUT_B16 = RMUX_T3_WEST_B16_O;
assign SB_T4_EAST_SB_OUT_B16 = RMUX_T4_EAST_B16_O;
assign SB_T4_NORTH_SB_OUT_B16 = RMUX_T4_NORTH_B16_O;
assign SB_T4_SOUTH_SB_OUT_B16 = RMUX_T4_SOUTH_B16_O;
assign SB_T4_WEST_SB_OUT_B16 = RMUX_T4_WEST_B16_O;
assign read_config_data = MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0_out;
endmodule

module SB_ID0_5TRACKS_B16_MemCore (
    input [15:0] SB_T0_EAST_SB_IN_B16,
    output [15:0] SB_T0_EAST_SB_OUT_B16,
    input [15:0] SB_T0_NORTH_SB_IN_B16,
    output [15:0] SB_T0_NORTH_SB_OUT_B16,
    input [15:0] SB_T0_SOUTH_SB_IN_B16,
    output [15:0] SB_T0_SOUTH_SB_OUT_B16,
    input [15:0] SB_T0_WEST_SB_IN_B16,
    output [15:0] SB_T0_WEST_SB_OUT_B16,
    input [15:0] SB_T1_EAST_SB_IN_B16,
    output [15:0] SB_T1_EAST_SB_OUT_B16,
    input [15:0] SB_T1_NORTH_SB_IN_B16,
    output [15:0] SB_T1_NORTH_SB_OUT_B16,
    input [15:0] SB_T1_SOUTH_SB_IN_B16,
    output [15:0] SB_T1_SOUTH_SB_OUT_B16,
    input [15:0] SB_T1_WEST_SB_IN_B16,
    output [15:0] SB_T1_WEST_SB_OUT_B16,
    input [15:0] SB_T2_EAST_SB_IN_B16,
    output [15:0] SB_T2_EAST_SB_OUT_B16,
    input [15:0] SB_T2_NORTH_SB_IN_B16,
    output [15:0] SB_T2_NORTH_SB_OUT_B16,
    input [15:0] SB_T2_SOUTH_SB_IN_B16,
    output [15:0] SB_T2_SOUTH_SB_OUT_B16,
    input [15:0] SB_T2_WEST_SB_IN_B16,
    output [15:0] SB_T2_WEST_SB_OUT_B16,
    input [15:0] SB_T3_EAST_SB_IN_B16,
    output [15:0] SB_T3_EAST_SB_OUT_B16,
    input [15:0] SB_T3_NORTH_SB_IN_B16,
    output [15:0] SB_T3_NORTH_SB_OUT_B16,
    input [15:0] SB_T3_SOUTH_SB_IN_B16,
    output [15:0] SB_T3_SOUTH_SB_OUT_B16,
    input [15:0] SB_T3_WEST_SB_IN_B16,
    output [15:0] SB_T3_WEST_SB_OUT_B16,
    input [15:0] SB_T4_EAST_SB_IN_B16,
    output [15:0] SB_T4_EAST_SB_OUT_B16,
    input [15:0] SB_T4_NORTH_SB_IN_B16,
    output [15:0] SB_T4_NORTH_SB_OUT_B16,
    input [15:0] SB_T4_SOUTH_SB_IN_B16,
    output [15:0] SB_T4_SOUTH_SB_OUT_B16,
    input [15:0] SB_T4_WEST_SB_IN_B16,
    output [15:0] SB_T4_WEST_SB_OUT_B16,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    input [15:0] output_width_16_num_0,
    input [15:0] output_width_16_num_1,
    output [31:0] read_config_data,
    input reset,
    input [0:0] stall
);
wire [0:0] Invert1_inst0_out;
wire [15:0] MUX_SB_T0_EAST_SB_OUT_B16_O;
wire [15:0] MUX_SB_T0_NORTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T0_SOUTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T0_WEST_SB_OUT_B16_O;
wire [15:0] MUX_SB_T1_EAST_SB_OUT_B16_O;
wire [15:0] MUX_SB_T1_NORTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T1_SOUTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T1_WEST_SB_OUT_B16_O;
wire [15:0] MUX_SB_T2_EAST_SB_OUT_B16_O;
wire [15:0] MUX_SB_T2_NORTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T2_SOUTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T2_WEST_SB_OUT_B16_O;
wire [15:0] MUX_SB_T3_EAST_SB_OUT_B16_O;
wire [15:0] MUX_SB_T3_NORTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T3_SOUTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T3_WEST_SB_OUT_B16_O;
wire [15:0] MUX_SB_T4_EAST_SB_OUT_B16_O;
wire [15:0] MUX_SB_T4_NORTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T4_SOUTH_SB_OUT_B16_O;
wire [15:0] MUX_SB_T4_WEST_SB_OUT_B16_O;
wire [31:0] MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0_out;
wire [15:0] REG_T0_EAST_B16_O;
wire [15:0] REG_T0_NORTH_B16_O;
wire [15:0] REG_T0_SOUTH_B16_O;
wire [15:0] REG_T0_WEST_B16_O;
wire [15:0] REG_T1_EAST_B16_O;
wire [15:0] REG_T1_NORTH_B16_O;
wire [15:0] REG_T1_SOUTH_B16_O;
wire [15:0] REG_T1_WEST_B16_O;
wire [15:0] REG_T2_EAST_B16_O;
wire [15:0] REG_T2_NORTH_B16_O;
wire [15:0] REG_T2_SOUTH_B16_O;
wire [15:0] REG_T2_WEST_B16_O;
wire [15:0] REG_T3_EAST_B16_O;
wire [15:0] REG_T3_NORTH_B16_O;
wire [15:0] REG_T3_SOUTH_B16_O;
wire [15:0] REG_T3_WEST_B16_O;
wire [15:0] REG_T4_EAST_B16_O;
wire [15:0] REG_T4_NORTH_B16_O;
wire [15:0] REG_T4_SOUTH_B16_O;
wire [15:0] REG_T4_WEST_B16_O;
wire [15:0] RMUX_T0_EAST_B16_O;
wire [0:0] RMUX_T0_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T0_NORTH_B16_O;
wire [0:0] RMUX_T0_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T0_SOUTH_B16_O;
wire [0:0] RMUX_T0_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T0_WEST_B16_O;
wire [0:0] RMUX_T0_WEST_B16_sel_inst0_O;
wire [15:0] RMUX_T1_EAST_B16_O;
wire [0:0] RMUX_T1_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T1_NORTH_B16_O;
wire [0:0] RMUX_T1_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T1_SOUTH_B16_O;
wire [0:0] RMUX_T1_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T1_WEST_B16_O;
wire [0:0] RMUX_T1_WEST_B16_sel_inst0_O;
wire [15:0] RMUX_T2_EAST_B16_O;
wire [0:0] RMUX_T2_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T2_NORTH_B16_O;
wire [0:0] RMUX_T2_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T2_SOUTH_B16_O;
wire [0:0] RMUX_T2_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T2_WEST_B16_O;
wire [0:0] RMUX_T2_WEST_B16_sel_inst0_O;
wire [15:0] RMUX_T3_EAST_B16_O;
wire [0:0] RMUX_T3_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T3_NORTH_B16_O;
wire [0:0] RMUX_T3_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T3_SOUTH_B16_O;
wire [0:0] RMUX_T3_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T3_WEST_B16_O;
wire [0:0] RMUX_T3_WEST_B16_sel_inst0_O;
wire [15:0] RMUX_T4_EAST_B16_O;
wire [0:0] RMUX_T4_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T4_NORTH_B16_O;
wire [0:0] RMUX_T4_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T4_SOUTH_B16_O;
wire [0:0] RMUX_T4_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T4_WEST_B16_O;
wire [0:0] RMUX_T4_WEST_B16_sel_inst0_O;
wire [2:0] SB_T0_EAST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T0_NORTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T0_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T0_WEST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T1_EAST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T1_NORTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T1_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T1_WEST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T2_EAST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T2_NORTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T2_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T2_WEST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T3_EAST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T3_NORTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T3_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T3_WEST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T4_EAST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T4_NORTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T4_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T4_WEST_SB_OUT_B16_sel_inst0_O;
wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T3_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T3_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T3_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T3_WEST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T4_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T4_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T4_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T4_WEST_SB_IN_B16_O;
wire ZextWrapper_18_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_18_32_inst0$self_O_in;
wire ZextWrapper_30_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_30_32_inst0$self_O_in;
wire [0:0] and1_inst0_out;
wire [0:0] and1_inst1_out;
wire [0:0] and1_inst10_out;
wire [0:0] and1_inst11_out;
wire [0:0] and1_inst12_out;
wire [0:0] and1_inst13_out;
wire [0:0] and1_inst14_out;
wire [0:0] and1_inst15_out;
wire [0:0] and1_inst16_out;
wire [0:0] and1_inst17_out;
wire [0:0] and1_inst18_out;
wire [0:0] and1_inst19_out;
wire [0:0] and1_inst2_out;
wire [0:0] and1_inst3_out;
wire [0:0] and1_inst4_out;
wire [0:0] and1_inst5_out;
wire [0:0] and1_inst6_out;
wire [0:0] and1_inst7_out;
wire [0:0] and1_inst8_out;
wire [0:0] and1_inst9_out;
wire [31:0] config_reg_0_O;
wire [29:0] config_reg_1_O;
wire [17:0] config_reg_2_O;
wire [0:0] const_1_1_out;
wire coreir_eq_1_inst0_out;
wire coreir_eq_1_inst1_out;
wire coreir_eq_1_inst10_out;
wire coreir_eq_1_inst11_out;
wire coreir_eq_1_inst12_out;
wire coreir_eq_1_inst13_out;
wire coreir_eq_1_inst14_out;
wire coreir_eq_1_inst15_out;
wire coreir_eq_1_inst16_out;
wire coreir_eq_1_inst17_out;
wire coreir_eq_1_inst18_out;
wire coreir_eq_1_inst19_out;
wire coreir_eq_1_inst2_out;
wire coreir_eq_1_inst3_out;
wire coreir_eq_1_inst4_out;
wire coreir_eq_1_inst5_out;
wire coreir_eq_1_inst6_out;
wire coreir_eq_1_inst7_out;
wire coreir_eq_1_inst8_out;
wire coreir_eq_1_inst9_out;
wire [7:0] self_config_config_addr_out;
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(stall),
    .out(Invert1_inst0_out)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T0_EAST_SB_OUT_B16 (
    .I_0(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_1(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T0_EAST_SB_OUT_B16_O),
    .S(SB_T0_EAST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T0_NORTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_1(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T0_NORTH_SB_OUT_B16_O),
    .S(SB_T0_NORTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T0_SOUTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T0_SOUTH_SB_OUT_B16_O),
    .S(SB_T0_SOUTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T0_WEST_SB_OUT_B16 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T0_WEST_SB_OUT_B16_O),
    .S(SB_T0_WEST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T1_EAST_SB_OUT_B16 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T1_EAST_SB_OUT_B16_O),
    .S(SB_T1_EAST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T1_NORTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_1(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T1_NORTH_SB_OUT_B16_O),
    .S(SB_T1_NORTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T1_SOUTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_1(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T1_SOUTH_SB_OUT_B16_O),
    .S(SB_T1_SOUTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T1_WEST_SB_OUT_B16 (
    .I_0(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T1_WEST_SB_OUT_B16_O),
    .S(SB_T1_WEST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T2_EAST_SB_OUT_B16 (
    .I_0(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T2_EAST_SB_OUT_B16_O),
    .S(SB_T2_EAST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T2_NORTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_1(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T2_NORTH_SB_OUT_B16_O),
    .S(SB_T2_NORTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T2_SOUTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_1(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T2_SOUTH_SB_OUT_B16_O),
    .S(SB_T2_SOUTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T2_WEST_SB_OUT_B16 (
    .I_0(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T2_WEST_SB_OUT_B16_O),
    .S(SB_T2_WEST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T3_EAST_SB_OUT_B16 (
    .I_0(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T3_EAST_SB_OUT_B16_O),
    .S(SB_T3_EAST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T3_NORTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_1(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_2(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T3_NORTH_SB_OUT_B16_O),
    .S(SB_T3_NORTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T3_SOUTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_1(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T3_SOUTH_SB_OUT_B16_O),
    .S(SB_T3_SOUTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T3_WEST_SB_OUT_B16 (
    .I_0(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T3_WEST_SB_OUT_B16_O),
    .S(SB_T3_WEST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T4_EAST_SB_OUT_B16 (
    .I_0(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T4_EAST_SB_OUT_B16_O),
    .S(SB_T4_EAST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T4_NORTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_2(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T4_NORTH_SB_OUT_B16_O),
    .S(SB_T4_NORTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T4_SOUTH_SB_OUT_B16 (
    .I_0(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_1(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_2(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T4_SOUTH_SB_OUT_B16_O),
    .S(SB_T4_SOUTH_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_5_16 MUX_SB_T4_WEST_SB_OUT_B16 (
    .I_0(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_2(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_3(output_width_16_num_0),
    .I_4(output_width_16_num_1),
    .O(MUX_SB_T4_WEST_SB_OUT_B16_O),
    .S(SB_T4_WEST_SB_OUT_B16_sel_inst0_O)
);
commonlib_muxn__N3__width32 MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0 (
    .in_data_0(config_reg_0_O),
    .in_data_1(ZextWrapper_30_32_inst0$self_O_in),
    .in_data_2(ZextWrapper_18_32_inst0$self_O_in),
    .in_sel(self_config_config_addr_out[1:0]),
    .out(MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0_out)
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_EAST_B16 (
    .I(MUX_SB_T0_EAST_SB_OUT_B16_O),
    .O(REG_T0_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst2_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_NORTH_B16 (
    .I(MUX_SB_T0_NORTH_SB_OUT_B16_O),
    .O(REG_T0_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst0_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_SOUTH_B16 (
    .I(MUX_SB_T0_SOUTH_SB_OUT_B16_O),
    .O(REG_T0_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst1_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_WEST_B16 (
    .I(MUX_SB_T0_WEST_SB_OUT_B16_O),
    .O(REG_T0_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst3_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_EAST_B16 (
    .I(MUX_SB_T1_EAST_SB_OUT_B16_O),
    .O(REG_T1_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst6_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_NORTH_B16 (
    .I(MUX_SB_T1_NORTH_SB_OUT_B16_O),
    .O(REG_T1_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst4_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_SOUTH_B16 (
    .I(MUX_SB_T1_SOUTH_SB_OUT_B16_O),
    .O(REG_T1_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst5_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_WEST_B16 (
    .I(MUX_SB_T1_WEST_SB_OUT_B16_O),
    .O(REG_T1_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst7_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_EAST_B16 (
    .I(MUX_SB_T2_EAST_SB_OUT_B16_O),
    .O(REG_T2_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst10_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_NORTH_B16 (
    .I(MUX_SB_T2_NORTH_SB_OUT_B16_O),
    .O(REG_T2_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst8_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_SOUTH_B16 (
    .I(MUX_SB_T2_SOUTH_SB_OUT_B16_O),
    .O(REG_T2_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst9_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_WEST_B16 (
    .I(MUX_SB_T2_WEST_SB_OUT_B16_O),
    .O(REG_T2_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst11_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T3_EAST_B16 (
    .I(MUX_SB_T3_EAST_SB_OUT_B16_O),
    .O(REG_T3_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst14_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T3_NORTH_B16 (
    .I(MUX_SB_T3_NORTH_SB_OUT_B16_O),
    .O(REG_T3_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst12_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T3_SOUTH_B16 (
    .I(MUX_SB_T3_SOUTH_SB_OUT_B16_O),
    .O(REG_T3_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst13_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T3_WEST_B16 (
    .I(MUX_SB_T3_WEST_SB_OUT_B16_O),
    .O(REG_T3_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst15_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T4_EAST_B16 (
    .I(MUX_SB_T4_EAST_SB_OUT_B16_O),
    .O(REG_T4_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst18_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T4_NORTH_B16 (
    .I(MUX_SB_T4_NORTH_SB_OUT_B16_O),
    .O(REG_T4_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst16_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T4_SOUTH_B16 (
    .I(MUX_SB_T4_SOUTH_SB_OUT_B16_O),
    .O(REG_T4_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst17_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T4_WEST_B16 (
    .I(MUX_SB_T4_WEST_SB_OUT_B16_O),
    .O(REG_T4_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst19_out[0])
);
MuxWrapperAOIImpl_2_16 RMUX_T0_EAST_B16 (
    .I_0(MUX_SB_T0_EAST_SB_OUT_B16_O),
    .I_1(REG_T0_EAST_B16_O),
    .O(RMUX_T0_EAST_B16_O),
    .S(RMUX_T0_EAST_B16_sel_inst0_O)
);
RMUX_T0_EAST_B16_sel RMUX_T0_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_EAST_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T0_NORTH_B16 (
    .I_0(MUX_SB_T0_NORTH_SB_OUT_B16_O),
    .I_1(REG_T0_NORTH_B16_O),
    .O(RMUX_T0_NORTH_B16_O),
    .S(RMUX_T0_NORTH_B16_sel_inst0_O)
);
RMUX_T0_NORTH_B16_sel RMUX_T0_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_NORTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T0_SOUTH_B16 (
    .I_0(MUX_SB_T0_SOUTH_SB_OUT_B16_O),
    .I_1(REG_T0_SOUTH_B16_O),
    .O(RMUX_T0_SOUTH_B16_O),
    .S(RMUX_T0_SOUTH_B16_sel_inst0_O)
);
RMUX_T0_SOUTH_B16_sel RMUX_T0_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_SOUTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T0_WEST_B16 (
    .I_0(MUX_SB_T0_WEST_SB_OUT_B16_O),
    .I_1(REG_T0_WEST_B16_O),
    .O(RMUX_T0_WEST_B16_O),
    .S(RMUX_T0_WEST_B16_sel_inst0_O)
);
RMUX_T0_WEST_B16_sel RMUX_T0_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_WEST_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T1_EAST_B16 (
    .I_0(MUX_SB_T1_EAST_SB_OUT_B16_O),
    .I_1(REG_T1_EAST_B16_O),
    .O(RMUX_T1_EAST_B16_O),
    .S(RMUX_T1_EAST_B16_sel_inst0_O)
);
RMUX_T1_EAST_B16_sel RMUX_T1_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_EAST_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T1_NORTH_B16 (
    .I_0(MUX_SB_T1_NORTH_SB_OUT_B16_O),
    .I_1(REG_T1_NORTH_B16_O),
    .O(RMUX_T1_NORTH_B16_O),
    .S(RMUX_T1_NORTH_B16_sel_inst0_O)
);
RMUX_T1_NORTH_B16_sel RMUX_T1_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_NORTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T1_SOUTH_B16 (
    .I_0(MUX_SB_T1_SOUTH_SB_OUT_B16_O),
    .I_1(REG_T1_SOUTH_B16_O),
    .O(RMUX_T1_SOUTH_B16_O),
    .S(RMUX_T1_SOUTH_B16_sel_inst0_O)
);
RMUX_T1_SOUTH_B16_sel RMUX_T1_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_SOUTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T1_WEST_B16 (
    .I_0(MUX_SB_T1_WEST_SB_OUT_B16_O),
    .I_1(REG_T1_WEST_B16_O),
    .O(RMUX_T1_WEST_B16_O),
    .S(RMUX_T1_WEST_B16_sel_inst0_O)
);
RMUX_T1_WEST_B16_sel RMUX_T1_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_WEST_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T2_EAST_B16 (
    .I_0(MUX_SB_T2_EAST_SB_OUT_B16_O),
    .I_1(REG_T2_EAST_B16_O),
    .O(RMUX_T2_EAST_B16_O),
    .S(RMUX_T2_EAST_B16_sel_inst0_O)
);
RMUX_T2_EAST_B16_sel RMUX_T2_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_EAST_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T2_NORTH_B16 (
    .I_0(MUX_SB_T2_NORTH_SB_OUT_B16_O),
    .I_1(REG_T2_NORTH_B16_O),
    .O(RMUX_T2_NORTH_B16_O),
    .S(RMUX_T2_NORTH_B16_sel_inst0_O)
);
RMUX_T2_NORTH_B16_sel RMUX_T2_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_NORTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T2_SOUTH_B16 (
    .I_0(MUX_SB_T2_SOUTH_SB_OUT_B16_O),
    .I_1(REG_T2_SOUTH_B16_O),
    .O(RMUX_T2_SOUTH_B16_O),
    .S(RMUX_T2_SOUTH_B16_sel_inst0_O)
);
RMUX_T2_SOUTH_B16_sel RMUX_T2_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_SOUTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T2_WEST_B16 (
    .I_0(MUX_SB_T2_WEST_SB_OUT_B16_O),
    .I_1(REG_T2_WEST_B16_O),
    .O(RMUX_T2_WEST_B16_O),
    .S(RMUX_T2_WEST_B16_sel_inst0_O)
);
RMUX_T2_WEST_B16_sel RMUX_T2_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_WEST_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T3_EAST_B16 (
    .I_0(MUX_SB_T3_EAST_SB_OUT_B16_O),
    .I_1(REG_T3_EAST_B16_O),
    .O(RMUX_T3_EAST_B16_O),
    .S(RMUX_T3_EAST_B16_sel_inst0_O)
);
RMUX_T3_EAST_B16_sel RMUX_T3_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_EAST_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T3_NORTH_B16 (
    .I_0(MUX_SB_T3_NORTH_SB_OUT_B16_O),
    .I_1(REG_T3_NORTH_B16_O),
    .O(RMUX_T3_NORTH_B16_O),
    .S(RMUX_T3_NORTH_B16_sel_inst0_O)
);
RMUX_T3_NORTH_B16_sel RMUX_T3_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_NORTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T3_SOUTH_B16 (
    .I_0(MUX_SB_T3_SOUTH_SB_OUT_B16_O),
    .I_1(REG_T3_SOUTH_B16_O),
    .O(RMUX_T3_SOUTH_B16_O),
    .S(RMUX_T3_SOUTH_B16_sel_inst0_O)
);
RMUX_T3_SOUTH_B16_sel RMUX_T3_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_SOUTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T3_WEST_B16 (
    .I_0(MUX_SB_T3_WEST_SB_OUT_B16_O),
    .I_1(REG_T3_WEST_B16_O),
    .O(RMUX_T3_WEST_B16_O),
    .S(RMUX_T3_WEST_B16_sel_inst0_O)
);
RMUX_T3_WEST_B16_sel RMUX_T3_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_WEST_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T4_EAST_B16 (
    .I_0(MUX_SB_T4_EAST_SB_OUT_B16_O),
    .I_1(REG_T4_EAST_B16_O),
    .O(RMUX_T4_EAST_B16_O),
    .S(RMUX_T4_EAST_B16_sel_inst0_O)
);
RMUX_T4_EAST_B16_sel RMUX_T4_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_EAST_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T4_NORTH_B16 (
    .I_0(MUX_SB_T4_NORTH_SB_OUT_B16_O),
    .I_1(REG_T4_NORTH_B16_O),
    .O(RMUX_T4_NORTH_B16_O),
    .S(RMUX_T4_NORTH_B16_sel_inst0_O)
);
RMUX_T4_NORTH_B16_sel RMUX_T4_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_NORTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T4_SOUTH_B16 (
    .I_0(MUX_SB_T4_SOUTH_SB_OUT_B16_O),
    .I_1(REG_T4_SOUTH_B16_O),
    .O(RMUX_T4_SOUTH_B16_O),
    .S(RMUX_T4_SOUTH_B16_sel_inst0_O)
);
RMUX_T4_SOUTH_B16_sel RMUX_T4_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_SOUTH_B16_sel_inst0_O)
);
MuxWrapperAOIImpl_2_16 RMUX_T4_WEST_B16 (
    .I_0(MUX_SB_T4_WEST_SB_OUT_B16_O),
    .I_1(REG_T4_WEST_B16_O),
    .O(RMUX_T4_WEST_B16_O),
    .S(RMUX_T4_WEST_B16_sel_inst0_O)
);
RMUX_T4_WEST_B16_sel RMUX_T4_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_WEST_B16_sel_inst0_O)
);
SB_T0_EAST_SB_OUT_B16_sel SB_T0_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T0_NORTH_SB_OUT_B16_sel SB_T0_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T0_SOUTH_SB_OUT_B16_sel SB_T0_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T0_WEST_SB_OUT_B16_sel SB_T0_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_WEST_SB_OUT_B16_sel_inst0_O)
);
SB_T1_EAST_SB_OUT_B16_sel SB_T1_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T1_NORTH_SB_OUT_B16_sel SB_T1_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T1_SOUTH_SB_OUT_B16_sel SB_T1_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T1_WEST_SB_OUT_B16_sel SB_T1_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_WEST_SB_OUT_B16_sel_inst0_O)
);
SB_T2_EAST_SB_OUT_B16_sel SB_T2_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T2_NORTH_SB_OUT_B16_sel SB_T2_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T2_SOUTH_SB_OUT_B16_sel SB_T2_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T2_WEST_SB_OUT_B16_sel SB_T2_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_WEST_SB_OUT_B16_sel_inst0_O)
);
SB_T3_EAST_SB_OUT_B16_sel SB_T3_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T3_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T3_NORTH_SB_OUT_B16_sel SB_T3_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T3_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T3_SOUTH_SB_OUT_B16_sel SB_T3_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T3_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T3_WEST_SB_OUT_B16_sel SB_T3_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T3_WEST_SB_OUT_B16_sel_inst0_O)
);
SB_T4_EAST_SB_OUT_B16_sel SB_T4_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T4_NORTH_SB_OUT_B16_sel SB_T4_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T4_SOUTH_SB_OUT_B16_sel SB_T4_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T4_WEST_SB_OUT_B16_sel SB_T4_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_WEST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T0_EAST_SB_IN_B16 (
    .I(SB_T0_EAST_SB_IN_B16),
    .O(WIRE_SB_T0_EAST_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T0_NORTH_SB_IN_B16 (
    .I(SB_T0_NORTH_SB_IN_B16),
    .O(WIRE_SB_T0_NORTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T0_SOUTH_SB_IN_B16 (
    .I(SB_T0_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T0_WEST_SB_IN_B16 (
    .I(SB_T0_WEST_SB_IN_B16),
    .O(WIRE_SB_T0_WEST_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T1_EAST_SB_IN_B16 (
    .I(SB_T1_EAST_SB_IN_B16),
    .O(WIRE_SB_T1_EAST_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T1_NORTH_SB_IN_B16 (
    .I(SB_T1_NORTH_SB_IN_B16),
    .O(WIRE_SB_T1_NORTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T1_SOUTH_SB_IN_B16 (
    .I(SB_T1_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T1_WEST_SB_IN_B16 (
    .I(SB_T1_WEST_SB_IN_B16),
    .O(WIRE_SB_T1_WEST_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T2_EAST_SB_IN_B16 (
    .I(SB_T2_EAST_SB_IN_B16),
    .O(WIRE_SB_T2_EAST_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T2_NORTH_SB_IN_B16 (
    .I(SB_T2_NORTH_SB_IN_B16),
    .O(WIRE_SB_T2_NORTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T2_SOUTH_SB_IN_B16 (
    .I(SB_T2_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T2_WEST_SB_IN_B16 (
    .I(SB_T2_WEST_SB_IN_B16),
    .O(WIRE_SB_T2_WEST_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T3_EAST_SB_IN_B16 (
    .I(SB_T3_EAST_SB_IN_B16),
    .O(WIRE_SB_T3_EAST_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T3_NORTH_SB_IN_B16 (
    .I(SB_T3_NORTH_SB_IN_B16),
    .O(WIRE_SB_T3_NORTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T3_SOUTH_SB_IN_B16 (
    .I(SB_T3_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T3_WEST_SB_IN_B16 (
    .I(SB_T3_WEST_SB_IN_B16),
    .O(WIRE_SB_T3_WEST_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T4_EAST_SB_IN_B16 (
    .I(SB_T4_EAST_SB_IN_B16),
    .O(WIRE_SB_T4_EAST_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T4_NORTH_SB_IN_B16 (
    .I(SB_T4_NORTH_SB_IN_B16),
    .O(WIRE_SB_T4_NORTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T4_SOUTH_SB_IN_B16 (
    .I(SB_T4_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B16_O)
);
MuxWrapperAOI_1_16_Regular WIRE_SB_T4_WEST_SB_IN_B16 (
    .I(SB_T4_WEST_SB_IN_B16),
    .O(WIRE_SB_T4_WEST_SB_IN_B16_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_18_32_inst0$bit_const_0_None (
    .out(ZextWrapper_18_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_18_32_inst0$self_O_out;
assign ZextWrapper_18_32_inst0$self_O_out = {ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,config_reg_2_O};
mantle_wire__typeBitIn32 ZextWrapper_18_32_inst0$self_O (
    .in(ZextWrapper_18_32_inst0$self_O_in),
    .out(ZextWrapper_18_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_30_32_inst0$bit_const_0_None (
    .out(ZextWrapper_30_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_30_32_inst0$self_O_out;
assign ZextWrapper_30_32_inst0$self_O_out = {ZextWrapper_30_32_inst0$bit_const_0_None_out,ZextWrapper_30_32_inst0$bit_const_0_None_out,config_reg_1_O};
mantle_wire__typeBitIn32 ZextWrapper_30_32_inst0$self_O (
    .in(ZextWrapper_30_32_inst0$self_O_in),
    .out(ZextWrapper_30_32_inst0$self_O_out)
);
coreir_and #(
    .width(1)
) and1_inst0 (
    .in0(coreir_eq_1_inst0_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst0_out)
);
coreir_and #(
    .width(1)
) and1_inst1 (
    .in0(coreir_eq_1_inst1_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst1_out)
);
coreir_and #(
    .width(1)
) and1_inst10 (
    .in0(coreir_eq_1_inst10_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst10_out)
);
coreir_and #(
    .width(1)
) and1_inst11 (
    .in0(coreir_eq_1_inst11_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst11_out)
);
coreir_and #(
    .width(1)
) and1_inst12 (
    .in0(coreir_eq_1_inst12_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst12_out)
);
coreir_and #(
    .width(1)
) and1_inst13 (
    .in0(coreir_eq_1_inst13_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst13_out)
);
coreir_and #(
    .width(1)
) and1_inst14 (
    .in0(coreir_eq_1_inst14_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst14_out)
);
coreir_and #(
    .width(1)
) and1_inst15 (
    .in0(coreir_eq_1_inst15_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst15_out)
);
coreir_and #(
    .width(1)
) and1_inst16 (
    .in0(coreir_eq_1_inst16_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst16_out)
);
coreir_and #(
    .width(1)
) and1_inst17 (
    .in0(coreir_eq_1_inst17_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst17_out)
);
coreir_and #(
    .width(1)
) and1_inst18 (
    .in0(coreir_eq_1_inst18_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst18_out)
);
coreir_and #(
    .width(1)
) and1_inst19 (
    .in0(coreir_eq_1_inst19_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst19_out)
);
coreir_and #(
    .width(1)
) and1_inst2 (
    .in0(coreir_eq_1_inst2_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst2_out)
);
coreir_and #(
    .width(1)
) and1_inst3 (
    .in0(coreir_eq_1_inst3_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst3_out)
);
coreir_and #(
    .width(1)
) and1_inst4 (
    .in0(coreir_eq_1_inst4_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst4_out)
);
coreir_and #(
    .width(1)
) and1_inst5 (
    .in0(coreir_eq_1_inst5_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst5_out)
);
coreir_and #(
    .width(1)
) and1_inst6 (
    .in0(coreir_eq_1_inst6_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst6_out)
);
coreir_and #(
    .width(1)
) and1_inst7 (
    .in0(coreir_eq_1_inst7_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst7_out)
);
coreir_and #(
    .width(1)
) and1_inst8 (
    .in0(coreir_eq_1_inst8_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst8_out)
);
coreir_and #(
    .width(1)
) and1_inst9 (
    .in0(coreir_eq_1_inst9_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst9_out)
);
wire [7:0] config_reg_0_config_addr;
assign config_reg_0_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2],self_config_config_addr_out[1:0]};
ConfigRegister_32_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_reg_0_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_1_config_addr;
assign config_reg_1_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2],self_config_config_addr_out[1:0]};
ConfigRegister_30_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_reg_1_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_2_config_addr;
assign config_reg_2_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2],self_config_config_addr_out[1:0]};
ConfigRegister_18_8_32_2 config_reg_2 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_2_O),
    .config_addr(config_reg_2_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst0 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst0_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst1 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst10 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst10_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst11 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst11_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst12 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst12_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst13 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst13_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst14 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst14_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst15 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst15_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst16 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst16_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst17 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst17_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst18 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst18_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst19 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst19_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst2 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst2_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst3 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst3_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst4 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst4_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst5 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst5_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst6 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst6_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst7 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst7_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst8 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst8_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst9 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst9_out)
);
mantle_wire__typeBit8 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
assign SB_T0_EAST_SB_OUT_B16 = RMUX_T0_EAST_B16_O;
assign SB_T0_NORTH_SB_OUT_B16 = RMUX_T0_NORTH_B16_O;
assign SB_T0_SOUTH_SB_OUT_B16 = RMUX_T0_SOUTH_B16_O;
assign SB_T0_WEST_SB_OUT_B16 = RMUX_T0_WEST_B16_O;
assign SB_T1_EAST_SB_OUT_B16 = RMUX_T1_EAST_B16_O;
assign SB_T1_NORTH_SB_OUT_B16 = RMUX_T1_NORTH_B16_O;
assign SB_T1_SOUTH_SB_OUT_B16 = RMUX_T1_SOUTH_B16_O;
assign SB_T1_WEST_SB_OUT_B16 = RMUX_T1_WEST_B16_O;
assign SB_T2_EAST_SB_OUT_B16 = RMUX_T2_EAST_B16_O;
assign SB_T2_NORTH_SB_OUT_B16 = RMUX_T2_NORTH_B16_O;
assign SB_T2_SOUTH_SB_OUT_B16 = RMUX_T2_SOUTH_B16_O;
assign SB_T2_WEST_SB_OUT_B16 = RMUX_T2_WEST_B16_O;
assign SB_T3_EAST_SB_OUT_B16 = RMUX_T3_EAST_B16_O;
assign SB_T3_NORTH_SB_OUT_B16 = RMUX_T3_NORTH_B16_O;
assign SB_T3_SOUTH_SB_OUT_B16 = RMUX_T3_SOUTH_B16_O;
assign SB_T3_WEST_SB_OUT_B16 = RMUX_T3_WEST_B16_O;
assign SB_T4_EAST_SB_OUT_B16 = RMUX_T4_EAST_B16_O;
assign SB_T4_NORTH_SB_OUT_B16 = RMUX_T4_NORTH_B16_O;
assign SB_T4_SOUTH_SB_OUT_B16 = RMUX_T4_SOUTH_B16_O;
assign SB_T4_WEST_SB_OUT_B16 = RMUX_T4_WEST_B16_O;
assign read_config_data = MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0_out;
endmodule

module ConfigRegister_17_8_32_78 (
    input clk,
    input reset,
    output [16:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [16:0] Register_inst0_O;
wire [7:0] const_78_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq3 Register_inst0 (
    .I(config_data[16:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h4e),
    .width(8)
) const_78_8 (
    .out(const_78_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_78_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_17_8_32_7 (
    input clk,
    input reset,
    output [16:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [16:0] Register_inst0_O;
wire [7:0] const_7_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq3 Register_inst0 (
    .I(config_data[16:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h07),
    .width(8)
) const_7_8 (
    .out(const_7_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_7_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_17_8_32_61 (
    input clk,
    input reset,
    output [16:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [16:0] Register_inst0_O;
wire [7:0] const_61_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq3 Register_inst0 (
    .I(config_data[16:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h3d),
    .width(8)
) const_61_8 (
    .out(const_61_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_61_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_17_8_32_57 (
    input clk,
    input reset,
    output [16:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [16:0] Register_inst0_O;
wire [7:0] const_57_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq3 Register_inst0 (
    .I(config_data[16:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h39),
    .width(8)
) const_57_8 (
    .out(const_57_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_57_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_17_8_32_30 (
    input clk,
    input reset,
    output [16:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [16:0] Register_inst0_O;
wire [7:0] const_30_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq3 Register_inst0 (
    .I(config_data[16:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h1e),
    .width(8)
) const_30_8 (
    .out(const_30_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_30_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_17_8_32_3 (
    input clk,
    input reset,
    output [16:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [16:0] Register_inst0_O;
wire [7:0] const_3_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq3 Register_inst0 (
    .I(config_data[16:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h03),
    .width(8)
) const_3_8 (
    .out(const_3_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_3_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_17_8_32_26 (
    input clk,
    input reset,
    output [16:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [16:0] Register_inst0_O;
wire [7:0] const_26_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq3 Register_inst0 (
    .I(config_data[16:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h1a),
    .width(8)
) const_26_8 (
    .out(const_26_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_26_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_17_8_32_2 (
    input clk,
    input reset,
    output [16:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [16:0] Register_inst0_O;
wire [7:0] const_2_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq3 Register_inst0 (
    .I(config_data[16:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h02),
    .width(8)
) const_2_8 (
    .out(const_2_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_2_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module PondCore (
    input clk,
    input [7:0] config_1_config_addr,
    input [31:0] config_1_config_data,
    input [0:0] config_1_read,
    input [0:0] config_1_write,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input config_en_0,
    input [0:0] config_read,
    input [0:0] config_write,
    input [15:0] data_in_pond,
    output [15:0] data_out_pond,
    input [0:0] flush,
    input [0:0] flush_core,
    output [31:0] read_config_data,
    output [31:0] read_config_data_1,
    input reset,
    input [0:0] stall,
    output [0:0] valid_out_pond
);
wire [0:0] AND_CONFIG_EN_SRAM_0_out;
wire [0:0] Invert1_inst0_out;
wire [0:0] Invert1_inst1_out;
wire [31:0] MuxWrapper_11_32_inst0$Mux11xBits32_inst0$coreir_commonlib_mux11x32_inst0_out;
wire [0:0] OR_CONFIG_EN_SRAM_0_out;
wire OR_CONFIG_RD_SRAM$orr_inst0_out;
wire OR_CONFIG_WR_SRAM$orr_inst0_out;
wire [7:0] OR_config_addr_FEATURE_out;
wire [31:0] OR_config_data_FEATURE_out;
wire ZextWrapper_17_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_17_32_inst0$self_O_in;
wire ZextWrapper_17_32_inst1$bit_const_0_None_out;
wire [31:0] ZextWrapper_17_32_inst1$self_O_in;
wire ZextWrapper_1_32_inst0$bit_const_0_None_out;
wire ZextWrapper_23_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_23_32_inst0$self_O_in;
wire ZextWrapper_24_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_24_32_inst0$self_O_in;
wire [23:0] config_reg_0_O;
wire [31:0] config_reg_1_O;
wire [0:0] config_reg_10_O;
wire [16:0] config_reg_2_O;
wire [31:0] config_reg_3_O;
wire [31:0] config_reg_4_O;
wire [22:0] config_reg_5_O;
wire [31:0] config_reg_6_O;
wire [16:0] config_reg_7_O;
wire [31:0] config_reg_8_O;
wire [31:0] config_reg_9_O;
wire coreir_wrapInAsyncReset_inst0_out;
wire coreir_wrapOutAsyncReset_inst0_out;
wire [0:0] flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] flush_mux_sel_inst0_O;
wire [31:0] pond_W_inst0_config_data_out;
wire [0:0] pond_W_inst0_valid_out_pond;
wire [15:0] pond_W_inst0_data_out_pond;
wire [4:0] rf_read_addr_0_starting_addr_inst0_O;
wire [4:0] rf_read_addr_0_strides_0_inst0_O;
wire [4:0] rf_read_addr_0_strides_1_inst0_O;
wire [4:0] rf_read_addr_0_strides_2_inst0_O;
wire [2:0] rf_read_iter_0_dimensionality_inst0_O;
wire [15:0] rf_read_iter_0_ranges_0_inst0_O;
wire [15:0] rf_read_iter_0_ranges_1_inst0_O;
wire [15:0] rf_read_iter_0_ranges_2_inst0_O;
wire [0:0] rf_read_sched_0_enable_inst0_O;
wire [15:0] rf_read_sched_0_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] rf_read_sched_0_sched_addr_gen_strides_0_inst0_O;
wire [15:0] rf_read_sched_0_sched_addr_gen_strides_1_inst0_O;
wire [15:0] rf_read_sched_0_sched_addr_gen_strides_2_inst0_O;
wire [4:0] rf_write_addr_0_starting_addr_inst0_O;
wire [4:0] rf_write_addr_0_strides_0_inst0_O;
wire [4:0] rf_write_addr_0_strides_1_inst0_O;
wire [4:0] rf_write_addr_0_strides_2_inst0_O;
wire [2:0] rf_write_iter_0_dimensionality_inst0_O;
wire [15:0] rf_write_iter_0_ranges_0_inst0_O;
wire [15:0] rf_write_iter_0_ranges_1_inst0_O;
wire [15:0] rf_write_iter_0_ranges_2_inst0_O;
wire [0:0] rf_write_sched_0_enable_inst0_O;
wire [15:0] rf_write_sched_0_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] rf_write_sched_0_sched_addr_gen_strides_0_inst0_O;
wire [15:0] rf_write_sched_0_sched_addr_gen_strides_1_inst0_O;
wire [15:0] rf_write_sched_0_sched_addr_gen_strides_2_inst0_O;
wire [7:0] self_config_config_addr_out;
wire [0:0] tile_en_inst0_O;
coreir_and #(
    .width(1)
) AND_CONFIG_EN_SRAM_0 (
    .in0(OR_CONFIG_EN_SRAM_0_out),
    .in1(config_en_0),
    .out(AND_CONFIG_EN_SRAM_0_out)
);
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(coreir_wrapInAsyncReset_inst0_out),
    .out(Invert1_inst0_out)
);
coreir_not #(
    .width(1)
) Invert1_inst1 (
    .in(stall),
    .out(Invert1_inst1_out)
);
wire [31:0] MuxWrapper_11_32_inst0$Mux11xBits32_inst0$coreir_commonlib_mux11x32_inst0_in_data_10;
assign MuxWrapper_11_32_inst0$Mux11xBits32_inst0$coreir_commonlib_mux11x32_inst0_in_data_10 = {ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,config_reg_10_O[0]};
commonlib_muxn__N11__width32 MuxWrapper_11_32_inst0$Mux11xBits32_inst0$coreir_commonlib_mux11x32_inst0 (
    .in_data_0(ZextWrapper_24_32_inst0$self_O_in),
    .in_data_1(config_reg_1_O),
    .in_data_10(MuxWrapper_11_32_inst0$Mux11xBits32_inst0$coreir_commonlib_mux11x32_inst0_in_data_10),
    .in_data_2(ZextWrapper_17_32_inst0$self_O_in),
    .in_data_3(config_reg_3_O),
    .in_data_4(config_reg_4_O),
    .in_data_5(ZextWrapper_23_32_inst0$self_O_in),
    .in_data_6(config_reg_6_O),
    .in_data_7(ZextWrapper_17_32_inst1$self_O_in),
    .in_data_8(config_reg_8_O),
    .in_data_9(config_reg_9_O),
    .in_sel(self_config_config_addr_out[3:0]),
    .out(MuxWrapper_11_32_inst0$Mux11xBits32_inst0$coreir_commonlib_mux11x32_inst0_out)
);
coreir_or #(
    .width(1)
) OR_CONFIG_EN_SRAM_0 (
    .in0(config_1_write),
    .in1(config_1_read),
    .out(OR_CONFIG_EN_SRAM_0_out)
);
coreir_orr #(
    .width(1)
) OR_CONFIG_RD_SRAM$orr_inst0 (
    .in(config_1_write),
    .out(OR_CONFIG_RD_SRAM$orr_inst0_out)
);
coreir_orr #(
    .width(1)
) OR_CONFIG_WR_SRAM$orr_inst0 (
    .in(config_1_read),
    .out(OR_CONFIG_WR_SRAM$orr_inst0_out)
);
wire [7:0] OR_config_addr_FEATURE_in0;
assign OR_config_addr_FEATURE_in0 = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3:0]};
coreir_or #(
    .width(8)
) OR_config_addr_FEATURE (
    .in0(OR_config_addr_FEATURE_in0),
    .in1(config_1_config_addr),
    .out(OR_config_addr_FEATURE_out)
);
coreir_or #(
    .width(32)
) OR_config_data_FEATURE (
    .in0(config_config_data),
    .in1(config_1_config_data),
    .out(OR_config_data_FEATURE_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_17_32_inst0$bit_const_0_None (
    .out(ZextWrapper_17_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_17_32_inst0$self_O_out;
assign ZextWrapper_17_32_inst0$self_O_out = {ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,config_reg_2_O};
mantle_wire__typeBitIn32 ZextWrapper_17_32_inst0$self_O (
    .in(ZextWrapper_17_32_inst0$self_O_in),
    .out(ZextWrapper_17_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_17_32_inst1$bit_const_0_None (
    .out(ZextWrapper_17_32_inst1$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_17_32_inst1$self_O_out;
assign ZextWrapper_17_32_inst1$self_O_out = {ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,config_reg_7_O};
mantle_wire__typeBitIn32 ZextWrapper_17_32_inst1$self_O (
    .in(ZextWrapper_17_32_inst1$self_O_in),
    .out(ZextWrapper_17_32_inst1$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_1_32_inst0$bit_const_0_None (
    .out(ZextWrapper_1_32_inst0$bit_const_0_None_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_23_32_inst0$bit_const_0_None (
    .out(ZextWrapper_23_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_23_32_inst0$self_O_out;
assign ZextWrapper_23_32_inst0$self_O_out = {ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,config_reg_5_O};
mantle_wire__typeBitIn32 ZextWrapper_23_32_inst0$self_O (
    .in(ZextWrapper_23_32_inst0$self_O_in),
    .out(ZextWrapper_23_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_24_32_inst0$bit_const_0_None (
    .out(ZextWrapper_24_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_24_32_inst0$self_O_out;
assign ZextWrapper_24_32_inst0$self_O_out = {ZextWrapper_24_32_inst0$bit_const_0_None_out,ZextWrapper_24_32_inst0$bit_const_0_None_out,ZextWrapper_24_32_inst0$bit_const_0_None_out,ZextWrapper_24_32_inst0$bit_const_0_None_out,ZextWrapper_24_32_inst0$bit_const_0_None_out,ZextWrapper_24_32_inst0$bit_const_0_None_out,ZextWrapper_24_32_inst0$bit_const_0_None_out,ZextWrapper_24_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_24_32_inst0$self_O (
    .in(ZextWrapper_24_32_inst0$self_O_in),
    .out(ZextWrapper_24_32_inst0$self_O_out)
);
wire [7:0] config_reg_0_config_addr;
assign config_reg_0_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3:0]};
ConfigRegister_24_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_reg_0_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_1_config_addr;
assign config_reg_1_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3:0]};
ConfigRegister_32_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_reg_1_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_10_config_addr;
assign config_reg_10_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3:0]};
ConfigRegister_1_8_32_10 config_reg_10 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_10_O),
    .config_addr(config_reg_10_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_2_config_addr;
assign config_reg_2_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3:0]};
ConfigRegister_17_8_32_2 config_reg_2 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_2_O),
    .config_addr(config_reg_2_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_3_config_addr;
assign config_reg_3_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3:0]};
ConfigRegister_32_8_32_3 config_reg_3 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_3_O),
    .config_addr(config_reg_3_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_4_config_addr;
assign config_reg_4_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3:0]};
ConfigRegister_32_8_32_4 config_reg_4 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_4_O),
    .config_addr(config_reg_4_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_5_config_addr;
assign config_reg_5_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3:0]};
ConfigRegister_23_8_32_5 config_reg_5 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_5_O),
    .config_addr(config_reg_5_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_6_config_addr;
assign config_reg_6_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3:0]};
ConfigRegister_32_8_32_6 config_reg_6 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_6_O),
    .config_addr(config_reg_6_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_7_config_addr;
assign config_reg_7_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3:0]};
ConfigRegister_17_8_32_7 config_reg_7 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_7_O),
    .config_addr(config_reg_7_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_8_config_addr;
assign config_reg_8_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3:0]};
ConfigRegister_32_8_32_8 config_reg_8 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_8_O),
    .config_addr(config_reg_8_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_9_config_addr;
assign config_reg_9_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3:0]};
ConfigRegister_32_8_32_9 config_reg_9 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_9_O),
    .config_addr(config_reg_9_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_wrap coreir_wrapInAsyncReset_inst0 (
    .in(reset),
    .out(coreir_wrapInAsyncReset_inst0_out)
);
coreir_wrap coreir_wrapOutAsyncReset_inst0 (
    .in(Invert1_inst0_out[0]),
    .out(coreir_wrapOutAsyncReset_inst0_out)
);
coreir_mux #(
    .width(1)
) flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(flush_core),
    .in1(flush),
    .sel(flush_mux_sel_inst0_O[0]),
    .out(flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
flush_mux_sel flush_mux_sel_inst0 (
    .I(config_reg_0_O),
    .O(flush_mux_sel_inst0_O)
);
pond_W pond_W_inst0 (
    .rf_write_addr_0_strides_1(rf_write_addr_0_strides_1_inst0_O),
    .rf_read_sched_0_sched_addr_gen_strides_1(rf_read_sched_0_sched_addr_gen_strides_1_inst0_O),
    .rf_read_addr_0_starting_addr(rf_read_addr_0_starting_addr_inst0_O),
    .rf_read_sched_0_sched_addr_gen_starting_addr(rf_read_sched_0_sched_addr_gen_starting_addr_inst0_O),
    .config_data_out(pond_W_inst0_config_data_out),
    .rf_write_iter_0_ranges_2(rf_write_iter_0_ranges_2_inst0_O),
    .clk(clk),
    .rf_read_sched_0_sched_addr_gen_strides_0(rf_read_sched_0_sched_addr_gen_strides_0_inst0_O),
    .rf_read_iter_0_ranges_2(rf_read_iter_0_ranges_2_inst0_O),
    .rf_write_sched_0_sched_addr_gen_strides_1(rf_write_sched_0_sched_addr_gen_strides_1_inst0_O),
    .rf_read_sched_0_enable(rf_read_sched_0_enable_inst0_O),
    .rf_write_iter_0_ranges_0(rf_write_iter_0_ranges_0_inst0_O),
    .rf_read_iter_0_dimensionality(rf_read_iter_0_dimensionality_inst0_O),
    .rf_write_iter_0_ranges_1(rf_write_iter_0_ranges_1_inst0_O),
    .rf_write_sched_0_sched_addr_gen_starting_addr(rf_write_sched_0_sched_addr_gen_starting_addr_inst0_O),
    .config_write(OR_CONFIG_RD_SRAM$orr_inst0_out),
    .rf_read_sched_0_sched_addr_gen_strides_2(rf_read_sched_0_sched_addr_gen_strides_2_inst0_O),
    .rf_write_addr_0_starting_addr(rf_write_addr_0_starting_addr_inst0_O),
    .rf_read_iter_0_ranges_1(rf_read_iter_0_ranges_1_inst0_O),
    .rf_write_addr_0_strides_0(rf_write_addr_0_strides_0_inst0_O),
    .config_data_in(OR_config_data_FEATURE_out),
    .valid_out_pond(pond_W_inst0_valid_out_pond),
    .rf_write_sched_0_sched_addr_gen_strides_0(rf_write_sched_0_sched_addr_gen_strides_0_inst0_O),
    .config_read(OR_CONFIG_WR_SRAM$orr_inst0_out),
    .clk_en(Invert1_inst1_out),
    .rf_read_addr_0_strides_0(rf_read_addr_0_strides_0_inst0_O),
    .data_out_pond(pond_W_inst0_data_out_pond),
    .config_addr_in(OR_config_addr_FEATURE_out),
    .rf_read_addr_0_strides_1(rf_read_addr_0_strides_1_inst0_O),
    .rf_write_sched_0_enable(rf_write_sched_0_enable_inst0_O),
    .rst_n(coreir_wrapOutAsyncReset_inst0_out),
    .rf_read_addr_0_strides_2(rf_read_addr_0_strides_2_inst0_O),
    .data_in_pond(data_in_pond),
    .rf_write_addr_0_strides_2(rf_write_addr_0_strides_2_inst0_O),
    .tile_en(tile_en_inst0_O),
    .config_en(AND_CONFIG_EN_SRAM_0_out),
    .rf_read_iter_0_ranges_0(rf_read_iter_0_ranges_0_inst0_O),
    .flush(flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .rf_write_iter_0_dimensionality(rf_write_iter_0_dimensionality_inst0_O),
    .rf_write_sched_0_sched_addr_gen_strides_2(rf_write_sched_0_sched_addr_gen_strides_2_inst0_O)
);
rf_read_addr_0_starting_addr rf_read_addr_0_starting_addr_inst0 (
    .I(config_reg_0_O),
    .O(rf_read_addr_0_starting_addr_inst0_O)
);
rf_read_addr_0_strides_0 rf_read_addr_0_strides_0_inst0 (
    .I(config_reg_0_O),
    .O(rf_read_addr_0_strides_0_inst0_O)
);
rf_read_addr_0_strides_1 rf_read_addr_0_strides_1_inst0 (
    .I(config_reg_0_O),
    .O(rf_read_addr_0_strides_1_inst0_O)
);
rf_read_addr_0_strides_2 rf_read_addr_0_strides_2_inst0 (
    .I(config_reg_0_O),
    .O(rf_read_addr_0_strides_2_inst0_O)
);
rf_read_iter_0_dimensionality rf_read_iter_0_dimensionality_inst0 (
    .I(config_reg_0_O),
    .O(rf_read_iter_0_dimensionality_inst0_O)
);
rf_read_iter_0_ranges_0 rf_read_iter_0_ranges_0_inst0 (
    .I(config_reg_1_O),
    .O(rf_read_iter_0_ranges_0_inst0_O)
);
rf_read_iter_0_ranges_1 rf_read_iter_0_ranges_1_inst0 (
    .I(config_reg_1_O),
    .O(rf_read_iter_0_ranges_1_inst0_O)
);
rf_read_iter_0_ranges_2 rf_read_iter_0_ranges_2_inst0 (
    .I(config_reg_2_O),
    .O(rf_read_iter_0_ranges_2_inst0_O)
);
rf_read_sched_0_enable rf_read_sched_0_enable_inst0 (
    .I(config_reg_2_O),
    .O(rf_read_sched_0_enable_inst0_O)
);
rf_read_sched_0_sched_addr_gen_starting_addr rf_read_sched_0_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_3_O),
    .O(rf_read_sched_0_sched_addr_gen_starting_addr_inst0_O)
);
rf_read_sched_0_sched_addr_gen_strides_0 rf_read_sched_0_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_3_O),
    .O(rf_read_sched_0_sched_addr_gen_strides_0_inst0_O)
);
rf_read_sched_0_sched_addr_gen_strides_1 rf_read_sched_0_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_4_O),
    .O(rf_read_sched_0_sched_addr_gen_strides_1_inst0_O)
);
rf_read_sched_0_sched_addr_gen_strides_2 rf_read_sched_0_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_4_O),
    .O(rf_read_sched_0_sched_addr_gen_strides_2_inst0_O)
);
rf_write_addr_0_starting_addr rf_write_addr_0_starting_addr_inst0 (
    .I(config_reg_5_O),
    .O(rf_write_addr_0_starting_addr_inst0_O)
);
rf_write_addr_0_strides_0 rf_write_addr_0_strides_0_inst0 (
    .I(config_reg_5_O),
    .O(rf_write_addr_0_strides_0_inst0_O)
);
rf_write_addr_0_strides_1 rf_write_addr_0_strides_1_inst0 (
    .I(config_reg_5_O),
    .O(rf_write_addr_0_strides_1_inst0_O)
);
rf_write_addr_0_strides_2 rf_write_addr_0_strides_2_inst0 (
    .I(config_reg_5_O),
    .O(rf_write_addr_0_strides_2_inst0_O)
);
rf_write_iter_0_dimensionality rf_write_iter_0_dimensionality_inst0 (
    .I(config_reg_5_O),
    .O(rf_write_iter_0_dimensionality_inst0_O)
);
rf_write_iter_0_ranges_0 rf_write_iter_0_ranges_0_inst0 (
    .I(config_reg_6_O),
    .O(rf_write_iter_0_ranges_0_inst0_O)
);
rf_write_iter_0_ranges_1 rf_write_iter_0_ranges_1_inst0 (
    .I(config_reg_6_O),
    .O(rf_write_iter_0_ranges_1_inst0_O)
);
rf_write_iter_0_ranges_2 rf_write_iter_0_ranges_2_inst0 (
    .I(config_reg_7_O),
    .O(rf_write_iter_0_ranges_2_inst0_O)
);
rf_write_sched_0_enable rf_write_sched_0_enable_inst0 (
    .I(config_reg_7_O),
    .O(rf_write_sched_0_enable_inst0_O)
);
rf_write_sched_0_sched_addr_gen_starting_addr rf_write_sched_0_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_8_O),
    .O(rf_write_sched_0_sched_addr_gen_starting_addr_inst0_O)
);
rf_write_sched_0_sched_addr_gen_strides_0 rf_write_sched_0_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_8_O),
    .O(rf_write_sched_0_sched_addr_gen_strides_0_inst0_O)
);
rf_write_sched_0_sched_addr_gen_strides_1 rf_write_sched_0_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_9_O),
    .O(rf_write_sched_0_sched_addr_gen_strides_1_inst0_O)
);
rf_write_sched_0_sched_addr_gen_strides_2 rf_write_sched_0_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_9_O),
    .O(rf_write_sched_0_sched_addr_gen_strides_2_inst0_O)
);
mantle_wire__typeBit8 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
tile_en tile_en_inst0 (
    .I(config_reg_10_O),
    .O(tile_en_inst0_O)
);
assign data_out_pond = pond_W_inst0_data_out_pond;
assign read_config_data = MuxWrapper_11_32_inst0$Mux11xBits32_inst0$coreir_commonlib_mux11x32_inst0_out;
assign read_config_data_1 = pond_W_inst0_config_data_out;
assign valid_out_pond = pond_W_inst0_valid_out_pond;
endmodule

module ConfigRegister_17_8_32_15 (
    input clk,
    input reset,
    output [16:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [16:0] Register_inst0_O;
wire [7:0] const_15_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq3 Register_inst0 (
    .I(config_data[16:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0f),
    .width(8)
) const_15_8 (
    .out(const_15_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_15_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_17_8_32_11 (
    input clk,
    input reset,
    output [16:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [16:0] Register_inst0_O;
wire [7:0] const_11_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq3 Register_inst0 (
    .I(config_data[16:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0b),
    .width(8)
) const_11_8 (
    .out(const_11_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_11_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module MemCore (
    input clk,
    input [7:0] config_1_config_addr,
    input [31:0] config_1_config_data,
    input [0:0] config_1_read,
    input [0:0] config_1_write,
    input [7:0] config_2_config_addr,
    input [31:0] config_2_config_data,
    input [0:0] config_2_read,
    input [0:0] config_2_write,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input config_en_0,
    input config_en_1,
    input [0:0] config_read,
    input [0:0] config_write,
    input [0:0] flush,
    input [0:0] flush_core,
    input [15:0] input_width_16_num_0,
    input [15:0] input_width_16_num_1,
    input [15:0] input_width_16_num_2,
    input [15:0] input_width_16_num_3,
    input [0:0] input_width_1_num_0,
    input [0:0] input_width_1_num_1,
    output [15:0] output_width_16_num_0,
    output [15:0] output_width_16_num_1,
    output [0:0] output_width_1_num_0,
    output [0:0] output_width_1_num_1,
    output [0:0] output_width_1_num_2,
    output [0:0] output_width_1_num_3,
    output [31:0] read_config_data,
    output [31:0] read_config_data_1,
    output [31:0] read_config_data_2,
    input reset,
    input [0:0] stall
);
wire [0:0] AND_CONFIG_EN_SRAM_0_out;
wire [0:0] AND_CONFIG_EN_SRAM_1_out;
wire [0:0] Invert1_inst0_out;
wire [0:0] Invert1_inst1_out;
wire [0:0] LakeTop_W_inst0_output_width_1_num_3;
wire [31:0] LakeTop_W_inst0_config_data_out_1;
wire [15:0] LakeTop_W_inst0_output_width_16_num_1;
wire [0:0] LakeTop_W_inst0_output_width_1_num_0;
wire [15:0] LakeTop_W_inst0_output_width_16_num_0;
wire [31:0] LakeTop_W_inst0_config_data_out_0;
wire [0:0] LakeTop_W_inst0_output_width_1_num_2;
wire [0:0] LakeTop_W_inst0_output_width_1_num_1;
wire [31:0] MuxWrapper_84_32_inst0$Mux84xBits32_inst0$coreir_commonlib_mux84x32_inst0_out;
wire [0:0] OR_CONFIG_EN_SRAM_0_out;
wire [0:0] OR_CONFIG_EN_SRAM_1_out;
wire [0:0] OR_CONFIG_RD_SRAM_out;
wire [0:0] OR_CONFIG_WR_SRAM_out;
wire [7:0] OR_config_addr_FEATURE_O;
wire [31:0] OR_config_data_FEATURE_O;
wire ZextWrapper_17_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_17_32_inst0$self_O_in;
wire ZextWrapper_17_32_inst1$bit_const_0_None_out;
wire [31:0] ZextWrapper_17_32_inst1$self_O_in;
wire ZextWrapper_17_32_inst2$bit_const_0_None_out;
wire [31:0] ZextWrapper_17_32_inst2$self_O_in;
wire ZextWrapper_17_32_inst3$bit_const_0_None_out;
wire [31:0] ZextWrapper_17_32_inst3$self_O_in;
wire ZextWrapper_17_32_inst4$bit_const_0_None_out;
wire [31:0] ZextWrapper_17_32_inst4$self_O_in;
wire ZextWrapper_17_32_inst5$bit_const_0_None_out;
wire [31:0] ZextWrapper_17_32_inst5$self_O_in;
wire ZextWrapper_17_32_inst6$bit_const_0_None_out;
wire [31:0] ZextWrapper_17_32_inst6$self_O_in;
wire ZextWrapper_17_32_inst7$bit_const_0_None_out;
wire [31:0] ZextWrapper_17_32_inst7$self_O_in;
wire ZextWrapper_20_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_20_32_inst0$self_O_in;
wire ZextWrapper_20_32_inst1$bit_const_0_None_out;
wire [31:0] ZextWrapper_20_32_inst1$self_O_in;
wire ZextWrapper_20_32_inst2$bit_const_0_None_out;
wire [31:0] ZextWrapper_20_32_inst2$self_O_in;
wire ZextWrapper_20_32_inst3$bit_const_0_None_out;
wire [31:0] ZextWrapper_20_32_inst3$self_O_in;
wire ZextWrapper_20_32_inst4$bit_const_0_None_out;
wire [31:0] ZextWrapper_20_32_inst4$self_O_in;
wire ZextWrapper_20_32_inst5$bit_const_0_None_out;
wire [31:0] ZextWrapper_20_32_inst5$self_O_in;
wire ZextWrapper_20_32_inst6$bit_const_0_None_out;
wire [31:0] ZextWrapper_20_32_inst6$self_O_in;
wire ZextWrapper_25_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_25_32_inst0$self_O_in;
wire ZextWrapper_25_32_inst1$bit_const_0_None_out;
wire [31:0] ZextWrapper_25_32_inst1$self_O_in;
wire ZextWrapper_26_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_26_32_inst0$self_O_in;
wire ZextWrapper_27_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_27_32_inst0$self_O_in;
wire ZextWrapper_27_32_inst1$bit_const_0_None_out;
wire [31:0] ZextWrapper_27_32_inst1$self_O_in;
wire ZextWrapper_27_32_inst2$bit_const_0_None_out;
wire [31:0] ZextWrapper_27_32_inst2$self_O_in;
wire ZextWrapper_27_32_inst3$bit_const_0_None_out;
wire [31:0] ZextWrapper_27_32_inst3$self_O_in;
wire ZextWrapper_27_32_inst4$bit_const_0_None_out;
wire [31:0] ZextWrapper_27_32_inst4$self_O_in;
wire ZextWrapper_27_32_inst5$bit_const_0_None_out;
wire [31:0] ZextWrapper_27_32_inst5$self_O_in;
wire ZextWrapper_27_32_inst6$bit_const_0_None_out;
wire [31:0] ZextWrapper_27_32_inst6$self_O_in;
wire ZextWrapper_27_32_inst7$bit_const_0_None_out;
wire [31:0] ZextWrapper_27_32_inst7$self_O_in;
wire ZextWrapper_27_32_inst8$bit_const_0_None_out;
wire [31:0] ZextWrapper_27_32_inst8$self_O_in;
wire ZextWrapper_31_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_31_32_inst0$self_O_in;
wire [24:0] config_reg_0_O;
wire [31:0] config_reg_1_O;
wire [31:0] config_reg_10_O;
wire [16:0] config_reg_11_O;
wire [31:0] config_reg_12_O;
wire [31:0] config_reg_13_O;
wire [31:0] config_reg_14_O;
wire [16:0] config_reg_15_O;
wire [31:0] config_reg_16_O;
wire [31:0] config_reg_17_O;
wire [31:0] config_reg_18_O;
wire [19:0] config_reg_19_O;
wire [31:0] config_reg_2_O;
wire [31:0] config_reg_20_O;
wire [31:0] config_reg_21_O;
wire [31:0] config_reg_22_O;
wire [19:0] config_reg_23_O;
wire [31:0] config_reg_24_O;
wire [31:0] config_reg_25_O;
wire [16:0] config_reg_26_O;
wire [31:0] config_reg_27_O;
wire [31:0] config_reg_28_O;
wire [31:0] config_reg_29_O;
wire [16:0] config_reg_3_O;
wire [16:0] config_reg_30_O;
wire [31:0] config_reg_31_O;
wire [31:0] config_reg_32_O;
wire [31:0] config_reg_33_O;
wire [19:0] config_reg_34_O;
wire [31:0] config_reg_35_O;
wire [31:0] config_reg_36_O;
wire [31:0] config_reg_37_O;
wire [19:0] config_reg_38_O;
wire [31:0] config_reg_39_O;
wire [31:0] config_reg_4_O;
wire [31:0] config_reg_40_O;
wire [25:0] config_reg_41_O;
wire [26:0] config_reg_42_O;
wire [26:0] config_reg_43_O;
wire [26:0] config_reg_44_O;
wire [26:0] config_reg_45_O;
wire [26:0] config_reg_46_O;
wire [26:0] config_reg_47_O;
wire [26:0] config_reg_48_O;
wire [26:0] config_reg_49_O;
wire [31:0] config_reg_5_O;
wire [30:0] config_reg_50_O;
wire [31:0] config_reg_51_O;
wire [31:0] config_reg_52_O;
wire [31:0] config_reg_53_O;
wire [19:0] config_reg_54_O;
wire [31:0] config_reg_55_O;
wire [31:0] config_reg_56_O;
wire [16:0] config_reg_57_O;
wire [31:0] config_reg_58_O;
wire [31:0] config_reg_59_O;
wire [31:0] config_reg_6_O;
wire [31:0] config_reg_60_O;
wire [16:0] config_reg_61_O;
wire [31:0] config_reg_62_O;
wire [31:0] config_reg_63_O;
wire [31:0] config_reg_64_O;
wire [19:0] config_reg_65_O;
wire [31:0] config_reg_66_O;
wire [31:0] config_reg_67_O;
wire [31:0] config_reg_68_O;
wire [19:0] config_reg_69_O;
wire [31:0] config_reg_7_O;
wire [31:0] config_reg_70_O;
wire [31:0] config_reg_71_O;
wire [31:0] config_reg_72_O;
wire [31:0] config_reg_73_O;
wire [24:0] config_reg_74_O;
wire [31:0] config_reg_75_O;
wire [31:0] config_reg_76_O;
wire [31:0] config_reg_77_O;
wire [16:0] config_reg_78_O;
wire [31:0] config_reg_79_O;
wire [31:0] config_reg_8_O;
wire [31:0] config_reg_80_O;
wire [31:0] config_reg_81_O;
wire [31:0] config_reg_82_O;
wire [26:0] config_reg_83_O;
wire [31:0] config_reg_9_O;
wire coreir_wrapInAsyncReset_inst0_out;
wire coreir_wrapOutAsyncReset_inst0_out;
wire [0:0] flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] flush_mux_sel_inst0_O;
wire [0:0] input_width_1_num_0_reg_sel_inst0_O;
wire [0:0] input_width_1_num_0_reg_value_inst0_O;
wire [0:0] input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] input_width_1_num_1_reg_sel_inst0_O;
wire [0:0] input_width_1_num_1_reg_value_inst0_O;
wire [0:0] input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [3:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality_inst0_O;
wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0_inst0_O;
wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1_inst0_O;
wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2_inst0_O;
wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3_inst0_O;
wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4_inst0_O;
wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5_inst0_O;
wire [0:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable_inst0_O;
wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0_inst0_O;
wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1_inst0_O;
wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2_inst0_O;
wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3_inst0_O;
wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4_inst0_O;
wire [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5_inst0_O;
wire [15:0] mem_ctrl_strg_fifo_flat_strg_fifo_inst_fifo_depth_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5_inst0_O;
wire [0:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5_inst0_O;
wire [0:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5_inst0_O;
wire [0:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5_inst0_O;
wire [0:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5_inst0_O;
wire [0:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4_inst0_O;
wire [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5_inst0_O;
wire [0:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5_inst0_O;
wire [0:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5_inst0_O;
wire [0:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5_inst0_O;
wire [0:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4_inst0_O;
wire [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4_inst0_O;
wire [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5_inst0_O;
wire [1:0] mode_inst0_O;
wire [7:0] self_config_config_addr_out;
wire [0:0] tile_en_inst0_O;
coreir_and #(
    .width(1)
) AND_CONFIG_EN_SRAM_0 (
    .in0(OR_CONFIG_EN_SRAM_0_out),
    .in1(config_en_0),
    .out(AND_CONFIG_EN_SRAM_0_out)
);
coreir_and #(
    .width(1)
) AND_CONFIG_EN_SRAM_1 (
    .in0(OR_CONFIG_EN_SRAM_1_out),
    .in1(config_en_1),
    .out(AND_CONFIG_EN_SRAM_1_out)
);
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(coreir_wrapInAsyncReset_inst0_out),
    .out(Invert1_inst0_out)
);
coreir_not #(
    .width(1)
) Invert1_inst1 (
    .in(stall),
    .out(Invert1_inst1_out)
);
wire [1:0] LakeTop_W_inst0_config_en;
assign LakeTop_W_inst0_config_en = {AND_CONFIG_EN_SRAM_1_out[0],AND_CONFIG_EN_SRAM_0_out[0]};
LakeTop_W LakeTop_W_inst0 (
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr_inst0_O),
    .input_width_16_num_1(input_width_16_num_1),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2_inst0_O),
    .input_width_16_num_3(input_width_16_num_3),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2_inst0_O),
    .output_width_1_num_3(LakeTop_W_inst0_output_width_1_num_3),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5_inst0_O),
    .config_write(OR_CONFIG_RD_SRAM_out),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1_inst0_O),
    .mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0_inst0_O),
    .mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1_inst0_O),
    .mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2_inst0_O),
    .mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2_inst0_O),
    .mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4_inst0_O),
    .config_data_out_1(LakeTop_W_inst0_config_data_out_1),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr_inst0_O),
    .mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2_inst0_O),
    .input_width_16_num_2(input_width_16_num_2),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1_inst0_O),
    .input_width_1_num_1(input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0_inst0_O),
    .mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0_inst0_O),
    .output_width_16_num_1(LakeTop_W_inst0_output_width_16_num_1),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4_inst0_O),
    .output_width_1_num_0(LakeTop_W_inst0_output_width_1_num_0),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5_inst0_O),
    .output_width_16_num_0(LakeTop_W_inst0_output_width_16_num_0),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5_inst0_O),
    .mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0_inst0_O),
    .mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2_inst0_O),
    .flush(flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0_inst0_O),
    .input_width_1_num_0(input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr_inst0_O),
    .config_data_out_0(LakeTop_W_inst0_config_data_out_0),
    .clk(clk),
    .mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3_inst0_O),
    .mem_ctrl_strg_fifo_flat_strg_fifo_inst_fifo_depth(mem_ctrl_strg_fifo_flat_strg_fifo_inst_fifo_depth_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5_inst0_O),
    .clk_en(Invert1_inst1_out),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0_inst0_O),
    .output_width_1_num_2(LakeTop_W_inst0_output_width_1_num_2),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3_inst0_O),
    .output_width_1_num_1(LakeTop_W_inst0_output_width_1_num_1),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4_inst0_O),
    .mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality_inst0_O),
    .config_en(LakeTop_W_inst0_config_en),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0_inst0_O),
    .mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en_inst0_O),
    .mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0_inst0_O),
    .mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1_inst0_O),
    .config_data_in(OR_config_data_FEATURE_O),
    .mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3_inst0_O),
    .input_width_16_num_0(input_width_16_num_0),
    .config_read(OR_CONFIG_WR_SRAM_out),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0_inst0_O),
    .config_addr_in(OR_config_addr_FEATURE_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4_inst0_O),
    .rst_n(coreir_wrapOutAsyncReset_inst0_out),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1_inst0_O),
    .tile_en(tile_en_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr_inst0_O),
    .mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2_inst0_O),
    .mode(mode_inst0_O)
);
commonlib_muxn__N84__width32 MuxWrapper_84_32_inst0$Mux84xBits32_inst0$coreir_commonlib_mux84x32_inst0 (
    .in_data_0(ZextWrapper_25_32_inst0$self_O_in),
    .in_data_1(config_reg_1_O),
    .in_data_10(config_reg_10_O),
    .in_data_11(ZextWrapper_17_32_inst1$self_O_in),
    .in_data_12(config_reg_12_O),
    .in_data_13(config_reg_13_O),
    .in_data_14(config_reg_14_O),
    .in_data_15(ZextWrapper_17_32_inst2$self_O_in),
    .in_data_16(config_reg_16_O),
    .in_data_17(config_reg_17_O),
    .in_data_18(config_reg_18_O),
    .in_data_19(ZextWrapper_20_32_inst0$self_O_in),
    .in_data_2(config_reg_2_O),
    .in_data_20(config_reg_20_O),
    .in_data_21(config_reg_21_O),
    .in_data_22(config_reg_22_O),
    .in_data_23(ZextWrapper_20_32_inst1$self_O_in),
    .in_data_24(config_reg_24_O),
    .in_data_25(config_reg_25_O),
    .in_data_26(ZextWrapper_17_32_inst3$self_O_in),
    .in_data_27(config_reg_27_O),
    .in_data_28(config_reg_28_O),
    .in_data_29(config_reg_29_O),
    .in_data_3(ZextWrapper_17_32_inst0$self_O_in),
    .in_data_30(ZextWrapper_17_32_inst4$self_O_in),
    .in_data_31(config_reg_31_O),
    .in_data_32(config_reg_32_O),
    .in_data_33(config_reg_33_O),
    .in_data_34(ZextWrapper_20_32_inst2$self_O_in),
    .in_data_35(config_reg_35_O),
    .in_data_36(config_reg_36_O),
    .in_data_37(config_reg_37_O),
    .in_data_38(ZextWrapper_20_32_inst3$self_O_in),
    .in_data_39(config_reg_39_O),
    .in_data_4(config_reg_4_O),
    .in_data_40(config_reg_40_O),
    .in_data_41(ZextWrapper_26_32_inst0$self_O_in),
    .in_data_42(ZextWrapper_27_32_inst0$self_O_in),
    .in_data_43(ZextWrapper_27_32_inst1$self_O_in),
    .in_data_44(ZextWrapper_27_32_inst2$self_O_in),
    .in_data_45(ZextWrapper_27_32_inst3$self_O_in),
    .in_data_46(ZextWrapper_27_32_inst4$self_O_in),
    .in_data_47(ZextWrapper_27_32_inst5$self_O_in),
    .in_data_48(ZextWrapper_27_32_inst6$self_O_in),
    .in_data_49(ZextWrapper_27_32_inst7$self_O_in),
    .in_data_5(config_reg_5_O),
    .in_data_50(ZextWrapper_31_32_inst0$self_O_in),
    .in_data_51(config_reg_51_O),
    .in_data_52(config_reg_52_O),
    .in_data_53(config_reg_53_O),
    .in_data_54(ZextWrapper_20_32_inst4$self_O_in),
    .in_data_55(config_reg_55_O),
    .in_data_56(config_reg_56_O),
    .in_data_57(ZextWrapper_17_32_inst5$self_O_in),
    .in_data_58(config_reg_58_O),
    .in_data_59(config_reg_59_O),
    .in_data_6(config_reg_6_O),
    .in_data_60(config_reg_60_O),
    .in_data_61(ZextWrapper_17_32_inst6$self_O_in),
    .in_data_62(config_reg_62_O),
    .in_data_63(config_reg_63_O),
    .in_data_64(config_reg_64_O),
    .in_data_65(ZextWrapper_20_32_inst5$self_O_in),
    .in_data_66(config_reg_66_O),
    .in_data_67(config_reg_67_O),
    .in_data_68(config_reg_68_O),
    .in_data_69(ZextWrapper_20_32_inst6$self_O_in),
    .in_data_7(config_reg_7_O),
    .in_data_70(config_reg_70_O),
    .in_data_71(config_reg_71_O),
    .in_data_72(config_reg_72_O),
    .in_data_73(config_reg_73_O),
    .in_data_74(ZextWrapper_25_32_inst1$self_O_in),
    .in_data_75(config_reg_75_O),
    .in_data_76(config_reg_76_O),
    .in_data_77(config_reg_77_O),
    .in_data_78(ZextWrapper_17_32_inst7$self_O_in),
    .in_data_79(config_reg_79_O),
    .in_data_8(config_reg_8_O),
    .in_data_80(config_reg_80_O),
    .in_data_81(config_reg_81_O),
    .in_data_82(config_reg_82_O),
    .in_data_83(ZextWrapper_27_32_inst8$self_O_in),
    .in_data_9(config_reg_9_O),
    .in_sel(self_config_config_addr_out[6:0]),
    .out(MuxWrapper_84_32_inst0$Mux84xBits32_inst0$coreir_commonlib_mux84x32_inst0_out)
);
coreir_or #(
    .width(1)
) OR_CONFIG_EN_SRAM_0 (
    .in0(config_1_write),
    .in1(config_1_read),
    .out(OR_CONFIG_EN_SRAM_0_out)
);
coreir_or #(
    .width(1)
) OR_CONFIG_EN_SRAM_1 (
    .in0(config_2_write),
    .in1(config_2_read),
    .out(OR_CONFIG_EN_SRAM_1_out)
);
coreir_or #(
    .width(1)
) OR_CONFIG_RD_SRAM (
    .in0(config_1_write),
    .in1(config_2_write),
    .out(OR_CONFIG_RD_SRAM_out)
);
coreir_or #(
    .width(1)
) OR_CONFIG_WR_SRAM (
    .in0(config_1_read),
    .in1(config_2_read),
    .out(OR_CONFIG_WR_SRAM_out)
);
wire [7:0] OR_config_addr_FEATURE_I0;
assign OR_config_addr_FEATURE_I0 = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
Or3x8 OR_config_addr_FEATURE (
    .I0(OR_config_addr_FEATURE_I0),
    .I1(config_1_config_addr),
    .I2(config_2_config_addr),
    .O(OR_config_addr_FEATURE_O)
);
Or3x32 OR_config_data_FEATURE (
    .I0(config_config_data),
    .I1(config_1_config_data),
    .I2(config_2_config_data),
    .O(OR_config_data_FEATURE_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_17_32_inst0$bit_const_0_None (
    .out(ZextWrapper_17_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_17_32_inst0$self_O_out;
assign ZextWrapper_17_32_inst0$self_O_out = {ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,config_reg_3_O};
mantle_wire__typeBitIn32 ZextWrapper_17_32_inst0$self_O (
    .in(ZextWrapper_17_32_inst0$self_O_in),
    .out(ZextWrapper_17_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_17_32_inst1$bit_const_0_None (
    .out(ZextWrapper_17_32_inst1$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_17_32_inst1$self_O_out;
assign ZextWrapper_17_32_inst1$self_O_out = {ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,config_reg_11_O};
mantle_wire__typeBitIn32 ZextWrapper_17_32_inst1$self_O (
    .in(ZextWrapper_17_32_inst1$self_O_in),
    .out(ZextWrapper_17_32_inst1$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_17_32_inst2$bit_const_0_None (
    .out(ZextWrapper_17_32_inst2$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_17_32_inst2$self_O_out;
assign ZextWrapper_17_32_inst2$self_O_out = {ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,config_reg_15_O};
mantle_wire__typeBitIn32 ZextWrapper_17_32_inst2$self_O (
    .in(ZextWrapper_17_32_inst2$self_O_in),
    .out(ZextWrapper_17_32_inst2$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_17_32_inst3$bit_const_0_None (
    .out(ZextWrapper_17_32_inst3$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_17_32_inst3$self_O_out;
assign ZextWrapper_17_32_inst3$self_O_out = {ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,config_reg_26_O};
mantle_wire__typeBitIn32 ZextWrapper_17_32_inst3$self_O (
    .in(ZextWrapper_17_32_inst3$self_O_in),
    .out(ZextWrapper_17_32_inst3$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_17_32_inst4$bit_const_0_None (
    .out(ZextWrapper_17_32_inst4$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_17_32_inst4$self_O_out;
assign ZextWrapper_17_32_inst4$self_O_out = {ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,config_reg_30_O};
mantle_wire__typeBitIn32 ZextWrapper_17_32_inst4$self_O (
    .in(ZextWrapper_17_32_inst4$self_O_in),
    .out(ZextWrapper_17_32_inst4$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_17_32_inst5$bit_const_0_None (
    .out(ZextWrapper_17_32_inst5$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_17_32_inst5$self_O_out;
assign ZextWrapper_17_32_inst5$self_O_out = {ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,config_reg_57_O};
mantle_wire__typeBitIn32 ZextWrapper_17_32_inst5$self_O (
    .in(ZextWrapper_17_32_inst5$self_O_in),
    .out(ZextWrapper_17_32_inst5$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_17_32_inst6$bit_const_0_None (
    .out(ZextWrapper_17_32_inst6$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_17_32_inst6$self_O_out;
assign ZextWrapper_17_32_inst6$self_O_out = {ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,config_reg_61_O};
mantle_wire__typeBitIn32 ZextWrapper_17_32_inst6$self_O (
    .in(ZextWrapper_17_32_inst6$self_O_in),
    .out(ZextWrapper_17_32_inst6$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_17_32_inst7$bit_const_0_None (
    .out(ZextWrapper_17_32_inst7$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_17_32_inst7$self_O_out;
assign ZextWrapper_17_32_inst7$self_O_out = {ZextWrapper_17_32_inst7$bit_const_0_None_out,ZextWrapper_17_32_inst7$bit_const_0_None_out,ZextWrapper_17_32_inst7$bit_const_0_None_out,ZextWrapper_17_32_inst7$bit_const_0_None_out,ZextWrapper_17_32_inst7$bit_const_0_None_out,ZextWrapper_17_32_inst7$bit_const_0_None_out,ZextWrapper_17_32_inst7$bit_const_0_None_out,ZextWrapper_17_32_inst7$bit_const_0_None_out,ZextWrapper_17_32_inst7$bit_const_0_None_out,ZextWrapper_17_32_inst7$bit_const_0_None_out,ZextWrapper_17_32_inst7$bit_const_0_None_out,ZextWrapper_17_32_inst7$bit_const_0_None_out,ZextWrapper_17_32_inst7$bit_const_0_None_out,ZextWrapper_17_32_inst7$bit_const_0_None_out,ZextWrapper_17_32_inst7$bit_const_0_None_out,config_reg_78_O};
mantle_wire__typeBitIn32 ZextWrapper_17_32_inst7$self_O (
    .in(ZextWrapper_17_32_inst7$self_O_in),
    .out(ZextWrapper_17_32_inst7$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_20_32_inst0$bit_const_0_None (
    .out(ZextWrapper_20_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_20_32_inst0$self_O_out;
assign ZextWrapper_20_32_inst0$self_O_out = {ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,config_reg_19_O};
mantle_wire__typeBitIn32 ZextWrapper_20_32_inst0$self_O (
    .in(ZextWrapper_20_32_inst0$self_O_in),
    .out(ZextWrapper_20_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_20_32_inst1$bit_const_0_None (
    .out(ZextWrapper_20_32_inst1$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_20_32_inst1$self_O_out;
assign ZextWrapper_20_32_inst1$self_O_out = {ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,config_reg_23_O};
mantle_wire__typeBitIn32 ZextWrapper_20_32_inst1$self_O (
    .in(ZextWrapper_20_32_inst1$self_O_in),
    .out(ZextWrapper_20_32_inst1$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_20_32_inst2$bit_const_0_None (
    .out(ZextWrapper_20_32_inst2$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_20_32_inst2$self_O_out;
assign ZextWrapper_20_32_inst2$self_O_out = {ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,config_reg_34_O};
mantle_wire__typeBitIn32 ZextWrapper_20_32_inst2$self_O (
    .in(ZextWrapper_20_32_inst2$self_O_in),
    .out(ZextWrapper_20_32_inst2$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_20_32_inst3$bit_const_0_None (
    .out(ZextWrapper_20_32_inst3$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_20_32_inst3$self_O_out;
assign ZextWrapper_20_32_inst3$self_O_out = {ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,config_reg_38_O};
mantle_wire__typeBitIn32 ZextWrapper_20_32_inst3$self_O (
    .in(ZextWrapper_20_32_inst3$self_O_in),
    .out(ZextWrapper_20_32_inst3$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_20_32_inst4$bit_const_0_None (
    .out(ZextWrapper_20_32_inst4$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_20_32_inst4$self_O_out;
assign ZextWrapper_20_32_inst4$self_O_out = {ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,config_reg_54_O};
mantle_wire__typeBitIn32 ZextWrapper_20_32_inst4$self_O (
    .in(ZextWrapper_20_32_inst4$self_O_in),
    .out(ZextWrapper_20_32_inst4$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_20_32_inst5$bit_const_0_None (
    .out(ZextWrapper_20_32_inst5$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_20_32_inst5$self_O_out;
assign ZextWrapper_20_32_inst5$self_O_out = {ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,config_reg_65_O};
mantle_wire__typeBitIn32 ZextWrapper_20_32_inst5$self_O (
    .in(ZextWrapper_20_32_inst5$self_O_in),
    .out(ZextWrapper_20_32_inst5$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_20_32_inst6$bit_const_0_None (
    .out(ZextWrapper_20_32_inst6$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_20_32_inst6$self_O_out;
assign ZextWrapper_20_32_inst6$self_O_out = {ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,config_reg_69_O};
mantle_wire__typeBitIn32 ZextWrapper_20_32_inst6$self_O (
    .in(ZextWrapper_20_32_inst6$self_O_in),
    .out(ZextWrapper_20_32_inst6$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_25_32_inst0$bit_const_0_None (
    .out(ZextWrapper_25_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_25_32_inst0$self_O_out;
assign ZextWrapper_25_32_inst0$self_O_out = {ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_25_32_inst0$self_O (
    .in(ZextWrapper_25_32_inst0$self_O_in),
    .out(ZextWrapper_25_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_25_32_inst1$bit_const_0_None (
    .out(ZextWrapper_25_32_inst1$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_25_32_inst1$self_O_out;
assign ZextWrapper_25_32_inst1$self_O_out = {ZextWrapper_25_32_inst1$bit_const_0_None_out,ZextWrapper_25_32_inst1$bit_const_0_None_out,ZextWrapper_25_32_inst1$bit_const_0_None_out,ZextWrapper_25_32_inst1$bit_const_0_None_out,ZextWrapper_25_32_inst1$bit_const_0_None_out,ZextWrapper_25_32_inst1$bit_const_0_None_out,ZextWrapper_25_32_inst1$bit_const_0_None_out,config_reg_74_O};
mantle_wire__typeBitIn32 ZextWrapper_25_32_inst1$self_O (
    .in(ZextWrapper_25_32_inst1$self_O_in),
    .out(ZextWrapper_25_32_inst1$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_26_32_inst0$bit_const_0_None (
    .out(ZextWrapper_26_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_26_32_inst0$self_O_out;
assign ZextWrapper_26_32_inst0$self_O_out = {ZextWrapper_26_32_inst0$bit_const_0_None_out,ZextWrapper_26_32_inst0$bit_const_0_None_out,ZextWrapper_26_32_inst0$bit_const_0_None_out,ZextWrapper_26_32_inst0$bit_const_0_None_out,ZextWrapper_26_32_inst0$bit_const_0_None_out,ZextWrapper_26_32_inst0$bit_const_0_None_out,config_reg_41_O};
mantle_wire__typeBitIn32 ZextWrapper_26_32_inst0$self_O (
    .in(ZextWrapper_26_32_inst0$self_O_in),
    .out(ZextWrapper_26_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_27_32_inst0$bit_const_0_None (
    .out(ZextWrapper_27_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_27_32_inst0$self_O_out;
assign ZextWrapper_27_32_inst0$self_O_out = {ZextWrapper_27_32_inst0$bit_const_0_None_out,ZextWrapper_27_32_inst0$bit_const_0_None_out,ZextWrapper_27_32_inst0$bit_const_0_None_out,ZextWrapper_27_32_inst0$bit_const_0_None_out,ZextWrapper_27_32_inst0$bit_const_0_None_out,config_reg_42_O};
mantle_wire__typeBitIn32 ZextWrapper_27_32_inst0$self_O (
    .in(ZextWrapper_27_32_inst0$self_O_in),
    .out(ZextWrapper_27_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_27_32_inst1$bit_const_0_None (
    .out(ZextWrapper_27_32_inst1$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_27_32_inst1$self_O_out;
assign ZextWrapper_27_32_inst1$self_O_out = {ZextWrapper_27_32_inst1$bit_const_0_None_out,ZextWrapper_27_32_inst1$bit_const_0_None_out,ZextWrapper_27_32_inst1$bit_const_0_None_out,ZextWrapper_27_32_inst1$bit_const_0_None_out,ZextWrapper_27_32_inst1$bit_const_0_None_out,config_reg_43_O};
mantle_wire__typeBitIn32 ZextWrapper_27_32_inst1$self_O (
    .in(ZextWrapper_27_32_inst1$self_O_in),
    .out(ZextWrapper_27_32_inst1$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_27_32_inst2$bit_const_0_None (
    .out(ZextWrapper_27_32_inst2$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_27_32_inst2$self_O_out;
assign ZextWrapper_27_32_inst2$self_O_out = {ZextWrapper_27_32_inst2$bit_const_0_None_out,ZextWrapper_27_32_inst2$bit_const_0_None_out,ZextWrapper_27_32_inst2$bit_const_0_None_out,ZextWrapper_27_32_inst2$bit_const_0_None_out,ZextWrapper_27_32_inst2$bit_const_0_None_out,config_reg_44_O};
mantle_wire__typeBitIn32 ZextWrapper_27_32_inst2$self_O (
    .in(ZextWrapper_27_32_inst2$self_O_in),
    .out(ZextWrapper_27_32_inst2$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_27_32_inst3$bit_const_0_None (
    .out(ZextWrapper_27_32_inst3$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_27_32_inst3$self_O_out;
assign ZextWrapper_27_32_inst3$self_O_out = {ZextWrapper_27_32_inst3$bit_const_0_None_out,ZextWrapper_27_32_inst3$bit_const_0_None_out,ZextWrapper_27_32_inst3$bit_const_0_None_out,ZextWrapper_27_32_inst3$bit_const_0_None_out,ZextWrapper_27_32_inst3$bit_const_0_None_out,config_reg_45_O};
mantle_wire__typeBitIn32 ZextWrapper_27_32_inst3$self_O (
    .in(ZextWrapper_27_32_inst3$self_O_in),
    .out(ZextWrapper_27_32_inst3$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_27_32_inst4$bit_const_0_None (
    .out(ZextWrapper_27_32_inst4$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_27_32_inst4$self_O_out;
assign ZextWrapper_27_32_inst4$self_O_out = {ZextWrapper_27_32_inst4$bit_const_0_None_out,ZextWrapper_27_32_inst4$bit_const_0_None_out,ZextWrapper_27_32_inst4$bit_const_0_None_out,ZextWrapper_27_32_inst4$bit_const_0_None_out,ZextWrapper_27_32_inst4$bit_const_0_None_out,config_reg_46_O};
mantle_wire__typeBitIn32 ZextWrapper_27_32_inst4$self_O (
    .in(ZextWrapper_27_32_inst4$self_O_in),
    .out(ZextWrapper_27_32_inst4$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_27_32_inst5$bit_const_0_None (
    .out(ZextWrapper_27_32_inst5$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_27_32_inst5$self_O_out;
assign ZextWrapper_27_32_inst5$self_O_out = {ZextWrapper_27_32_inst5$bit_const_0_None_out,ZextWrapper_27_32_inst5$bit_const_0_None_out,ZextWrapper_27_32_inst5$bit_const_0_None_out,ZextWrapper_27_32_inst5$bit_const_0_None_out,ZextWrapper_27_32_inst5$bit_const_0_None_out,config_reg_47_O};
mantle_wire__typeBitIn32 ZextWrapper_27_32_inst5$self_O (
    .in(ZextWrapper_27_32_inst5$self_O_in),
    .out(ZextWrapper_27_32_inst5$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_27_32_inst6$bit_const_0_None (
    .out(ZextWrapper_27_32_inst6$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_27_32_inst6$self_O_out;
assign ZextWrapper_27_32_inst6$self_O_out = {ZextWrapper_27_32_inst6$bit_const_0_None_out,ZextWrapper_27_32_inst6$bit_const_0_None_out,ZextWrapper_27_32_inst6$bit_const_0_None_out,ZextWrapper_27_32_inst6$bit_const_0_None_out,ZextWrapper_27_32_inst6$bit_const_0_None_out,config_reg_48_O};
mantle_wire__typeBitIn32 ZextWrapper_27_32_inst6$self_O (
    .in(ZextWrapper_27_32_inst6$self_O_in),
    .out(ZextWrapper_27_32_inst6$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_27_32_inst7$bit_const_0_None (
    .out(ZextWrapper_27_32_inst7$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_27_32_inst7$self_O_out;
assign ZextWrapper_27_32_inst7$self_O_out = {ZextWrapper_27_32_inst7$bit_const_0_None_out,ZextWrapper_27_32_inst7$bit_const_0_None_out,ZextWrapper_27_32_inst7$bit_const_0_None_out,ZextWrapper_27_32_inst7$bit_const_0_None_out,ZextWrapper_27_32_inst7$bit_const_0_None_out,config_reg_49_O};
mantle_wire__typeBitIn32 ZextWrapper_27_32_inst7$self_O (
    .in(ZextWrapper_27_32_inst7$self_O_in),
    .out(ZextWrapper_27_32_inst7$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_27_32_inst8$bit_const_0_None (
    .out(ZextWrapper_27_32_inst8$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_27_32_inst8$self_O_out;
assign ZextWrapper_27_32_inst8$self_O_out = {ZextWrapper_27_32_inst8$bit_const_0_None_out,ZextWrapper_27_32_inst8$bit_const_0_None_out,ZextWrapper_27_32_inst8$bit_const_0_None_out,ZextWrapper_27_32_inst8$bit_const_0_None_out,ZextWrapper_27_32_inst8$bit_const_0_None_out,config_reg_83_O};
mantle_wire__typeBitIn32 ZextWrapper_27_32_inst8$self_O (
    .in(ZextWrapper_27_32_inst8$self_O_in),
    .out(ZextWrapper_27_32_inst8$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_31_32_inst0$bit_const_0_None (
    .out(ZextWrapper_31_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_31_32_inst0$self_O_out;
assign ZextWrapper_31_32_inst0$self_O_out = {ZextWrapper_31_32_inst0$bit_const_0_None_out,config_reg_50_O};
mantle_wire__typeBitIn32 ZextWrapper_31_32_inst0$self_O (
    .in(ZextWrapper_31_32_inst0$self_O_in),
    .out(ZextWrapper_31_32_inst0$self_O_out)
);
wire [7:0] config_reg_0_config_addr;
assign config_reg_0_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_25_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_reg_0_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_1_config_addr;
assign config_reg_1_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_reg_1_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_10_config_addr;
assign config_reg_10_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_10 config_reg_10 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_10_O),
    .config_addr(config_reg_10_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_11_config_addr;
assign config_reg_11_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_17_8_32_11 config_reg_11 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_11_O),
    .config_addr(config_reg_11_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_12_config_addr;
assign config_reg_12_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_12 config_reg_12 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_12_O),
    .config_addr(config_reg_12_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_13_config_addr;
assign config_reg_13_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_13 config_reg_13 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_13_O),
    .config_addr(config_reg_13_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_14_config_addr;
assign config_reg_14_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_14 config_reg_14 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_14_O),
    .config_addr(config_reg_14_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_15_config_addr;
assign config_reg_15_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_17_8_32_15 config_reg_15 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_15_O),
    .config_addr(config_reg_15_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_16_config_addr;
assign config_reg_16_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_16 config_reg_16 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_16_O),
    .config_addr(config_reg_16_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_17_config_addr;
assign config_reg_17_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_17 config_reg_17 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_17_O),
    .config_addr(config_reg_17_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_18_config_addr;
assign config_reg_18_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_18 config_reg_18 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_18_O),
    .config_addr(config_reg_18_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_19_config_addr;
assign config_reg_19_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_20_8_32_19 config_reg_19 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_19_O),
    .config_addr(config_reg_19_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_2_config_addr;
assign config_reg_2_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_2 config_reg_2 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_2_O),
    .config_addr(config_reg_2_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_20_config_addr;
assign config_reg_20_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_20 config_reg_20 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_20_O),
    .config_addr(config_reg_20_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_21_config_addr;
assign config_reg_21_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_21 config_reg_21 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_21_O),
    .config_addr(config_reg_21_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_22_config_addr;
assign config_reg_22_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_22 config_reg_22 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_22_O),
    .config_addr(config_reg_22_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_23_config_addr;
assign config_reg_23_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_20_8_32_23 config_reg_23 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_23_O),
    .config_addr(config_reg_23_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_24_config_addr;
assign config_reg_24_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_24 config_reg_24 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_24_O),
    .config_addr(config_reg_24_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_25_config_addr;
assign config_reg_25_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_25 config_reg_25 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_25_O),
    .config_addr(config_reg_25_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_26_config_addr;
assign config_reg_26_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_17_8_32_26 config_reg_26 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_26_O),
    .config_addr(config_reg_26_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_27_config_addr;
assign config_reg_27_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_27 config_reg_27 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_27_O),
    .config_addr(config_reg_27_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_28_config_addr;
assign config_reg_28_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_28 config_reg_28 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_28_O),
    .config_addr(config_reg_28_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_29_config_addr;
assign config_reg_29_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_29 config_reg_29 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_29_O),
    .config_addr(config_reg_29_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_3_config_addr;
assign config_reg_3_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_17_8_32_3 config_reg_3 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_3_O),
    .config_addr(config_reg_3_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_30_config_addr;
assign config_reg_30_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_17_8_32_30 config_reg_30 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_30_O),
    .config_addr(config_reg_30_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_31_config_addr;
assign config_reg_31_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_31 config_reg_31 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_31_O),
    .config_addr(config_reg_31_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_32_config_addr;
assign config_reg_32_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_32 config_reg_32 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_32_O),
    .config_addr(config_reg_32_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_33_config_addr;
assign config_reg_33_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_33 config_reg_33 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_33_O),
    .config_addr(config_reg_33_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_34_config_addr;
assign config_reg_34_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_20_8_32_34 config_reg_34 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_34_O),
    .config_addr(config_reg_34_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_35_config_addr;
assign config_reg_35_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_35 config_reg_35 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_35_O),
    .config_addr(config_reg_35_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_36_config_addr;
assign config_reg_36_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_36 config_reg_36 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_36_O),
    .config_addr(config_reg_36_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_37_config_addr;
assign config_reg_37_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_37 config_reg_37 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_37_O),
    .config_addr(config_reg_37_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_38_config_addr;
assign config_reg_38_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_20_8_32_38 config_reg_38 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_38_O),
    .config_addr(config_reg_38_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_39_config_addr;
assign config_reg_39_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_39 config_reg_39 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_39_O),
    .config_addr(config_reg_39_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_4_config_addr;
assign config_reg_4_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_4 config_reg_4 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_4_O),
    .config_addr(config_reg_4_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_40_config_addr;
assign config_reg_40_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_40 config_reg_40 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_40_O),
    .config_addr(config_reg_40_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_41_config_addr;
assign config_reg_41_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_26_8_32_41 config_reg_41 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_41_O),
    .config_addr(config_reg_41_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_42_config_addr;
assign config_reg_42_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_27_8_32_42 config_reg_42 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_42_O),
    .config_addr(config_reg_42_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_43_config_addr;
assign config_reg_43_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_27_8_32_43 config_reg_43 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_43_O),
    .config_addr(config_reg_43_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_44_config_addr;
assign config_reg_44_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_27_8_32_44 config_reg_44 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_44_O),
    .config_addr(config_reg_44_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_45_config_addr;
assign config_reg_45_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_27_8_32_45 config_reg_45 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_45_O),
    .config_addr(config_reg_45_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_46_config_addr;
assign config_reg_46_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_27_8_32_46 config_reg_46 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_46_O),
    .config_addr(config_reg_46_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_47_config_addr;
assign config_reg_47_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_27_8_32_47 config_reg_47 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_47_O),
    .config_addr(config_reg_47_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_48_config_addr;
assign config_reg_48_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_27_8_32_48 config_reg_48 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_48_O),
    .config_addr(config_reg_48_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_49_config_addr;
assign config_reg_49_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_27_8_32_49 config_reg_49 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_49_O),
    .config_addr(config_reg_49_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_5_config_addr;
assign config_reg_5_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_5 config_reg_5 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_5_O),
    .config_addr(config_reg_5_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_50_config_addr;
assign config_reg_50_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_31_8_32_50 config_reg_50 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_50_O),
    .config_addr(config_reg_50_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_51_config_addr;
assign config_reg_51_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_51 config_reg_51 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_51_O),
    .config_addr(config_reg_51_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_52_config_addr;
assign config_reg_52_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_52 config_reg_52 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_52_O),
    .config_addr(config_reg_52_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_53_config_addr;
assign config_reg_53_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_53 config_reg_53 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_53_O),
    .config_addr(config_reg_53_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_54_config_addr;
assign config_reg_54_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_20_8_32_54 config_reg_54 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_54_O),
    .config_addr(config_reg_54_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_55_config_addr;
assign config_reg_55_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_55 config_reg_55 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_55_O),
    .config_addr(config_reg_55_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_56_config_addr;
assign config_reg_56_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_56 config_reg_56 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_56_O),
    .config_addr(config_reg_56_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_57_config_addr;
assign config_reg_57_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_17_8_32_57 config_reg_57 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_57_O),
    .config_addr(config_reg_57_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_58_config_addr;
assign config_reg_58_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_58 config_reg_58 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_58_O),
    .config_addr(config_reg_58_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_59_config_addr;
assign config_reg_59_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_59 config_reg_59 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_59_O),
    .config_addr(config_reg_59_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_6_config_addr;
assign config_reg_6_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_6 config_reg_6 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_6_O),
    .config_addr(config_reg_6_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_60_config_addr;
assign config_reg_60_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_60 config_reg_60 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_60_O),
    .config_addr(config_reg_60_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_61_config_addr;
assign config_reg_61_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_17_8_32_61 config_reg_61 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_61_O),
    .config_addr(config_reg_61_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_62_config_addr;
assign config_reg_62_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_62 config_reg_62 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_62_O),
    .config_addr(config_reg_62_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_63_config_addr;
assign config_reg_63_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_63 config_reg_63 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_63_O),
    .config_addr(config_reg_63_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_64_config_addr;
assign config_reg_64_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_64 config_reg_64 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_64_O),
    .config_addr(config_reg_64_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_65_config_addr;
assign config_reg_65_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_20_8_32_65 config_reg_65 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_65_O),
    .config_addr(config_reg_65_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_66_config_addr;
assign config_reg_66_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_66 config_reg_66 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_66_O),
    .config_addr(config_reg_66_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_67_config_addr;
assign config_reg_67_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_67 config_reg_67 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_67_O),
    .config_addr(config_reg_67_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_68_config_addr;
assign config_reg_68_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_68 config_reg_68 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_68_O),
    .config_addr(config_reg_68_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_69_config_addr;
assign config_reg_69_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_20_8_32_69 config_reg_69 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_69_O),
    .config_addr(config_reg_69_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_7_config_addr;
assign config_reg_7_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_7 config_reg_7 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_7_O),
    .config_addr(config_reg_7_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_70_config_addr;
assign config_reg_70_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_70 config_reg_70 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_70_O),
    .config_addr(config_reg_70_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_71_config_addr;
assign config_reg_71_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_71 config_reg_71 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_71_O),
    .config_addr(config_reg_71_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_72_config_addr;
assign config_reg_72_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_72 config_reg_72 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_72_O),
    .config_addr(config_reg_72_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_73_config_addr;
assign config_reg_73_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_73 config_reg_73 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_73_O),
    .config_addr(config_reg_73_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_74_config_addr;
assign config_reg_74_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_25_8_32_74 config_reg_74 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_74_O),
    .config_addr(config_reg_74_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_75_config_addr;
assign config_reg_75_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_75 config_reg_75 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_75_O),
    .config_addr(config_reg_75_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_76_config_addr;
assign config_reg_76_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_76 config_reg_76 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_76_O),
    .config_addr(config_reg_76_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_77_config_addr;
assign config_reg_77_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_77 config_reg_77 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_77_O),
    .config_addr(config_reg_77_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_78_config_addr;
assign config_reg_78_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_17_8_32_78 config_reg_78 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_78_O),
    .config_addr(config_reg_78_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_79_config_addr;
assign config_reg_79_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_79 config_reg_79 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_79_O),
    .config_addr(config_reg_79_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_8_config_addr;
assign config_reg_8_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_8 config_reg_8 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_8_O),
    .config_addr(config_reg_8_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_80_config_addr;
assign config_reg_80_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_80 config_reg_80 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_80_O),
    .config_addr(config_reg_80_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_81_config_addr;
assign config_reg_81_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_81 config_reg_81 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_81_O),
    .config_addr(config_reg_81_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_82_config_addr;
assign config_reg_82_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_82 config_reg_82 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_82_O),
    .config_addr(config_reg_82_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_83_config_addr;
assign config_reg_83_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_27_8_32_83 config_reg_83 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_83_O),
    .config_addr(config_reg_83_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_9_config_addr;
assign config_reg_9_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6:0]};
ConfigRegister_32_8_32_9 config_reg_9 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_9_O),
    .config_addr(config_reg_9_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_wrap coreir_wrapInAsyncReset_inst0 (
    .in(reset),
    .out(coreir_wrapInAsyncReset_inst0_out)
);
coreir_wrap coreir_wrapOutAsyncReset_inst0 (
    .in(Invert1_inst0_out[0]),
    .out(coreir_wrapOutAsyncReset_inst0_out)
);
coreir_mux #(
    .width(1)
) flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(flush_core),
    .in1(flush),
    .sel(flush_mux_sel_inst0_O[0]),
    .out(flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
flush_mux_sel_unq1 flush_mux_sel_inst0 (
    .I(config_reg_0_O),
    .O(flush_mux_sel_inst0_O)
);
input_width_1_num_0_reg_sel input_width_1_num_0_reg_sel_inst0 (
    .I(config_reg_0_O),
    .O(input_width_1_num_0_reg_sel_inst0_O)
);
input_width_1_num_0_reg_value input_width_1_num_0_reg_value_inst0 (
    .I(config_reg_0_O),
    .O(input_width_1_num_0_reg_value_inst0_O)
);
coreir_mux #(
    .width(1)
) input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(input_width_1_num_0),
    .in1(input_width_1_num_0_reg_value_inst0_O),
    .sel(input_width_1_num_0_reg_sel_inst0_O[0]),
    .out(input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
input_width_1_num_1_reg_sel input_width_1_num_1_reg_sel_inst0 (
    .I(config_reg_0_O),
    .O(input_width_1_num_1_reg_sel_inst0_O)
);
input_width_1_num_1_reg_value input_width_1_num_1_reg_value_inst0 (
    .I(config_reg_0_O),
    .O(input_width_1_num_1_reg_value_inst0_O)
);
coreir_mux #(
    .width(1)
) input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(input_width_1_num_1),
    .in1(input_width_1_num_1_reg_value_inst0_O),
    .sel(input_width_1_num_1_reg_sel_inst0_O[0]),
    .out(input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality_inst0 (
    .I(config_reg_0_O),
    .O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality_inst0_O)
);
mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0 mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0_inst0 (
    .I(config_reg_0_O),
    .O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0_inst0_O)
);
mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1 mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1_inst0 (
    .I(config_reg_1_O),
    .O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1_inst0_O)
);
mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2 mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2_inst0 (
    .I(config_reg_1_O),
    .O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2_inst0_O)
);
mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3 mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3_inst0 (
    .I(config_reg_2_O),
    .O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3_inst0_O)
);
mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4 mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4_inst0 (
    .I(config_reg_2_O),
    .O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4_inst0_O)
);
mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5 mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5_inst0 (
    .I(config_reg_3_O),
    .O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5_inst0_O)
);
mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable_inst0 (
    .I(config_reg_3_O),
    .O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable_inst0_O)
);
mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_4_O),
    .O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr_inst0_O)
);
mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0 mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_4_O),
    .O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0_inst0_O)
);
mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1 mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_5_O),
    .O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1_inst0_O)
);
mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2 mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_5_O),
    .O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2_inst0_O)
);
mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3 mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3_inst0 (
    .I(config_reg_6_O),
    .O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3_inst0_O)
);
mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4 mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4_inst0 (
    .I(config_reg_6_O),
    .O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4_inst0_O)
);
mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5 mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5_inst0 (
    .I(config_reg_7_O),
    .O(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5_inst0_O)
);
mem_ctrl_strg_fifo_flat_strg_fifo_inst_fifo_depth mem_ctrl_strg_fifo_flat_strg_fifo_inst_fifo_depth_inst0 (
    .I(config_reg_7_O),
    .O(mem_ctrl_strg_fifo_flat_strg_fifo_inst_fifo_depth_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr_inst0 (
    .I(config_reg_8_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0_inst0 (
    .I(config_reg_8_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1_inst0 (
    .I(config_reg_8_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2_inst0 (
    .I(config_reg_8_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3_inst0 (
    .I(config_reg_8_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4_inst0 (
    .I(config_reg_8_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5_inst0 (
    .I(config_reg_8_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_0_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr_inst0 (
    .I(config_reg_8_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0_inst0 (
    .I(config_reg_9_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1_inst0 (
    .I(config_reg_9_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2_inst0 (
    .I(config_reg_9_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3_inst0 (
    .I(config_reg_9_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4_inst0 (
    .I(config_reg_9_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5_inst0 (
    .I(config_reg_9_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_read_addr_gen_1_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr_inst0 (
    .I(config_reg_9_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0_inst0 (
    .I(config_reg_9_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1_inst0 (
    .I(config_reg_10_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2_inst0 (
    .I(config_reg_10_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3_inst0 (
    .I(config_reg_10_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4_inst0 (
    .I(config_reg_10_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5_inst0 (
    .I(config_reg_10_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr_inst0 (
    .I(config_reg_10_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0_inst0 (
    .I(config_reg_10_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1_inst0 (
    .I(config_reg_10_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2_inst0 (
    .I(config_reg_11_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3_inst0 (
    .I(config_reg_11_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4_inst0 (
    .I(config_reg_11_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5_inst0 (
    .I(config_reg_11_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable_inst0 (
    .I(config_reg_11_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_12_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_12_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_13_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_13_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3_inst0 (
    .I(config_reg_14_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4_inst0 (
    .I(config_reg_14_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5_inst0 (
    .I(config_reg_15_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable_inst0 (
    .I(config_reg_15_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_16_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_16_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_17_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_17_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3_inst0 (
    .I(config_reg_18_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4_inst0 (
    .I(config_reg_18_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5_inst0 (
    .I(config_reg_19_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality_inst0 (
    .I(config_reg_19_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0_inst0 (
    .I(config_reg_20_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1_inst0 (
    .I(config_reg_20_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2_inst0 (
    .I(config_reg_21_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3_inst0 (
    .I(config_reg_21_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4_inst0 (
    .I(config_reg_22_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5_inst0 (
    .I(config_reg_22_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality_inst0 (
    .I(config_reg_23_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0_inst0 (
    .I(config_reg_23_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1_inst0 (
    .I(config_reg_24_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2_inst0 (
    .I(config_reg_24_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3_inst0 (
    .I(config_reg_25_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4_inst0 (
    .I(config_reg_25_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5_inst0 (
    .I(config_reg_26_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable_inst0 (
    .I(config_reg_26_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_enable_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_27_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_27_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_28_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_28_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3_inst0 (
    .I(config_reg_29_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4_inst0 (
    .I(config_reg_29_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5_inst0 (
    .I(config_reg_30_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable_inst0 (
    .I(config_reg_30_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_enable_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_31_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_31_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_32_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_32_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3_inst0 (
    .I(config_reg_33_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4_inst0 (
    .I(config_reg_33_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5_inst0 (
    .I(config_reg_34_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality_inst0 (
    .I(config_reg_34_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0_inst0 (
    .I(config_reg_35_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1_inst0 (
    .I(config_reg_35_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2_inst0 (
    .I(config_reg_36_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3_inst0 (
    .I(config_reg_36_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4_inst0 (
    .I(config_reg_37_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5_inst0 (
    .I(config_reg_37_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality_inst0 (
    .I(config_reg_38_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0_inst0 (
    .I(config_reg_38_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1_inst0 (
    .I(config_reg_39_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2_inst0 (
    .I(config_reg_39_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3_inst0 (
    .I(config_reg_40_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4_inst0 (
    .I(config_reg_40_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5_inst0 (
    .I(config_reg_41_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en_inst0 (
    .I(config_reg_41_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr_inst0 (
    .I(config_reg_41_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0_inst0 (
    .I(config_reg_42_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1_inst0 (
    .I(config_reg_42_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2_inst0 (
    .I(config_reg_42_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3_inst0 (
    .I(config_reg_43_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4_inst0 (
    .I(config_reg_43_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5_inst0 (
    .I(config_reg_43_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_0_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr_inst0 (
    .I(config_reg_44_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0_inst0 (
    .I(config_reg_44_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1_inst0 (
    .I(config_reg_44_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2_inst0 (
    .I(config_reg_45_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3_inst0 (
    .I(config_reg_45_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4_inst0 (
    .I(config_reg_45_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5_inst0 (
    .I(config_reg_46_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_input_addr_gen_1_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr_inst0 (
    .I(config_reg_46_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0_inst0 (
    .I(config_reg_46_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1_inst0 (
    .I(config_reg_47_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2_inst0 (
    .I(config_reg_47_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3_inst0 (
    .I(config_reg_47_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4_inst0 (
    .I(config_reg_48_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5_inst0 (
    .I(config_reg_48_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr_inst0 (
    .I(config_reg_48_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0_inst0 (
    .I(config_reg_49_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1_inst0 (
    .I(config_reg_49_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2_inst0 (
    .I(config_reg_49_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3_inst0 (
    .I(config_reg_50_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4_inst0 (
    .I(config_reg_50_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5_inst0 (
    .I(config_reg_50_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality_inst0 (
    .I(config_reg_50_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0_inst0 (
    .I(config_reg_51_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1_inst0 (
    .I(config_reg_51_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2_inst0 (
    .I(config_reg_52_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3_inst0 (
    .I(config_reg_52_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4_inst0 (
    .I(config_reg_53_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5_inst0 (
    .I(config_reg_53_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality_inst0 (
    .I(config_reg_54_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0_inst0 (
    .I(config_reg_54_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1_inst0 (
    .I(config_reg_55_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2_inst0 (
    .I(config_reg_55_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3_inst0 (
    .I(config_reg_56_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4_inst0 (
    .I(config_reg_56_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5_inst0 (
    .I(config_reg_57_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable_inst0 (
    .I(config_reg_57_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_58_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_58_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_59_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_59_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3_inst0 (
    .I(config_reg_60_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4_inst0 (
    .I(config_reg_60_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5_inst0 (
    .I(config_reg_61_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable_inst0 (
    .I(config_reg_61_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_62_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_62_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_63_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_63_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3_inst0 (
    .I(config_reg_64_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4_inst0 (
    .I(config_reg_64_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5_inst0 (
    .I(config_reg_65_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality_inst0 (
    .I(config_reg_65_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0_inst0 (
    .I(config_reg_66_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1_inst0 (
    .I(config_reg_66_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2_inst0 (
    .I(config_reg_67_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3_inst0 (
    .I(config_reg_67_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4_inst0 (
    .I(config_reg_68_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5_inst0 (
    .I(config_reg_68_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality_inst0 (
    .I(config_reg_69_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0_inst0 (
    .I(config_reg_69_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1_inst0 (
    .I(config_reg_70_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2_inst0 (
    .I(config_reg_70_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3_inst0 (
    .I(config_reg_71_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4_inst0 (
    .I(config_reg_71_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5_inst0 (
    .I(config_reg_72_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr_inst0 (
    .I(config_reg_72_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0_inst0 (
    .I(config_reg_72_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1_inst0 (
    .I(config_reg_72_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2_inst0 (
    .I(config_reg_72_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3_inst0 (
    .I(config_reg_73_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4_inst0 (
    .I(config_reg_73_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5_inst0 (
    .I(config_reg_73_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr_inst0 (
    .I(config_reg_73_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0_inst0 (
    .I(config_reg_73_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1_inst0 (
    .I(config_reg_73_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2_inst0 (
    .I(config_reg_73_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3_inst0 (
    .I(config_reg_73_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4_inst0 (
    .I(config_reg_74_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5_inst0 (
    .I(config_reg_74_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable_inst0 (
    .I(config_reg_74_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_74_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_75_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_75_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_76_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3_inst0 (
    .I(config_reg_76_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4_inst0 (
    .I(config_reg_77_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5_inst0 (
    .I(config_reg_77_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable_inst0 (
    .I(config_reg_78_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_78_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_79_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_79_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_80_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3_inst0 (
    .I(config_reg_80_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4_inst0 (
    .I(config_reg_81_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5_inst0 (
    .I(config_reg_81_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr_inst0 (
    .I(config_reg_82_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0_inst0 (
    .I(config_reg_82_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1_inst0 (
    .I(config_reg_82_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2_inst0 (
    .I(config_reg_82_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3_inst0 (
    .I(config_reg_82_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4_inst0 (
    .I(config_reg_82_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5_inst0 (
    .I(config_reg_82_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr_inst0 (
    .I(config_reg_82_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0_inst0 (
    .I(config_reg_83_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1_inst0 (
    .I(config_reg_83_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2_inst0 (
    .I(config_reg_83_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3_inst0 (
    .I(config_reg_83_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4_inst0 (
    .I(config_reg_83_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4_inst0_O)
);
mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5 mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5_inst0 (
    .I(config_reg_83_O),
    .O(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5_inst0_O)
);
mode mode_inst0 (
    .I(config_reg_83_O),
    .O(mode_inst0_O)
);
mantle_wire__typeBit8 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
tile_en_unq1 tile_en_inst0 (
    .I(config_reg_83_O),
    .O(tile_en_inst0_O)
);
assign output_width_16_num_0 = LakeTop_W_inst0_output_width_16_num_0;
assign output_width_16_num_1 = LakeTop_W_inst0_output_width_16_num_1;
assign output_width_1_num_0 = LakeTop_W_inst0_output_width_1_num_0;
assign output_width_1_num_1 = LakeTop_W_inst0_output_width_1_num_1;
assign output_width_1_num_2 = LakeTop_W_inst0_output_width_1_num_2;
assign output_width_1_num_3 = LakeTop_W_inst0_output_width_1_num_3;
assign read_config_data = MuxWrapper_84_32_inst0$Mux84xBits32_inst0$coreir_commonlib_mux84x32_inst0_out;
assign read_config_data_1 = LakeTop_W_inst0_config_data_out_0;
assign read_config_data_2 = LakeTop_W_inst0_config_data_out_1;
endmodule

module Cond (
    input [4:0] code,
    input alu,
    input Z,
    input N,
    input C,
    input V,
    output O,
    input CLK,
    input ASYNCRESET
);
wire [0:0] Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst13$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst14$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst15$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst16$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst17$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst9$coreir_commonlib_mux2x1_inst0$_join_out;
wire [4:0] const_0_5_out;
wire [4:0] const_10_5_out;
wire [4:0] const_11_5_out;
wire [4:0] const_12_5_out;
wire [4:0] const_13_5_out;
wire [4:0] const_14_5_out;
wire [4:0] const_15_5_out;
wire [4:0] const_16_5_out;
wire [4:0] const_17_5_out;
wire [4:0] const_1_5_out;
wire [4:0] const_2_5_out;
wire [4:0] const_3_5_out;
wire [4:0] const_4_5_out;
wire [4:0] const_5_5_out;
wire [4:0] const_6_5_out;
wire [4:0] const_7_5_out;
wire [4:0] const_8_5_out;
wire [4:0] const_9_5_out;
wire magma_Bit_and_inst0_out;
wire magma_Bit_and_inst1_out;
wire magma_Bit_and_inst2_out;
wire magma_Bit_and_inst3_out;
wire magma_Bit_not_inst0_out;
wire magma_Bit_not_inst1_out;
wire magma_Bit_not_inst10_out;
wire magma_Bit_not_inst11_out;
wire magma_Bit_not_inst12_out;
wire magma_Bit_not_inst2_out;
wire magma_Bit_not_inst3_out;
wire magma_Bit_not_inst4_out;
wire magma_Bit_not_inst5_out;
wire magma_Bit_not_inst6_out;
wire magma_Bit_not_inst7_out;
wire magma_Bit_not_inst8_out;
wire magma_Bit_not_inst9_out;
wire magma_Bit_or_inst0_out;
wire magma_Bit_or_inst1_out;
wire magma_Bit_or_inst2_out;
wire magma_Bit_or_inst3_out;
wire magma_Bit_or_inst4_out;
wire magma_Bit_or_inst5_out;
wire magma_Bit_xor_inst0_out;
wire magma_Bit_xor_inst1_out;
wire magma_Bit_xor_inst2_out;
wire magma_Bit_xor_inst3_out;
wire magma_Bits_5_eq_inst0_out;
wire magma_Bits_5_eq_inst1_out;
wire magma_Bits_5_eq_inst10_out;
wire magma_Bits_5_eq_inst11_out;
wire magma_Bits_5_eq_inst12_out;
wire magma_Bits_5_eq_inst13_out;
wire magma_Bits_5_eq_inst14_out;
wire magma_Bits_5_eq_inst15_out;
wire magma_Bits_5_eq_inst16_out;
wire magma_Bits_5_eq_inst17_out;
wire magma_Bits_5_eq_inst18_out;
wire magma_Bits_5_eq_inst19_out;
wire magma_Bits_5_eq_inst2_out;
wire magma_Bits_5_eq_inst3_out;
wire magma_Bits_5_eq_inst4_out;
wire magma_Bits_5_eq_inst5_out;
wire magma_Bits_5_eq_inst6_out;
wire magma_Bits_5_eq_inst7_out;
wire magma_Bits_5_eq_inst8_out;
wire magma_Bits_5_eq_inst9_out;
coreir_mux #(
    .width(1)
) Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(magma_Bit_and_inst3_out),
    .in1(magma_Bit_or_inst5_out),
    .sel(magma_Bits_5_eq_inst19_out),
    .out(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_and_inst2_out),
    .sel(magma_Bits_5_eq_inst18_out),
    .out(Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst10$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst9$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_not_inst3_out),
    .sel(magma_Bits_5_eq_inst9_out),
    .out(Mux2xBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst11$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(V),
    .sel(magma_Bits_5_eq_inst8_out),
    .out(Mux2xBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst12$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_not_inst2_out),
    .sel(magma_Bits_5_eq_inst7_out),
    .out(Mux2xBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst13$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(N),
    .sel(magma_Bits_5_eq_inst6_out),
    .out(Mux2xBit_inst13$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst14$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst13$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_not_inst1_out),
    .sel(magma_Bit_or_inst1_out),
    .out(Mux2xBit_inst14$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst15$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst14$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(C),
    .sel(magma_Bit_or_inst0_out),
    .out(Mux2xBit_inst15$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst16$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst15$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_not_inst0_out),
    .sel(magma_Bits_5_eq_inst1_out),
    .out(Mux2xBit_inst16$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst17$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst16$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(Z),
    .sel(magma_Bits_5_eq_inst0_out),
    .out(Mux2xBit_inst17$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_or_inst4_out),
    .sel(magma_Bits_5_eq_inst17_out),
    .out(Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(alu),
    .sel(magma_Bits_5_eq_inst16_out),
    .out(Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_or_inst3_out),
    .sel(magma_Bits_5_eq_inst15_out),
    .out(Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_and_inst1_out),
    .sel(magma_Bits_5_eq_inst14_out),
    .out(Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_xor_inst1_out),
    .sel(magma_Bits_5_eq_inst13_out),
    .out(Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_not_inst6_out),
    .sel(magma_Bits_5_eq_inst12_out),
    .out(Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst8$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_or_inst2_out),
    .sel(magma_Bits_5_eq_inst11_out),
    .out(Mux2xBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst9$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_and_inst0_out),
    .sel(magma_Bits_5_eq_inst10_out),
    .out(Mux2xBit_inst9$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_const #(
    .value(5'h00),
    .width(5)
) const_0_5 (
    .out(const_0_5_out)
);
coreir_const #(
    .value(5'h0a),
    .width(5)
) const_10_5 (
    .out(const_10_5_out)
);
coreir_const #(
    .value(5'h0b),
    .width(5)
) const_11_5 (
    .out(const_11_5_out)
);
coreir_const #(
    .value(5'h0c),
    .width(5)
) const_12_5 (
    .out(const_12_5_out)
);
coreir_const #(
    .value(5'h0d),
    .width(5)
) const_13_5 (
    .out(const_13_5_out)
);
coreir_const #(
    .value(5'h0e),
    .width(5)
) const_14_5 (
    .out(const_14_5_out)
);
coreir_const #(
    .value(5'h0f),
    .width(5)
) const_15_5 (
    .out(const_15_5_out)
);
coreir_const #(
    .value(5'h10),
    .width(5)
) const_16_5 (
    .out(const_16_5_out)
);
coreir_const #(
    .value(5'h11),
    .width(5)
) const_17_5 (
    .out(const_17_5_out)
);
coreir_const #(
    .value(5'h01),
    .width(5)
) const_1_5 (
    .out(const_1_5_out)
);
coreir_const #(
    .value(5'h02),
    .width(5)
) const_2_5 (
    .out(const_2_5_out)
);
coreir_const #(
    .value(5'h03),
    .width(5)
) const_3_5 (
    .out(const_3_5_out)
);
coreir_const #(
    .value(5'h04),
    .width(5)
) const_4_5 (
    .out(const_4_5_out)
);
coreir_const #(
    .value(5'h05),
    .width(5)
) const_5_5 (
    .out(const_5_5_out)
);
coreir_const #(
    .value(5'h06),
    .width(5)
) const_6_5 (
    .out(const_6_5_out)
);
coreir_const #(
    .value(5'h07),
    .width(5)
) const_7_5 (
    .out(const_7_5_out)
);
coreir_const #(
    .value(5'h08),
    .width(5)
) const_8_5 (
    .out(const_8_5_out)
);
coreir_const #(
    .value(5'h09),
    .width(5)
) const_9_5 (
    .out(const_9_5_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(C),
    .in1(magma_Bit_not_inst4_out),
    .out(magma_Bit_and_inst0_out)
);
corebit_and magma_Bit_and_inst1 (
    .in0(magma_Bit_not_inst7_out),
    .in1(magma_Bit_not_inst8_out),
    .out(magma_Bit_and_inst1_out)
);
corebit_and magma_Bit_and_inst2 (
    .in0(magma_Bit_not_inst10_out),
    .in1(magma_Bit_not_inst11_out),
    .out(magma_Bit_and_inst2_out)
);
corebit_and magma_Bit_and_inst3 (
    .in0(N),
    .in1(magma_Bit_not_inst12_out),
    .out(magma_Bit_and_inst3_out)
);
corebit_not magma_Bit_not_inst0 (
    .in(Z),
    .out(magma_Bit_not_inst0_out)
);
corebit_not magma_Bit_not_inst1 (
    .in(C),
    .out(magma_Bit_not_inst1_out)
);
corebit_not magma_Bit_not_inst10 (
    .in(N),
    .out(magma_Bit_not_inst10_out)
);
corebit_not magma_Bit_not_inst11 (
    .in(Z),
    .out(magma_Bit_not_inst11_out)
);
corebit_not magma_Bit_not_inst12 (
    .in(Z),
    .out(magma_Bit_not_inst12_out)
);
corebit_not magma_Bit_not_inst2 (
    .in(N),
    .out(magma_Bit_not_inst2_out)
);
corebit_not magma_Bit_not_inst3 (
    .in(V),
    .out(magma_Bit_not_inst3_out)
);
corebit_not magma_Bit_not_inst4 (
    .in(Z),
    .out(magma_Bit_not_inst4_out)
);
corebit_not magma_Bit_not_inst5 (
    .in(C),
    .out(magma_Bit_not_inst5_out)
);
corebit_not magma_Bit_not_inst6 (
    .in(magma_Bit_xor_inst0_out),
    .out(magma_Bit_not_inst6_out)
);
corebit_not magma_Bit_not_inst7 (
    .in(Z),
    .out(magma_Bit_not_inst7_out)
);
corebit_not magma_Bit_not_inst8 (
    .in(magma_Bit_xor_inst2_out),
    .out(magma_Bit_not_inst8_out)
);
corebit_not magma_Bit_not_inst9 (
    .in(N),
    .out(magma_Bit_not_inst9_out)
);
corebit_or magma_Bit_or_inst0 (
    .in0(magma_Bits_5_eq_inst2_out),
    .in1(magma_Bits_5_eq_inst3_out),
    .out(magma_Bit_or_inst0_out)
);
corebit_or magma_Bit_or_inst1 (
    .in0(magma_Bits_5_eq_inst4_out),
    .in1(magma_Bits_5_eq_inst5_out),
    .out(magma_Bit_or_inst1_out)
);
corebit_or magma_Bit_or_inst2 (
    .in0(magma_Bit_not_inst5_out),
    .in1(Z),
    .out(magma_Bit_or_inst2_out)
);
corebit_or magma_Bit_or_inst3 (
    .in0(Z),
    .in1(magma_Bit_xor_inst3_out),
    .out(magma_Bit_or_inst3_out)
);
corebit_or magma_Bit_or_inst4 (
    .in0(magma_Bit_not_inst9_out),
    .in1(Z),
    .out(magma_Bit_or_inst4_out)
);
corebit_or magma_Bit_or_inst5 (
    .in0(N),
    .in1(Z),
    .out(magma_Bit_or_inst5_out)
);
corebit_xor magma_Bit_xor_inst0 (
    .in0(N),
    .in1(V),
    .out(magma_Bit_xor_inst0_out)
);
corebit_xor magma_Bit_xor_inst1 (
    .in0(N),
    .in1(V),
    .out(magma_Bit_xor_inst1_out)
);
corebit_xor magma_Bit_xor_inst2 (
    .in0(N),
    .in1(V),
    .out(magma_Bit_xor_inst2_out)
);
corebit_xor magma_Bit_xor_inst3 (
    .in0(N),
    .in1(V),
    .out(magma_Bit_xor_inst3_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst0 (
    .in0(code),
    .in1(const_0_5_out),
    .out(magma_Bits_5_eq_inst0_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst1 (
    .in0(code),
    .in1(const_1_5_out),
    .out(magma_Bits_5_eq_inst1_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst10 (
    .in0(code),
    .in1(const_8_5_out),
    .out(magma_Bits_5_eq_inst10_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst11 (
    .in0(code),
    .in1(const_9_5_out),
    .out(magma_Bits_5_eq_inst11_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst12 (
    .in0(code),
    .in1(const_10_5_out),
    .out(magma_Bits_5_eq_inst12_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst13 (
    .in0(code),
    .in1(const_11_5_out),
    .out(magma_Bits_5_eq_inst13_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst14 (
    .in0(code),
    .in1(const_12_5_out),
    .out(magma_Bits_5_eq_inst14_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst15 (
    .in0(code),
    .in1(const_13_5_out),
    .out(magma_Bits_5_eq_inst15_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst16 (
    .in0(code),
    .in1(const_14_5_out),
    .out(magma_Bits_5_eq_inst16_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst17 (
    .in0(code),
    .in1(const_15_5_out),
    .out(magma_Bits_5_eq_inst17_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst18 (
    .in0(code),
    .in1(const_16_5_out),
    .out(magma_Bits_5_eq_inst18_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst19 (
    .in0(code),
    .in1(const_17_5_out),
    .out(magma_Bits_5_eq_inst19_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst2 (
    .in0(code),
    .in1(const_2_5_out),
    .out(magma_Bits_5_eq_inst2_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst3 (
    .in0(code),
    .in1(const_2_5_out),
    .out(magma_Bits_5_eq_inst3_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst4 (
    .in0(code),
    .in1(const_3_5_out),
    .out(magma_Bits_5_eq_inst4_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst5 (
    .in0(code),
    .in1(const_3_5_out),
    .out(magma_Bits_5_eq_inst5_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst6 (
    .in0(code),
    .in1(const_4_5_out),
    .out(magma_Bits_5_eq_inst6_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst7 (
    .in0(code),
    .in1(const_5_5_out),
    .out(magma_Bits_5_eq_inst7_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst8 (
    .in0(code),
    .in1(const_6_5_out),
    .out(magma_Bits_5_eq_inst8_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst9 (
    .in0(code),
    .in1(const_7_5_out),
    .out(magma_Bits_5_eq_inst9_out)
);
assign O = Mux2xBit_inst17$coreir_commonlib_mux2x1_inst0$_join_out[0];
endmodule

module CB_inputs6_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_inputs6 (
    input [0:0] I_0,
    input [0:0] I_1,
    input [0:0] I_10,
    input [0:0] I_11,
    input [0:0] I_12,
    input [0:0] I_13,
    input [0:0] I_14,
    input [0:0] I_15,
    input [0:0] I_16,
    input [0:0] I_17,
    input [0:0] I_18,
    input [0:0] I_19,
    input [0:0] I_2,
    input [0:0] I_3,
    input [0:0] I_4,
    input [0:0] I_5,
    input [0:0] I_6,
    input [0:0] I_7,
    input [0:0] I_8,
    input [0:0] I_9,
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [0:0] CB_inputs6_O;
wire [4:0] CB_inputs6_sel_inst0_O;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
MuxWrapperAOIImpl_20_1 CB_inputs6 (
    .I_0(I_0),
    .I_1(I_1),
    .I_10(I_10),
    .I_11(I_11),
    .I_12(I_12),
    .I_13(I_13),
    .I_14(I_14),
    .I_15(I_15),
    .I_16(I_16),
    .I_17(I_17),
    .I_18(I_18),
    .I_19(I_19),
    .I_2(I_2),
    .I_3(I_3),
    .I_4(I_4),
    .I_5(I_5),
    .I_6(I_6),
    .I_7(I_7),
    .I_8(I_8),
    .I_9(I_9),
    .O(CB_inputs6_O),
    .S(CB_inputs6_sel_inst0_O)
);
CB_inputs6_sel CB_inputs6_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_inputs6_sel_inst0_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_inputs6_O;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_inputs5_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_inputs5 (
    input [0:0] I_0,
    input [0:0] I_1,
    input [0:0] I_10,
    input [0:0] I_11,
    input [0:0] I_12,
    input [0:0] I_13,
    input [0:0] I_14,
    input [0:0] I_15,
    input [0:0] I_16,
    input [0:0] I_17,
    input [0:0] I_18,
    input [0:0] I_19,
    input [0:0] I_2,
    input [0:0] I_3,
    input [0:0] I_4,
    input [0:0] I_5,
    input [0:0] I_6,
    input [0:0] I_7,
    input [0:0] I_8,
    input [0:0] I_9,
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [0:0] CB_inputs5_O;
wire [4:0] CB_inputs5_sel_inst0_O;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
MuxWrapperAOIImpl_20_1 CB_inputs5 (
    .I_0(I_0),
    .I_1(I_1),
    .I_10(I_10),
    .I_11(I_11),
    .I_12(I_12),
    .I_13(I_13),
    .I_14(I_14),
    .I_15(I_15),
    .I_16(I_16),
    .I_17(I_17),
    .I_18(I_18),
    .I_19(I_19),
    .I_2(I_2),
    .I_3(I_3),
    .I_4(I_4),
    .I_5(I_5),
    .I_6(I_6),
    .I_7(I_7),
    .I_8(I_8),
    .I_9(I_9),
    .O(CB_inputs5_O),
    .S(CB_inputs5_sel_inst0_O)
);
CB_inputs5_sel CB_inputs5_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_inputs5_sel_inst0_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_inputs5_O;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_inputs4_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_inputs4 (
    input [0:0] I_0,
    input [0:0] I_1,
    input [0:0] I_10,
    input [0:0] I_11,
    input [0:0] I_12,
    input [0:0] I_13,
    input [0:0] I_14,
    input [0:0] I_15,
    input [0:0] I_16,
    input [0:0] I_17,
    input [0:0] I_18,
    input [0:0] I_19,
    input [0:0] I_2,
    input [0:0] I_3,
    input [0:0] I_4,
    input [0:0] I_5,
    input [0:0] I_6,
    input [0:0] I_7,
    input [0:0] I_8,
    input [0:0] I_9,
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [0:0] CB_inputs4_O;
wire [4:0] CB_inputs4_sel_inst0_O;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
MuxWrapperAOIImpl_20_1 CB_inputs4 (
    .I_0(I_0),
    .I_1(I_1),
    .I_10(I_10),
    .I_11(I_11),
    .I_12(I_12),
    .I_13(I_13),
    .I_14(I_14),
    .I_15(I_15),
    .I_16(I_16),
    .I_17(I_17),
    .I_18(I_18),
    .I_19(I_19),
    .I_2(I_2),
    .I_3(I_3),
    .I_4(I_4),
    .I_5(I_5),
    .I_6(I_6),
    .I_7(I_7),
    .I_8(I_8),
    .I_9(I_9),
    .O(CB_inputs4_O),
    .S(CB_inputs4_sel_inst0_O)
);
CB_inputs4_sel CB_inputs4_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_inputs4_sel_inst0_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_inputs4_O;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_inputs3_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_inputs3 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [15:0] CB_inputs3_O;
wire [4:0] CB_inputs3_sel_inst0_O;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
MuxWrapperAOIImpl_20_16 CB_inputs3 (
    .I_0(I_0),
    .I_1(I_1),
    .I_10(I_10),
    .I_11(I_11),
    .I_12(I_12),
    .I_13(I_13),
    .I_14(I_14),
    .I_15(I_15),
    .I_16(I_16),
    .I_17(I_17),
    .I_18(I_18),
    .I_19(I_19),
    .I_2(I_2),
    .I_3(I_3),
    .I_4(I_4),
    .I_5(I_5),
    .I_6(I_6),
    .I_7(I_7),
    .I_8(I_8),
    .I_9(I_9),
    .O(CB_inputs3_O),
    .S(CB_inputs3_sel_inst0_O)
);
CB_inputs3_sel CB_inputs3_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_inputs3_sel_inst0_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_inputs3_O;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_inputs2_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_inputs2 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [15:0] CB_inputs2_O;
wire [4:0] CB_inputs2_sel_inst0_O;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
MuxWrapperAOIImpl_20_16 CB_inputs2 (
    .I_0(I_0),
    .I_1(I_1),
    .I_10(I_10),
    .I_11(I_11),
    .I_12(I_12),
    .I_13(I_13),
    .I_14(I_14),
    .I_15(I_15),
    .I_16(I_16),
    .I_17(I_17),
    .I_18(I_18),
    .I_19(I_19),
    .I_2(I_2),
    .I_3(I_3),
    .I_4(I_4),
    .I_5(I_5),
    .I_6(I_6),
    .I_7(I_7),
    .I_8(I_8),
    .I_9(I_9),
    .O(CB_inputs2_O),
    .S(CB_inputs2_sel_inst0_O)
);
CB_inputs2_sel CB_inputs2_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_inputs2_sel_inst0_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_inputs2_O;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_inputs1_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_inputs1 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [15:0] CB_inputs1_O;
wire [4:0] CB_inputs1_sel_inst0_O;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
MuxWrapperAOIImpl_20_16 CB_inputs1 (
    .I_0(I_0),
    .I_1(I_1),
    .I_10(I_10),
    .I_11(I_11),
    .I_12(I_12),
    .I_13(I_13),
    .I_14(I_14),
    .I_15(I_15),
    .I_16(I_16),
    .I_17(I_17),
    .I_18(I_18),
    .I_19(I_19),
    .I_2(I_2),
    .I_3(I_3),
    .I_4(I_4),
    .I_5(I_5),
    .I_6(I_6),
    .I_7(I_7),
    .I_8(I_8),
    .I_9(I_9),
    .O(CB_inputs1_O),
    .S(CB_inputs1_sel_inst0_O)
);
CB_inputs1_sel CB_inputs1_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_inputs1_sel_inst0_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_inputs1_O;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_inputs0_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_inputs0 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [15:0] CB_inputs0_O;
wire [4:0] CB_inputs0_sel_inst0_O;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
MuxWrapperAOIImpl_20_16 CB_inputs0 (
    .I_0(I_0),
    .I_1(I_1),
    .I_10(I_10),
    .I_11(I_11),
    .I_12(I_12),
    .I_13(I_13),
    .I_14(I_14),
    .I_15(I_15),
    .I_16(I_16),
    .I_17(I_17),
    .I_18(I_18),
    .I_19(I_19),
    .I_2(I_2),
    .I_3(I_3),
    .I_4(I_4),
    .I_5(I_5),
    .I_6(I_6),
    .I_7(I_7),
    .I_8(I_8),
    .I_9(I_9),
    .O(CB_inputs0_O),
    .S(CB_inputs0_sel_inst0_O)
);
CB_inputs0_sel CB_inputs0_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_inputs0_sel_inst0_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_inputs0_O;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_input_width_1_num_1_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_input_width_1_num_1 (
    input [0:0] I_0,
    input [0:0] I_1,
    input [0:0] I_10,
    input [0:0] I_11,
    input [0:0] I_12,
    input [0:0] I_13,
    input [0:0] I_14,
    input [0:0] I_15,
    input [0:0] I_16,
    input [0:0] I_17,
    input [0:0] I_18,
    input [0:0] I_19,
    input [0:0] I_2,
    input [0:0] I_3,
    input [0:0] I_4,
    input [0:0] I_5,
    input [0:0] I_6,
    input [0:0] I_7,
    input [0:0] I_8,
    input [0:0] I_9,
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [0:0] CB_input_width_1_num_1_O;
wire [4:0] CB_input_width_1_num_1_sel_inst0_O;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
MuxWrapperAOIImpl_20_1 CB_input_width_1_num_1 (
    .I_0(I_0),
    .I_1(I_1),
    .I_10(I_10),
    .I_11(I_11),
    .I_12(I_12),
    .I_13(I_13),
    .I_14(I_14),
    .I_15(I_15),
    .I_16(I_16),
    .I_17(I_17),
    .I_18(I_18),
    .I_19(I_19),
    .I_2(I_2),
    .I_3(I_3),
    .I_4(I_4),
    .I_5(I_5),
    .I_6(I_6),
    .I_7(I_7),
    .I_8(I_8),
    .I_9(I_9),
    .O(CB_input_width_1_num_1_O),
    .S(CB_input_width_1_num_1_sel_inst0_O)
);
CB_input_width_1_num_1_sel CB_input_width_1_num_1_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_input_width_1_num_1_sel_inst0_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_input_width_1_num_1_O;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_input_width_1_num_0_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_input_width_1_num_0 (
    input [0:0] I_0,
    input [0:0] I_1,
    input [0:0] I_10,
    input [0:0] I_11,
    input [0:0] I_12,
    input [0:0] I_13,
    input [0:0] I_14,
    input [0:0] I_15,
    input [0:0] I_16,
    input [0:0] I_17,
    input [0:0] I_18,
    input [0:0] I_19,
    input [0:0] I_2,
    input [0:0] I_3,
    input [0:0] I_4,
    input [0:0] I_5,
    input [0:0] I_6,
    input [0:0] I_7,
    input [0:0] I_8,
    input [0:0] I_9,
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [0:0] CB_input_width_1_num_0_O;
wire [4:0] CB_input_width_1_num_0_sel_inst0_O;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
MuxWrapperAOIImpl_20_1 CB_input_width_1_num_0 (
    .I_0(I_0),
    .I_1(I_1),
    .I_10(I_10),
    .I_11(I_11),
    .I_12(I_12),
    .I_13(I_13),
    .I_14(I_14),
    .I_15(I_15),
    .I_16(I_16),
    .I_17(I_17),
    .I_18(I_18),
    .I_19(I_19),
    .I_2(I_2),
    .I_3(I_3),
    .I_4(I_4),
    .I_5(I_5),
    .I_6(I_6),
    .I_7(I_7),
    .I_8(I_8),
    .I_9(I_9),
    .O(CB_input_width_1_num_0_O),
    .S(CB_input_width_1_num_0_sel_inst0_O)
);
CB_input_width_1_num_0_sel CB_input_width_1_num_0_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_input_width_1_num_0_sel_inst0_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_input_width_1_num_0_O;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_input_width_16_num_3_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_input_width_16_num_3 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [15:0] CB_input_width_16_num_3_O;
wire [4:0] CB_input_width_16_num_3_sel_inst0_O;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
MuxWrapperAOIImpl_20_16 CB_input_width_16_num_3 (
    .I_0(I_0),
    .I_1(I_1),
    .I_10(I_10),
    .I_11(I_11),
    .I_12(I_12),
    .I_13(I_13),
    .I_14(I_14),
    .I_15(I_15),
    .I_16(I_16),
    .I_17(I_17),
    .I_18(I_18),
    .I_19(I_19),
    .I_2(I_2),
    .I_3(I_3),
    .I_4(I_4),
    .I_5(I_5),
    .I_6(I_6),
    .I_7(I_7),
    .I_8(I_8),
    .I_9(I_9),
    .O(CB_input_width_16_num_3_O),
    .S(CB_input_width_16_num_3_sel_inst0_O)
);
CB_input_width_16_num_3_sel CB_input_width_16_num_3_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_input_width_16_num_3_sel_inst0_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_input_width_16_num_3_O;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_input_width_16_num_2_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_input_width_16_num_2 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [15:0] CB_input_width_16_num_2_O;
wire [4:0] CB_input_width_16_num_2_sel_inst0_O;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
MuxWrapperAOIImpl_20_16 CB_input_width_16_num_2 (
    .I_0(I_0),
    .I_1(I_1),
    .I_10(I_10),
    .I_11(I_11),
    .I_12(I_12),
    .I_13(I_13),
    .I_14(I_14),
    .I_15(I_15),
    .I_16(I_16),
    .I_17(I_17),
    .I_18(I_18),
    .I_19(I_19),
    .I_2(I_2),
    .I_3(I_3),
    .I_4(I_4),
    .I_5(I_5),
    .I_6(I_6),
    .I_7(I_7),
    .I_8(I_8),
    .I_9(I_9),
    .O(CB_input_width_16_num_2_O),
    .S(CB_input_width_16_num_2_sel_inst0_O)
);
CB_input_width_16_num_2_sel CB_input_width_16_num_2_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_input_width_16_num_2_sel_inst0_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_input_width_16_num_2_O;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_input_width_16_num_1_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_input_width_16_num_1 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [15:0] CB_input_width_16_num_1_O;
wire [4:0] CB_input_width_16_num_1_sel_inst0_O;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
MuxWrapperAOIImpl_20_16 CB_input_width_16_num_1 (
    .I_0(I_0),
    .I_1(I_1),
    .I_10(I_10),
    .I_11(I_11),
    .I_12(I_12),
    .I_13(I_13),
    .I_14(I_14),
    .I_15(I_15),
    .I_16(I_16),
    .I_17(I_17),
    .I_18(I_18),
    .I_19(I_19),
    .I_2(I_2),
    .I_3(I_3),
    .I_4(I_4),
    .I_5(I_5),
    .I_6(I_6),
    .I_7(I_7),
    .I_8(I_8),
    .I_9(I_9),
    .O(CB_input_width_16_num_1_O),
    .S(CB_input_width_16_num_1_sel_inst0_O)
);
CB_input_width_16_num_1_sel CB_input_width_16_num_1_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_input_width_16_num_1_sel_inst0_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_input_width_16_num_1_O;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_input_width_16_num_0_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_input_width_16_num_0 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [15:0] CB_input_width_16_num_0_O;
wire [4:0] CB_input_width_16_num_0_sel_inst0_O;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
MuxWrapperAOIImpl_20_16 CB_input_width_16_num_0 (
    .I_0(I_0),
    .I_1(I_1),
    .I_10(I_10),
    .I_11(I_11),
    .I_12(I_12),
    .I_13(I_13),
    .I_14(I_14),
    .I_15(I_15),
    .I_16(I_16),
    .I_17(I_17),
    .I_18(I_18),
    .I_19(I_19),
    .I_2(I_2),
    .I_3(I_3),
    .I_4(I_4),
    .I_5(I_5),
    .I_6(I_6),
    .I_7(I_7),
    .I_8(I_8),
    .I_9(I_9),
    .O(CB_input_width_16_num_0_O),
    .S(CB_input_width_16_num_0_sel_inst0_O)
);
CB_input_width_16_num_0_sel CB_input_width_16_num_0_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_input_width_16_num_0_sel_inst0_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_input_width_16_num_0_O;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_flush_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_flush (
    input [0:0] I_0,
    input [0:0] I_1,
    input [0:0] I_10,
    input [0:0] I_11,
    input [0:0] I_12,
    input [0:0] I_13,
    input [0:0] I_14,
    input [0:0] I_15,
    input [0:0] I_16,
    input [0:0] I_17,
    input [0:0] I_18,
    input [0:0] I_19,
    input [0:0] I_2,
    input [0:0] I_3,
    input [0:0] I_4,
    input [0:0] I_5,
    input [0:0] I_6,
    input [0:0] I_7,
    input [0:0] I_8,
    input [0:0] I_9,
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [0:0] CB_flush_O;
wire [4:0] CB_flush_sel_inst0_O;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
MuxWrapperAOIImpl_20_1 CB_flush (
    .I_0(I_0),
    .I_1(I_1),
    .I_10(I_10),
    .I_11(I_11),
    .I_12(I_12),
    .I_13(I_13),
    .I_14(I_14),
    .I_15(I_15),
    .I_16(I_16),
    .I_17(I_17),
    .I_18(I_18),
    .I_19(I_19),
    .I_2(I_2),
    .I_3(I_3),
    .I_4(I_4),
    .I_5(I_5),
    .I_6(I_6),
    .I_7(I_7),
    .I_8(I_8),
    .I_9(I_9),
    .O(CB_flush_O),
    .S(CB_flush_sel_inst0_O)
);
CB_flush_sel CB_flush_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_flush_sel_inst0_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_flush_O;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module Tile_MemCore (
    input [0:0] SB_T0_EAST_SB_IN_B1,
    input [15:0] SB_T0_EAST_SB_IN_B16,
    output [0:0] SB_T0_EAST_SB_OUT_B1,
    output [15:0] SB_T0_EAST_SB_OUT_B16,
    input [0:0] SB_T0_NORTH_SB_IN_B1,
    input [15:0] SB_T0_NORTH_SB_IN_B16,
    output [0:0] SB_T0_NORTH_SB_OUT_B1,
    output [15:0] SB_T0_NORTH_SB_OUT_B16,
    input [0:0] SB_T0_SOUTH_SB_IN_B1,
    input [15:0] SB_T0_SOUTH_SB_IN_B16,
    output [0:0] SB_T0_SOUTH_SB_OUT_B1,
    output [15:0] SB_T0_SOUTH_SB_OUT_B16,
    input [0:0] SB_T0_WEST_SB_IN_B1,
    input [15:0] SB_T0_WEST_SB_IN_B16,
    output [0:0] SB_T0_WEST_SB_OUT_B1,
    output [15:0] SB_T0_WEST_SB_OUT_B16,
    input [0:0] SB_T1_EAST_SB_IN_B1,
    input [15:0] SB_T1_EAST_SB_IN_B16,
    output [0:0] SB_T1_EAST_SB_OUT_B1,
    output [15:0] SB_T1_EAST_SB_OUT_B16,
    input [0:0] SB_T1_NORTH_SB_IN_B1,
    input [15:0] SB_T1_NORTH_SB_IN_B16,
    output [0:0] SB_T1_NORTH_SB_OUT_B1,
    output [15:0] SB_T1_NORTH_SB_OUT_B16,
    input [0:0] SB_T1_SOUTH_SB_IN_B1,
    input [15:0] SB_T1_SOUTH_SB_IN_B16,
    output [0:0] SB_T1_SOUTH_SB_OUT_B1,
    output [15:0] SB_T1_SOUTH_SB_OUT_B16,
    input [0:0] SB_T1_WEST_SB_IN_B1,
    input [15:0] SB_T1_WEST_SB_IN_B16,
    output [0:0] SB_T1_WEST_SB_OUT_B1,
    output [15:0] SB_T1_WEST_SB_OUT_B16,
    input [0:0] SB_T2_EAST_SB_IN_B1,
    input [15:0] SB_T2_EAST_SB_IN_B16,
    output [0:0] SB_T2_EAST_SB_OUT_B1,
    output [15:0] SB_T2_EAST_SB_OUT_B16,
    input [0:0] SB_T2_NORTH_SB_IN_B1,
    input [15:0] SB_T2_NORTH_SB_IN_B16,
    output [0:0] SB_T2_NORTH_SB_OUT_B1,
    output [15:0] SB_T2_NORTH_SB_OUT_B16,
    input [0:0] SB_T2_SOUTH_SB_IN_B1,
    input [15:0] SB_T2_SOUTH_SB_IN_B16,
    output [0:0] SB_T2_SOUTH_SB_OUT_B1,
    output [15:0] SB_T2_SOUTH_SB_OUT_B16,
    input [0:0] SB_T2_WEST_SB_IN_B1,
    input [15:0] SB_T2_WEST_SB_IN_B16,
    output [0:0] SB_T2_WEST_SB_OUT_B1,
    output [15:0] SB_T2_WEST_SB_OUT_B16,
    input [0:0] SB_T3_EAST_SB_IN_B1,
    input [15:0] SB_T3_EAST_SB_IN_B16,
    output [0:0] SB_T3_EAST_SB_OUT_B1,
    output [15:0] SB_T3_EAST_SB_OUT_B16,
    input [0:0] SB_T3_NORTH_SB_IN_B1,
    input [15:0] SB_T3_NORTH_SB_IN_B16,
    output [0:0] SB_T3_NORTH_SB_OUT_B1,
    output [15:0] SB_T3_NORTH_SB_OUT_B16,
    input [0:0] SB_T3_SOUTH_SB_IN_B1,
    input [15:0] SB_T3_SOUTH_SB_IN_B16,
    output [0:0] SB_T3_SOUTH_SB_OUT_B1,
    output [15:0] SB_T3_SOUTH_SB_OUT_B16,
    input [0:0] SB_T3_WEST_SB_IN_B1,
    input [15:0] SB_T3_WEST_SB_IN_B16,
    output [0:0] SB_T3_WEST_SB_OUT_B1,
    output [15:0] SB_T3_WEST_SB_OUT_B16,
    input [0:0] SB_T4_EAST_SB_IN_B1,
    input [15:0] SB_T4_EAST_SB_IN_B16,
    output [0:0] SB_T4_EAST_SB_OUT_B1,
    output [15:0] SB_T4_EAST_SB_OUT_B16,
    input [0:0] SB_T4_NORTH_SB_IN_B1,
    input [15:0] SB_T4_NORTH_SB_IN_B16,
    output [0:0] SB_T4_NORTH_SB_OUT_B1,
    output [15:0] SB_T4_NORTH_SB_OUT_B16,
    input [0:0] SB_T4_SOUTH_SB_IN_B1,
    input [15:0] SB_T4_SOUTH_SB_IN_B16,
    output [0:0] SB_T4_SOUTH_SB_OUT_B1,
    output [15:0] SB_T4_SOUTH_SB_OUT_B16,
    input [0:0] SB_T4_WEST_SB_IN_B1,
    input [15:0] SB_T4_WEST_SB_IN_B16,
    output [0:0] SB_T4_WEST_SB_OUT_B1,
    output [15:0] SB_T4_WEST_SB_OUT_B16,
    input clk,
    output clk_out,
    input [31:0] config_config_addr,
    input [31:0] config_config_data,
    output [31:0] config_out_config_addr,
    output [31:0] config_out_config_data,
    output [0:0] config_out_read,
    output [0:0] config_out_write,
    input [0:0] config_read,
    input [0:0] config_write,
    input [0:0] flush,
    output [0:0] flush_out,
    output [8:0] hi,
    output [7:0] lo,
    output [31:0] read_config_data,
    input [31:0] read_config_data_in,
    input reset,
    output reset_out,
    input [0:0] stall,
    output [0:0] stall_out,
    input [15:0] tile_id
);
wire [0:0] CB_flush_O;
wire [31:0] CB_flush_read_config_data;
wire [15:0] CB_input_width_16_num_0_O;
wire [31:0] CB_input_width_16_num_0_read_config_data;
wire [15:0] CB_input_width_16_num_1_O;
wire [31:0] CB_input_width_16_num_1_read_config_data;
wire [15:0] CB_input_width_16_num_2_O;
wire [31:0] CB_input_width_16_num_2_read_config_data;
wire [15:0] CB_input_width_16_num_3_O;
wire [31:0] CB_input_width_16_num_3_read_config_data;
wire [0:0] CB_input_width_1_num_0_O;
wire [31:0] CB_input_width_1_num_0_read_config_data;
wire [0:0] CB_input_width_1_num_1_O;
wire [31:0] CB_input_width_1_num_1_read_config_data;
wire DECODE_FEATURE_0_O;
wire DECODE_FEATURE_1_O;
wire DECODE_FEATURE_10_O;
wire DECODE_FEATURE_11_O;
wire DECODE_FEATURE_12_O;
wire DECODE_FEATURE_2_O;
wire DECODE_FEATURE_3_O;
wire DECODE_FEATURE_4_O;
wire DECODE_FEATURE_5_O;
wire DECODE_FEATURE_6_O;
wire DECODE_FEATURE_7_O;
wire DECODE_FEATURE_8_O;
wire DECODE_FEATURE_9_O;
wire FEATURE_AND_0_out;
wire FEATURE_AND_1_out;
wire FEATURE_AND_10_out;
wire FEATURE_AND_11_out;
wire FEATURE_AND_12_out;
wire FEATURE_AND_2_out;
wire FEATURE_AND_3_out;
wire FEATURE_AND_4_out;
wire FEATURE_AND_5_out;
wire FEATURE_AND_6_out;
wire FEATURE_AND_7_out;
wire FEATURE_AND_8_out;
wire FEATURE_AND_9_out;
wire [15:0] MemCore_inst0_output_width_16_num_0;
wire [15:0] MemCore_inst0_output_width_16_num_1;
wire [0:0] MemCore_inst0_output_width_1_num_0;
wire [0:0] MemCore_inst0_output_width_1_num_1;
wire [0:0] MemCore_inst0_output_width_1_num_2;
wire [0:0] MemCore_inst0_output_width_1_num_3;
wire [31:0] MemCore_inst0_read_config_data;
wire [31:0] MemCore_inst0_read_config_data_1;
wire [31:0] MemCore_inst0_read_config_data_2;
wire [0:0] PowerDomainConfigReg_inst0_ps_en_out;
wire [31:0] PowerDomainConfigReg_inst0_read_config_data;
wire [31:0] PowerDomainOR_O;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T0_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T0_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T0_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T0_WEST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T1_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T1_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T1_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T1_WEST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T2_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T2_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T2_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T2_WEST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T3_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T3_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T3_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T3_WEST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T4_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T4_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T4_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T4_WEST_SB_OUT_B16;
wire [31:0] SB_ID0_5TRACKS_B16_MemCore_read_config_data;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1;
wire [31:0] SB_ID0_5TRACKS_B1_MemCore_read_config_data;
wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T3_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T3_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T3_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T3_WEST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T4_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T4_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T4_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T4_WEST_SB_IN_B16_O;
wire and_inst0_out;
wire and_inst1_out;
wire [7:0] const_0_8_out;
wire [8:0] const_511_9_out;
wire coreir_eq_16_inst0_out;
wire [31:0] read_data_mux_O;
wire [7:0] CB_flush_config_config_addr;
assign CB_flush_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
CB_flush CB_flush (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .O(CB_flush_O),
    .clk(clk),
    .config_config_addr(CB_flush_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_3_out),
    .read_config_data(CB_flush_read_config_data),
    .reset(reset)
);
wire [7:0] CB_input_width_16_num_0_config_config_addr;
assign CB_input_width_16_num_0_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
CB_input_width_16_num_0 CB_input_width_16_num_0 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .O(CB_input_width_16_num_0_O),
    .clk(clk),
    .config_config_addr(CB_input_width_16_num_0_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_4_out),
    .read_config_data(CB_input_width_16_num_0_read_config_data),
    .reset(reset)
);
wire [7:0] CB_input_width_16_num_1_config_config_addr;
assign CB_input_width_16_num_1_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
CB_input_width_16_num_1 CB_input_width_16_num_1 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .O(CB_input_width_16_num_1_O),
    .clk(clk),
    .config_config_addr(CB_input_width_16_num_1_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_5_out),
    .read_config_data(CB_input_width_16_num_1_read_config_data),
    .reset(reset)
);
wire [7:0] CB_input_width_16_num_2_config_config_addr;
assign CB_input_width_16_num_2_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
CB_input_width_16_num_2 CB_input_width_16_num_2 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .O(CB_input_width_16_num_2_O),
    .clk(clk),
    .config_config_addr(CB_input_width_16_num_2_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_6_out),
    .read_config_data(CB_input_width_16_num_2_read_config_data),
    .reset(reset)
);
wire [7:0] CB_input_width_16_num_3_config_config_addr;
assign CB_input_width_16_num_3_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
CB_input_width_16_num_3 CB_input_width_16_num_3 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .O(CB_input_width_16_num_3_O),
    .clk(clk),
    .config_config_addr(CB_input_width_16_num_3_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_7_out),
    .read_config_data(CB_input_width_16_num_3_read_config_data),
    .reset(reset)
);
wire [7:0] CB_input_width_1_num_0_config_config_addr;
assign CB_input_width_1_num_0_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
CB_input_width_1_num_0 CB_input_width_1_num_0 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .O(CB_input_width_1_num_0_O),
    .clk(clk),
    .config_config_addr(CB_input_width_1_num_0_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_8_out),
    .read_config_data(CB_input_width_1_num_0_read_config_data),
    .reset(reset)
);
wire [7:0] CB_input_width_1_num_1_config_config_addr;
assign CB_input_width_1_num_1_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
CB_input_width_1_num_1 CB_input_width_1_num_1 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .O(CB_input_width_1_num_1_O),
    .clk(clk),
    .config_config_addr(CB_input_width_1_num_1_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_9_out),
    .read_config_data(CB_input_width_1_num_1_read_config_data),
    .reset(reset)
);
wire [7:0] DECODE_FEATURE_0_I;
assign DECODE_FEATURE_0_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode08 DECODE_FEATURE_0 (
    .I(DECODE_FEATURE_0_I),
    .O(DECODE_FEATURE_0_O)
);
wire [7:0] DECODE_FEATURE_1_I;
assign DECODE_FEATURE_1_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode18 DECODE_FEATURE_1 (
    .I(DECODE_FEATURE_1_I),
    .O(DECODE_FEATURE_1_O)
);
wire [7:0] DECODE_FEATURE_10_I;
assign DECODE_FEATURE_10_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode108 DECODE_FEATURE_10 (
    .I(DECODE_FEATURE_10_I),
    .O(DECODE_FEATURE_10_O)
);
wire [7:0] DECODE_FEATURE_11_I;
assign DECODE_FEATURE_11_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode118 DECODE_FEATURE_11 (
    .I(DECODE_FEATURE_11_I),
    .O(DECODE_FEATURE_11_O)
);
wire [7:0] DECODE_FEATURE_12_I;
assign DECODE_FEATURE_12_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode128 DECODE_FEATURE_12 (
    .I(DECODE_FEATURE_12_I),
    .O(DECODE_FEATURE_12_O)
);
wire [7:0] DECODE_FEATURE_2_I;
assign DECODE_FEATURE_2_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode28 DECODE_FEATURE_2 (
    .I(DECODE_FEATURE_2_I),
    .O(DECODE_FEATURE_2_O)
);
wire [7:0] DECODE_FEATURE_3_I;
assign DECODE_FEATURE_3_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode38 DECODE_FEATURE_3 (
    .I(DECODE_FEATURE_3_I),
    .O(DECODE_FEATURE_3_O)
);
wire [7:0] DECODE_FEATURE_4_I;
assign DECODE_FEATURE_4_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode48 DECODE_FEATURE_4 (
    .I(DECODE_FEATURE_4_I),
    .O(DECODE_FEATURE_4_O)
);
wire [7:0] DECODE_FEATURE_5_I;
assign DECODE_FEATURE_5_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode58 DECODE_FEATURE_5 (
    .I(DECODE_FEATURE_5_I),
    .O(DECODE_FEATURE_5_O)
);
wire [7:0] DECODE_FEATURE_6_I;
assign DECODE_FEATURE_6_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode68 DECODE_FEATURE_6 (
    .I(DECODE_FEATURE_6_I),
    .O(DECODE_FEATURE_6_O)
);
wire [7:0] DECODE_FEATURE_7_I;
assign DECODE_FEATURE_7_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode78 DECODE_FEATURE_7 (
    .I(DECODE_FEATURE_7_I),
    .O(DECODE_FEATURE_7_O)
);
wire [7:0] DECODE_FEATURE_8_I;
assign DECODE_FEATURE_8_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode88 DECODE_FEATURE_8 (
    .I(DECODE_FEATURE_8_I),
    .O(DECODE_FEATURE_8_O)
);
wire [7:0] DECODE_FEATURE_9_I;
assign DECODE_FEATURE_9_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode98 DECODE_FEATURE_9 (
    .I(DECODE_FEATURE_9_I),
    .O(DECODE_FEATURE_9_O)
);
corebit_and FEATURE_AND_0 (
    .in0(DECODE_FEATURE_0_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_0_out)
);
corebit_and FEATURE_AND_1 (
    .in0(DECODE_FEATURE_1_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_1_out)
);
corebit_and FEATURE_AND_10 (
    .in0(DECODE_FEATURE_10_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_10_out)
);
corebit_and FEATURE_AND_11 (
    .in0(DECODE_FEATURE_11_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_11_out)
);
corebit_and FEATURE_AND_12 (
    .in0(DECODE_FEATURE_12_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_12_out)
);
corebit_and FEATURE_AND_2 (
    .in0(DECODE_FEATURE_2_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_2_out)
);
corebit_and FEATURE_AND_3 (
    .in0(DECODE_FEATURE_3_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_3_out)
);
corebit_and FEATURE_AND_4 (
    .in0(DECODE_FEATURE_4_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_4_out)
);
corebit_and FEATURE_AND_5 (
    .in0(DECODE_FEATURE_5_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_5_out)
);
corebit_and FEATURE_AND_6 (
    .in0(DECODE_FEATURE_6_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_6_out)
);
corebit_and FEATURE_AND_7 (
    .in0(DECODE_FEATURE_7_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_7_out)
);
corebit_and FEATURE_AND_8 (
    .in0(DECODE_FEATURE_8_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_8_out)
);
corebit_and FEATURE_AND_9 (
    .in0(DECODE_FEATURE_9_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_9_out)
);
wire [7:0] MemCore_inst0_config_1_config_addr;
assign MemCore_inst0_config_1_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
wire [7:0] MemCore_inst0_config_2_config_addr;
assign MemCore_inst0_config_2_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
wire [7:0] MemCore_inst0_config_config_addr;
assign MemCore_inst0_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
MemCore MemCore_inst0 (
    .clk(clk),
    .config_1_config_addr(MemCore_inst0_config_1_config_addr),
    .config_1_config_data(config_config_data),
    .config_1_read(config_read),
    .config_1_write(FEATURE_AND_1_out),
    .config_2_config_addr(MemCore_inst0_config_2_config_addr),
    .config_2_config_data(config_config_data),
    .config_2_read(config_read),
    .config_2_write(FEATURE_AND_2_out),
    .config_config_addr(MemCore_inst0_config_config_addr),
    .config_config_data(config_config_data),
    .config_en_0(DECODE_FEATURE_1_O),
    .config_en_1(DECODE_FEATURE_2_O),
    .config_read(config_read),
    .config_write(FEATURE_AND_0_out),
    .flush(CB_flush_O),
    .flush_core(flush),
    .input_width_16_num_0(CB_input_width_16_num_0_O),
    .input_width_16_num_1(CB_input_width_16_num_1_O),
    .input_width_16_num_2(CB_input_width_16_num_2_O),
    .input_width_16_num_3(CB_input_width_16_num_3_O),
    .input_width_1_num_0(CB_input_width_1_num_0_O),
    .input_width_1_num_1(CB_input_width_1_num_1_O),
    .output_width_16_num_0(MemCore_inst0_output_width_16_num_0),
    .output_width_16_num_1(MemCore_inst0_output_width_16_num_1),
    .output_width_1_num_0(MemCore_inst0_output_width_1_num_0),
    .output_width_1_num_1(MemCore_inst0_output_width_1_num_1),
    .output_width_1_num_2(MemCore_inst0_output_width_1_num_2),
    .output_width_1_num_3(MemCore_inst0_output_width_1_num_3),
    .read_config_data(MemCore_inst0_read_config_data),
    .read_config_data_1(MemCore_inst0_read_config_data_1),
    .read_config_data_2(MemCore_inst0_read_config_data_2),
    .reset(reset),
    .stall(stall)
);
wire [7:0] PowerDomainConfigReg_inst0_config_config_addr;
assign PowerDomainConfigReg_inst0_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
PowerDomainConfigReg PowerDomainConfigReg_inst0 (
    .clk(clk),
    .config_config_addr(PowerDomainConfigReg_inst0_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_12_out),
    .ps_en_out(PowerDomainConfigReg_inst0_ps_en_out),
    .read_config_data(PowerDomainConfigReg_inst0_read_config_data),
    .reset(reset)
);
PowerDomainOR PowerDomainOR (
    .I0(read_data_mux_O),
    .I1(read_config_data_in),
    .O(PowerDomainOR_O),
    .I_not(PowerDomainConfigReg_inst0_ps_en_out)
);
wire [7:0] SB_ID0_5TRACKS_B16_MemCore_config_config_addr;
assign SB_ID0_5TRACKS_B16_MemCore_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
SB_ID0_5TRACKS_B16_MemCore SB_ID0_5TRACKS_B16_MemCore (
    .SB_T0_EAST_SB_IN_B16(SB_T0_EAST_SB_IN_B16),
    .SB_T0_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B16(SB_T0_NORTH_SB_IN_B16),
    .SB_T0_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B16(SB_T0_SOUTH_SB_IN_B16),
    .SB_T0_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B16(SB_T0_WEST_SB_IN_B16),
    .SB_T0_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B16(SB_T1_EAST_SB_IN_B16),
    .SB_T1_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B16(SB_T1_NORTH_SB_IN_B16),
    .SB_T1_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B16(SB_T1_SOUTH_SB_IN_B16),
    .SB_T1_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B16(SB_T1_WEST_SB_IN_B16),
    .SB_T1_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B16(SB_T2_EAST_SB_IN_B16),
    .SB_T2_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B16(SB_T2_NORTH_SB_IN_B16),
    .SB_T2_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B16(SB_T2_SOUTH_SB_IN_B16),
    .SB_T2_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B16(SB_T2_WEST_SB_IN_B16),
    .SB_T2_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B16(SB_T3_EAST_SB_IN_B16),
    .SB_T3_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B16(SB_T3_NORTH_SB_IN_B16),
    .SB_T3_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B16(SB_T3_SOUTH_SB_IN_B16),
    .SB_T3_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B16(SB_T3_WEST_SB_IN_B16),
    .SB_T3_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B16(SB_T4_EAST_SB_IN_B16),
    .SB_T4_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B16(SB_T4_NORTH_SB_IN_B16),
    .SB_T4_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B16(SB_T4_SOUTH_SB_IN_B16),
    .SB_T4_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B16(SB_T4_WEST_SB_IN_B16),
    .SB_T4_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .config_config_addr(SB_ID0_5TRACKS_B16_MemCore_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_11_out),
    .output_width_16_num_0(MemCore_inst0_output_width_16_num_0),
    .output_width_16_num_1(MemCore_inst0_output_width_16_num_1),
    .read_config_data(SB_ID0_5TRACKS_B16_MemCore_read_config_data),
    .reset(reset),
    .stall(stall)
);
wire [7:0] SB_ID0_5TRACKS_B1_MemCore_config_config_addr;
assign SB_ID0_5TRACKS_B1_MemCore_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
SB_ID0_5TRACKS_B1_MemCore SB_ID0_5TRACKS_B1_MemCore (
    .SB_T0_EAST_SB_IN_B1(SB_T0_EAST_SB_IN_B1),
    .SB_T0_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B1(SB_T0_NORTH_SB_IN_B1),
    .SB_T0_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B1(SB_T0_SOUTH_SB_IN_B1),
    .SB_T0_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B1(SB_T0_WEST_SB_IN_B1),
    .SB_T0_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B1(SB_T1_EAST_SB_IN_B1),
    .SB_T1_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B1(SB_T1_NORTH_SB_IN_B1),
    .SB_T1_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B1(SB_T1_SOUTH_SB_IN_B1),
    .SB_T1_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B1(SB_T1_WEST_SB_IN_B1),
    .SB_T1_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B1(SB_T2_EAST_SB_IN_B1),
    .SB_T2_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B1(SB_T2_NORTH_SB_IN_B1),
    .SB_T2_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B1(SB_T2_SOUTH_SB_IN_B1),
    .SB_T2_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B1(SB_T2_WEST_SB_IN_B1),
    .SB_T2_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B1(SB_T3_EAST_SB_IN_B1),
    .SB_T3_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B1(SB_T3_NORTH_SB_IN_B1),
    .SB_T3_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B1(SB_T3_SOUTH_SB_IN_B1),
    .SB_T3_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B1(SB_T3_WEST_SB_IN_B1),
    .SB_T3_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B1(SB_T4_EAST_SB_IN_B1),
    .SB_T4_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B1(SB_T4_NORTH_SB_IN_B1),
    .SB_T4_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B1(SB_T4_SOUTH_SB_IN_B1),
    .SB_T4_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B1(SB_T4_WEST_SB_IN_B1),
    .SB_T4_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1),
    .clk(clk),
    .config_config_addr(SB_ID0_5TRACKS_B1_MemCore_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_10_out),
    .output_width_1_num_0(MemCore_inst0_output_width_1_num_0),
    .output_width_1_num_1(MemCore_inst0_output_width_1_num_1),
    .output_width_1_num_2(MemCore_inst0_output_width_1_num_2),
    .output_width_1_num_3(MemCore_inst0_output_width_1_num_3),
    .read_config_data(SB_ID0_5TRACKS_B1_MemCore_read_config_data),
    .reset(reset),
    .stall(stall)
);
MuxWrapper_1_1 WIRE_SB_T0_EAST_SB_IN_B1 (
    .I(SB_T0_EAST_SB_IN_B1),
    .O(WIRE_SB_T0_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T0_EAST_SB_IN_B16 (
    .I(SB_T0_EAST_SB_IN_B16),
    .O(WIRE_SB_T0_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T0_NORTH_SB_IN_B1 (
    .I(SB_T0_NORTH_SB_IN_B1),
    .O(WIRE_SB_T0_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T0_NORTH_SB_IN_B16 (
    .I(SB_T0_NORTH_SB_IN_B16),
    .O(WIRE_SB_T0_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T0_SOUTH_SB_IN_B1 (
    .I(SB_T0_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T0_SOUTH_SB_IN_B16 (
    .I(SB_T0_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T0_WEST_SB_IN_B1 (
    .I(SB_T0_WEST_SB_IN_B1),
    .O(WIRE_SB_T0_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T0_WEST_SB_IN_B16 (
    .I(SB_T0_WEST_SB_IN_B16),
    .O(WIRE_SB_T0_WEST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T1_EAST_SB_IN_B1 (
    .I(SB_T1_EAST_SB_IN_B1),
    .O(WIRE_SB_T1_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T1_EAST_SB_IN_B16 (
    .I(SB_T1_EAST_SB_IN_B16),
    .O(WIRE_SB_T1_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T1_NORTH_SB_IN_B1 (
    .I(SB_T1_NORTH_SB_IN_B1),
    .O(WIRE_SB_T1_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T1_NORTH_SB_IN_B16 (
    .I(SB_T1_NORTH_SB_IN_B16),
    .O(WIRE_SB_T1_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T1_SOUTH_SB_IN_B1 (
    .I(SB_T1_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T1_SOUTH_SB_IN_B16 (
    .I(SB_T1_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T1_WEST_SB_IN_B1 (
    .I(SB_T1_WEST_SB_IN_B1),
    .O(WIRE_SB_T1_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T1_WEST_SB_IN_B16 (
    .I(SB_T1_WEST_SB_IN_B16),
    .O(WIRE_SB_T1_WEST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T2_EAST_SB_IN_B1 (
    .I(SB_T2_EAST_SB_IN_B1),
    .O(WIRE_SB_T2_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T2_EAST_SB_IN_B16 (
    .I(SB_T2_EAST_SB_IN_B16),
    .O(WIRE_SB_T2_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T2_NORTH_SB_IN_B1 (
    .I(SB_T2_NORTH_SB_IN_B1),
    .O(WIRE_SB_T2_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T2_NORTH_SB_IN_B16 (
    .I(SB_T2_NORTH_SB_IN_B16),
    .O(WIRE_SB_T2_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T2_SOUTH_SB_IN_B1 (
    .I(SB_T2_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T2_SOUTH_SB_IN_B16 (
    .I(SB_T2_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T2_WEST_SB_IN_B1 (
    .I(SB_T2_WEST_SB_IN_B1),
    .O(WIRE_SB_T2_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T2_WEST_SB_IN_B16 (
    .I(SB_T2_WEST_SB_IN_B16),
    .O(WIRE_SB_T2_WEST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T3_EAST_SB_IN_B1 (
    .I(SB_T3_EAST_SB_IN_B1),
    .O(WIRE_SB_T3_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T3_EAST_SB_IN_B16 (
    .I(SB_T3_EAST_SB_IN_B16),
    .O(WIRE_SB_T3_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T3_NORTH_SB_IN_B1 (
    .I(SB_T3_NORTH_SB_IN_B1),
    .O(WIRE_SB_T3_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T3_NORTH_SB_IN_B16 (
    .I(SB_T3_NORTH_SB_IN_B16),
    .O(WIRE_SB_T3_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T3_SOUTH_SB_IN_B1 (
    .I(SB_T3_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T3_SOUTH_SB_IN_B16 (
    .I(SB_T3_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T3_WEST_SB_IN_B1 (
    .I(SB_T3_WEST_SB_IN_B1),
    .O(WIRE_SB_T3_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T3_WEST_SB_IN_B16 (
    .I(SB_T3_WEST_SB_IN_B16),
    .O(WIRE_SB_T3_WEST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T4_EAST_SB_IN_B1 (
    .I(SB_T4_EAST_SB_IN_B1),
    .O(WIRE_SB_T4_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T4_EAST_SB_IN_B16 (
    .I(SB_T4_EAST_SB_IN_B16),
    .O(WIRE_SB_T4_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T4_NORTH_SB_IN_B1 (
    .I(SB_T4_NORTH_SB_IN_B1),
    .O(WIRE_SB_T4_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T4_NORTH_SB_IN_B16 (
    .I(SB_T4_NORTH_SB_IN_B16),
    .O(WIRE_SB_T4_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T4_SOUTH_SB_IN_B1 (
    .I(SB_T4_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T4_SOUTH_SB_IN_B16 (
    .I(SB_T4_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T4_WEST_SB_IN_B1 (
    .I(SB_T4_WEST_SB_IN_B1),
    .O(WIRE_SB_T4_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T4_WEST_SB_IN_B16 (
    .I(SB_T4_WEST_SB_IN_B16),
    .O(WIRE_SB_T4_WEST_SB_IN_B16_O)
);
corebit_and and_inst0 (
    .in0(coreir_eq_16_inst0_out),
    .in1(config_read[0]),
    .out(and_inst0_out)
);
corebit_and and_inst1 (
    .in0(coreir_eq_16_inst0_out),
    .in1(config_write[0]),
    .out(and_inst1_out)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
coreir_const #(
    .value(9'h1ff),
    .width(9)
) const_511_9 (
    .out(const_511_9_out)
);
wire [15:0] coreir_eq_16_inst0_in1;
assign coreir_eq_16_inst0_in1 = {config_config_addr[15],config_config_addr[14],config_config_addr[13],config_config_addr[12],config_config_addr[11],config_config_addr[10],config_config_addr[9],config_config_addr[8],config_config_addr[7],config_config_addr[6],config_config_addr[5],config_config_addr[4],config_config_addr[3],config_config_addr[2],config_config_addr[1],config_config_addr[0]};
coreir_eq #(
    .width(16)
) coreir_eq_16_inst0 (
    .in0(tile_id),
    .in1(coreir_eq_16_inst0_in1),
    .out(coreir_eq_16_inst0_out)
);
wire [7:0] read_data_mux_S;
assign read_data_mux_S = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
MuxWithDefaultWrapper_13_32_8_0 read_data_mux (
    .EN(and_inst0_out),
    .I_0(MemCore_inst0_read_config_data),
    .I_1(MemCore_inst0_read_config_data_1),
    .I_10(SB_ID0_5TRACKS_B1_MemCore_read_config_data),
    .I_11(SB_ID0_5TRACKS_B16_MemCore_read_config_data),
    .I_12(PowerDomainConfigReg_inst0_read_config_data),
    .I_2(MemCore_inst0_read_config_data_2),
    .I_3(CB_flush_read_config_data),
    .I_4(CB_input_width_16_num_0_read_config_data),
    .I_5(CB_input_width_16_num_1_read_config_data),
    .I_6(CB_input_width_16_num_2_read_config_data),
    .I_7(CB_input_width_16_num_3_read_config_data),
    .I_8(CB_input_width_1_num_0_read_config_data),
    .I_9(CB_input_width_1_num_1_read_config_data),
    .O(read_data_mux_O),
    .S(read_data_mux_S)
);
assign SB_T0_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1;
assign SB_T0_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T0_EAST_SB_OUT_B16;
assign SB_T0_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1;
assign SB_T0_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T0_NORTH_SB_OUT_B16;
assign SB_T0_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1;
assign SB_T0_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T0_SOUTH_SB_OUT_B16;
assign SB_T0_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1;
assign SB_T0_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T0_WEST_SB_OUT_B16;
assign SB_T1_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1;
assign SB_T1_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T1_EAST_SB_OUT_B16;
assign SB_T1_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1;
assign SB_T1_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T1_NORTH_SB_OUT_B16;
assign SB_T1_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1;
assign SB_T1_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T1_SOUTH_SB_OUT_B16;
assign SB_T1_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1;
assign SB_T1_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T1_WEST_SB_OUT_B16;
assign SB_T2_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1;
assign SB_T2_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T2_EAST_SB_OUT_B16;
assign SB_T2_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1;
assign SB_T2_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T2_NORTH_SB_OUT_B16;
assign SB_T2_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1;
assign SB_T2_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T2_SOUTH_SB_OUT_B16;
assign SB_T2_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1;
assign SB_T2_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T2_WEST_SB_OUT_B16;
assign SB_T3_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1;
assign SB_T3_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T3_EAST_SB_OUT_B16;
assign SB_T3_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1;
assign SB_T3_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T3_NORTH_SB_OUT_B16;
assign SB_T3_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1;
assign SB_T3_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T3_SOUTH_SB_OUT_B16;
assign SB_T3_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1;
assign SB_T3_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T3_WEST_SB_OUT_B16;
assign SB_T4_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1;
assign SB_T4_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T4_EAST_SB_OUT_B16;
assign SB_T4_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1;
assign SB_T4_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T4_NORTH_SB_OUT_B16;
assign SB_T4_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1;
assign SB_T4_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T4_SOUTH_SB_OUT_B16;
assign SB_T4_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1;
assign SB_T4_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T4_WEST_SB_OUT_B16;
assign clk_out = clk;
assign config_out_config_addr = config_config_addr;
assign config_out_config_data = config_config_data;
assign config_out_read = config_read;
assign config_out_write = config_write;
assign flush_out = flush;
assign hi = const_511_9_out;
assign lo = const_0_8_out;
assign read_config_data = PowerDomainOR_O;
assign reset_out = reset;
assign stall_out = stall;
endmodule

module CB_data_in_pond_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_data_in_pond (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [15:0] CB_data_in_pond_O;
wire [4:0] CB_data_in_pond_sel_inst0_O;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
MuxWrapperAOIImpl_20_16 CB_data_in_pond (
    .I_0(I_0),
    .I_1(I_1),
    .I_10(I_10),
    .I_11(I_11),
    .I_12(I_12),
    .I_13(I_13),
    .I_14(I_14),
    .I_15(I_15),
    .I_16(I_16),
    .I_17(I_17),
    .I_18(I_18),
    .I_19(I_19),
    .I_2(I_2),
    .I_3(I_3),
    .I_4(I_4),
    .I_5(I_5),
    .I_6(I_6),
    .I_7(I_7),
    .I_8(I_8),
    .I_9(I_9),
    .O(CB_data_in_pond_O),
    .S(CB_data_in_pond_sel_inst0_O)
);
CB_data_in_pond_sel CB_data_in_pond_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_data_in_pond_sel_inst0_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_data_in_pond_O;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module ADD (
    input [15:0] a,
    input [15:0] b,
    output [15:0] O0,
    output O1,
    output O2,
    output O3,
    output O4,
    output O5,
    input CLK,
    input ASYNCRESET
);
wire bit_const_0_None_out;
wire [15:0] const_0_16_out;
wire [16:0] const_0_17_out;
wire magma_Bit_and_inst0_out;
wire magma_Bit_and_inst1_out;
wire magma_Bit_and_inst2_out;
wire magma_Bit_and_inst3_out;
wire magma_Bit_not_inst0_out;
wire magma_Bit_not_inst1_out;
wire magma_Bit_not_inst2_out;
wire magma_Bit_or_inst0_out;
wire magma_UInt_16_eq_inst0_out;
wire [16:0] magma_UInt_17_add_inst0_out;
wire [16:0] magma_UInt_17_add_inst1_out;
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
coreir_const #(
    .value(17'h00000),
    .width(17)
) const_0_17 (
    .out(const_0_17_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(a[15]),
    .in1(b[15]),
    .out(magma_Bit_and_inst0_out)
);
corebit_and magma_Bit_and_inst1 (
    .in0(magma_Bit_and_inst0_out),
    .in1(magma_Bit_not_inst0_out),
    .out(magma_Bit_and_inst1_out)
);
corebit_and magma_Bit_and_inst2 (
    .in0(magma_Bit_not_inst1_out),
    .in1(magma_Bit_not_inst2_out),
    .out(magma_Bit_and_inst2_out)
);
corebit_and magma_Bit_and_inst3 (
    .in0(magma_Bit_and_inst2_out),
    .in1(magma_UInt_17_add_inst1_out[15]),
    .out(magma_Bit_and_inst3_out)
);
corebit_not magma_Bit_not_inst0 (
    .in(magma_UInt_17_add_inst1_out[15]),
    .out(magma_Bit_not_inst0_out)
);
corebit_not magma_Bit_not_inst1 (
    .in(a[15]),
    .out(magma_Bit_not_inst1_out)
);
corebit_not magma_Bit_not_inst2 (
    .in(b[15]),
    .out(magma_Bit_not_inst2_out)
);
corebit_or magma_Bit_or_inst0 (
    .in0(magma_Bit_and_inst1_out),
    .in1(magma_Bit_and_inst3_out),
    .out(magma_Bit_or_inst0_out)
);
wire [15:0] magma_UInt_16_eq_inst0_in0;
assign magma_UInt_16_eq_inst0_in0 = {magma_UInt_17_add_inst1_out[15],magma_UInt_17_add_inst1_out[14],magma_UInt_17_add_inst1_out[13],magma_UInt_17_add_inst1_out[12],magma_UInt_17_add_inst1_out[11],magma_UInt_17_add_inst1_out[10],magma_UInt_17_add_inst1_out[9],magma_UInt_17_add_inst1_out[8],magma_UInt_17_add_inst1_out[7],magma_UInt_17_add_inst1_out[6],magma_UInt_17_add_inst1_out[5],magma_UInt_17_add_inst1_out[4],magma_UInt_17_add_inst1_out[3],magma_UInt_17_add_inst1_out[2],magma_UInt_17_add_inst1_out[1],magma_UInt_17_add_inst1_out[0]};
coreir_eq #(
    .width(16)
) magma_UInt_16_eq_inst0 (
    .in0(magma_UInt_16_eq_inst0_in0),
    .in1(const_0_16_out),
    .out(magma_UInt_16_eq_inst0_out)
);
wire [16:0] magma_UInt_17_add_inst0_in0;
assign magma_UInt_17_add_inst0_in0 = {bit_const_0_None_out,a};
wire [16:0] magma_UInt_17_add_inst0_in1;
assign magma_UInt_17_add_inst0_in1 = {bit_const_0_None_out,b};
coreir_add #(
    .width(17)
) magma_UInt_17_add_inst0 (
    .in0(magma_UInt_17_add_inst0_in0),
    .in1(magma_UInt_17_add_inst0_in1),
    .out(magma_UInt_17_add_inst0_out)
);
coreir_add #(
    .width(17)
) magma_UInt_17_add_inst1 (
    .in0(magma_UInt_17_add_inst0_out),
    .in1(const_0_17_out),
    .out(magma_UInt_17_add_inst1_out)
);
assign O0 = {magma_UInt_17_add_inst1_out[15],magma_UInt_17_add_inst1_out[14],magma_UInt_17_add_inst1_out[13],magma_UInt_17_add_inst1_out[12],magma_UInt_17_add_inst1_out[11],magma_UInt_17_add_inst1_out[10],magma_UInt_17_add_inst1_out[9],magma_UInt_17_add_inst1_out[8],magma_UInt_17_add_inst1_out[7],magma_UInt_17_add_inst1_out[6],magma_UInt_17_add_inst1_out[5],magma_UInt_17_add_inst1_out[4],magma_UInt_17_add_inst1_out[3],magma_UInt_17_add_inst1_out[2],magma_UInt_17_add_inst1_out[1],magma_UInt_17_add_inst1_out[0]};
assign O1 = magma_UInt_17_add_inst1_out[16];
assign O2 = magma_UInt_16_eq_inst0_out;
assign O3 = magma_UInt_17_add_inst1_out[15];
assign O4 = magma_UInt_17_add_inst1_out[16];
assign O5 = magma_Bit_or_inst0_out;
endmodule

module ABSD (
    input [15:0] a,
    input [15:0] b,
    output [15:0] O0,
    output O1,
    output O2,
    output O3,
    output O4,
    output O5,
    input CLK,
    input ASYNCRESET
);
wire [15:0] Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire bit_const_0_None_out;
wire [15:0] const_0_16_out;
wire [16:0] const_1_17_out;
wire magma_Bits_16_eq_inst0_out;
wire [15:0] magma_Bits_16_not_inst0_out;
wire [15:0] magma_SInt_16_neg_inst0_out;
wire magma_SInt_16_sgt_inst0_out;
wire [16:0] magma_UInt_17_add_inst0_out;
wire [16:0] magma_UInt_17_add_inst1_out;
wire [15:0] Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_in0;
assign Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_in0 = {magma_UInt_17_add_inst1_out[15],magma_UInt_17_add_inst1_out[14],magma_UInt_17_add_inst1_out[13],magma_UInt_17_add_inst1_out[12],magma_UInt_17_add_inst1_out[11],magma_UInt_17_add_inst1_out[10],magma_UInt_17_add_inst1_out[9],magma_UInt_17_add_inst1_out[8],magma_UInt_17_add_inst1_out[7],magma_UInt_17_add_inst1_out[6],magma_UInt_17_add_inst1_out[5],magma_UInt_17_add_inst1_out[4],magma_UInt_17_add_inst1_out[3],magma_UInt_17_add_inst1_out[2],magma_UInt_17_add_inst1_out[1],magma_UInt_17_add_inst1_out[0]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_in0),
    .in1(magma_SInt_16_neg_inst0_out),
    .sel(magma_SInt_16_sgt_inst0_out),
    .out(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
coreir_const #(
    .value(17'h00001),
    .width(17)
) const_1_17 (
    .out(const_1_17_out)
);
coreir_eq #(
    .width(16)
) magma_Bits_16_eq_inst0 (
    .in0(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(const_0_16_out),
    .out(magma_Bits_16_eq_inst0_out)
);
coreir_not #(
    .width(16)
) magma_Bits_16_not_inst0 (
    .in(b),
    .out(magma_Bits_16_not_inst0_out)
);
wire [15:0] magma_SInt_16_neg_inst0_in;
assign magma_SInt_16_neg_inst0_in = {magma_UInt_17_add_inst1_out[15],magma_UInt_17_add_inst1_out[14],magma_UInt_17_add_inst1_out[13],magma_UInt_17_add_inst1_out[12],magma_UInt_17_add_inst1_out[11],magma_UInt_17_add_inst1_out[10],magma_UInt_17_add_inst1_out[9],magma_UInt_17_add_inst1_out[8],magma_UInt_17_add_inst1_out[7],magma_UInt_17_add_inst1_out[6],magma_UInt_17_add_inst1_out[5],magma_UInt_17_add_inst1_out[4],magma_UInt_17_add_inst1_out[3],magma_UInt_17_add_inst1_out[2],magma_UInt_17_add_inst1_out[1],magma_UInt_17_add_inst1_out[0]};
coreir_neg #(
    .width(16)
) magma_SInt_16_neg_inst0 (
    .in(magma_SInt_16_neg_inst0_in),
    .out(magma_SInt_16_neg_inst0_out)
);
wire [15:0] magma_SInt_16_sgt_inst0_in1;
assign magma_SInt_16_sgt_inst0_in1 = {magma_UInt_17_add_inst1_out[15],magma_UInt_17_add_inst1_out[14],magma_UInt_17_add_inst1_out[13],magma_UInt_17_add_inst1_out[12],magma_UInt_17_add_inst1_out[11],magma_UInt_17_add_inst1_out[10],magma_UInt_17_add_inst1_out[9],magma_UInt_17_add_inst1_out[8],magma_UInt_17_add_inst1_out[7],magma_UInt_17_add_inst1_out[6],magma_UInt_17_add_inst1_out[5],magma_UInt_17_add_inst1_out[4],magma_UInt_17_add_inst1_out[3],magma_UInt_17_add_inst1_out[2],magma_UInt_17_add_inst1_out[1],magma_UInt_17_add_inst1_out[0]};
coreir_sgt #(
    .width(16)
) magma_SInt_16_sgt_inst0 (
    .in0(const_0_16_out),
    .in1(magma_SInt_16_sgt_inst0_in1),
    .out(magma_SInt_16_sgt_inst0_out)
);
wire [16:0] magma_UInt_17_add_inst0_in0;
assign magma_UInt_17_add_inst0_in0 = {bit_const_0_None_out,a};
wire [16:0] magma_UInt_17_add_inst0_in1;
assign magma_UInt_17_add_inst0_in1 = {bit_const_0_None_out,magma_Bits_16_not_inst0_out};
coreir_add #(
    .width(17)
) magma_UInt_17_add_inst0 (
    .in0(magma_UInt_17_add_inst0_in0),
    .in1(magma_UInt_17_add_inst0_in1),
    .out(magma_UInt_17_add_inst0_out)
);
coreir_add #(
    .width(17)
) magma_UInt_17_add_inst1 (
    .in0(magma_UInt_17_add_inst0_out),
    .in1(const_1_17_out),
    .out(magma_UInt_17_add_inst1_out)
);
assign O0 = Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign O1 = bit_const_0_None_out;
assign O2 = magma_Bits_16_eq_inst0_out;
assign O3 = Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15];
assign O4 = bit_const_0_None_out;
assign O5 = bit_const_0_None_out;
endmodule

module PE_gen (
    input [80:0] inst,
    input [66:0] inputs,
    input clk_en,
    output [16:0] O,
    input CLK,
    input ASYNCRESET
);
wire [15:0] ABSD_inst0_O0;
wire ABSD_inst0_O1;
wire ABSD_inst0_O2;
wire ABSD_inst0_O3;
wire ABSD_inst0_O4;
wire ABSD_inst0_O5;
wire [15:0] ADD_inst0_O0;
wire ADD_inst0_O1;
wire ADD_inst0_O2;
wire ADD_inst0_O3;
wire ADD_inst0_O4;
wire ADD_inst0_O5;
wire [15:0] ADD_inst1_O0;
wire ADD_inst1_O1;
wire ADD_inst1_O2;
wire ADD_inst1_O3;
wire ADD_inst1_O4;
wire ADD_inst1_O5;
wire [15:0] ADD_inst2_O0;
wire ADD_inst2_O1;
wire ADD_inst2_O2;
wire ADD_inst2_O3;
wire ADD_inst2_O4;
wire ADD_inst2_O5;
wire Cond_inst0_O;
wire Cond_inst1_O;
wire Cond_inst2_O;
wire [15:0] GTE_inst0_O0;
wire GTE_inst0_O1;
wire GTE_inst0_O2;
wire GTE_inst0_O3;
wire GTE_inst0_O4;
wire GTE_inst0_O5;
wire [15:0] LTE_inst0_O0;
wire LTE_inst0_O1;
wire LTE_inst0_O2;
wire LTE_inst0_O3;
wire LTE_inst0_O4;
wire LTE_inst0_O5;
wire LUT_inst0_O;
wire [15:0] MUL_inst0_O;
wire [0:0] Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out;
wire [15:0] Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst10$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst11$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst13$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst14$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst15$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst16$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst17$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst18$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst19$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst20$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst21$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst22$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst23$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst24$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst25$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst26$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst27$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst28$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst29$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst30$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst31$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst32$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst6$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst8$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst9$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux_inst0$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] SHR_inst0_O0;
wire SHR_inst0_O1;
wire SHR_inst0_O2;
wire SHR_inst0_O3;
wire SHR_inst0_O4;
wire SHR_inst0_O5;
wire [15:0] SUB_inst0_O0;
wire SUB_inst0_O1;
wire SUB_inst0_O2;
wire SUB_inst0_O3;
wire SUB_inst0_O4;
wire SUB_inst0_O5;
wire [0:0] const_0_1_out;
wire [1:0] const_0_2_out;
wire [2:0] const_0_3_out;
wire [3:0] const_0_4_out;
wire [0:0] const_1_1_out;
wire [1:0] const_1_2_out;
wire [2:0] const_1_3_out;
wire [3:0] const_1_4_out;
wire [1:0] const_2_2_out;
wire [2:0] const_2_3_out;
wire [3:0] const_2_4_out;
wire [1:0] const_3_2_out;
wire [2:0] const_3_3_out;
wire [3:0] const_3_4_out;
wire [2:0] const_4_3_out;
wire [3:0] const_4_4_out;
wire [3:0] const_5_4_out;
wire [3:0] const_6_4_out;
wire [3:0] const_7_4_out;
wire [3:0] const_8_4_out;
wire magma_Bits_1_eq_inst0_out;
wire magma_Bits_1_eq_inst1_out;
wire magma_Bits_1_eq_inst10_out;
wire magma_Bits_1_eq_inst11_out;
wire magma_Bits_1_eq_inst12_out;
wire magma_Bits_1_eq_inst13_out;
wire magma_Bits_1_eq_inst14_out;
wire magma_Bits_1_eq_inst15_out;
wire magma_Bits_1_eq_inst16_out;
wire magma_Bits_1_eq_inst17_out;
wire magma_Bits_1_eq_inst18_out;
wire magma_Bits_1_eq_inst19_out;
wire magma_Bits_1_eq_inst2_out;
wire magma_Bits_1_eq_inst3_out;
wire magma_Bits_1_eq_inst4_out;
wire magma_Bits_1_eq_inst5_out;
wire magma_Bits_1_eq_inst6_out;
wire magma_Bits_1_eq_inst7_out;
wire magma_Bits_1_eq_inst8_out;
wire magma_Bits_1_eq_inst9_out;
wire magma_Bits_2_eq_inst0_out;
wire magma_Bits_2_eq_inst1_out;
wire magma_Bits_2_eq_inst2_out;
wire magma_Bits_2_eq_inst3_out;
wire magma_Bits_3_eq_inst0_out;
wire magma_Bits_3_eq_inst1_out;
wire magma_Bits_3_eq_inst2_out;
wire magma_Bits_3_eq_inst3_out;
wire magma_Bits_3_eq_inst4_out;
wire magma_Bits_4_eq_inst0_out;
wire magma_Bits_4_eq_inst1_out;
wire magma_Bits_4_eq_inst2_out;
wire magma_Bits_4_eq_inst3_out;
wire magma_Bits_4_eq_inst4_out;
wire magma_Bits_4_eq_inst5_out;
wire magma_Bits_4_eq_inst6_out;
wire magma_Bits_4_eq_inst7_out;
wire magma_Bits_4_eq_inst8_out;
wire [15:0] ABSD_inst0_a;
assign ABSD_inst0_a = {inputs[15],inputs[14],inputs[13],inputs[12],inputs[11],inputs[10],inputs[9],inputs[8],inputs[7],inputs[6],inputs[5],inputs[4],inputs[3],inputs[2],inputs[1],inputs[0]};
ABSD ABSD_inst0 (
    .a(ABSD_inst0_a),
    .b(Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join_out),
    .O0(ABSD_inst0_O0),
    .O1(ABSD_inst0_O1),
    .O2(ABSD_inst0_O2),
    .O3(ABSD_inst0_O3),
    .O4(ABSD_inst0_O4),
    .O5(ABSD_inst0_O5),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
wire [15:0] ADD_inst0_a;
assign ADD_inst0_a = {inputs[15],inputs[14],inputs[13],inputs[12],inputs[11],inputs[10],inputs[9],inputs[8],inputs[7],inputs[6],inputs[5],inputs[4],inputs[3],inputs[2],inputs[1],inputs[0]};
wire [15:0] ADD_inst0_b;
assign ADD_inst0_b = {inputs[47],inputs[46],inputs[45],inputs[44],inputs[43],inputs[42],inputs[41],inputs[40],inputs[39],inputs[38],inputs[37],inputs[36],inputs[35],inputs[34],inputs[33],inputs[32]};
ADD ADD_inst0 (
    .a(ADD_inst0_a),
    .b(ADD_inst0_b),
    .O0(ADD_inst0_O0),
    .O1(ADD_inst0_O1),
    .O2(ADD_inst0_O2),
    .O3(ADD_inst0_O3),
    .O4(ADD_inst0_O4),
    .O5(ADD_inst0_O5),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
wire [15:0] ADD_inst1_a;
assign ADD_inst1_a = {inputs[63],inputs[62],inputs[61],inputs[60],inputs[59],inputs[58],inputs[57],inputs[56],inputs[55],inputs[54],inputs[53],inputs[52],inputs[51],inputs[50],inputs[49],inputs[48]};
ADD ADD_inst1 (
    .a(ADD_inst1_a),
    .b(Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out),
    .O0(ADD_inst1_O0),
    .O1(ADD_inst1_O1),
    .O2(ADD_inst1_O2),
    .O3(ADD_inst1_O3),
    .O4(ADD_inst1_O4),
    .O5(ADD_inst1_O5),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
wire [15:0] ADD_inst2_b;
assign ADD_inst2_b = {inputs[31],inputs[30],inputs[29],inputs[28],inputs[27],inputs[26],inputs[25],inputs[24],inputs[23],inputs[22],inputs[21],inputs[20],inputs[19],inputs[18],inputs[17],inputs[16]};
ADD ADD_inst2 (
    .a(Mux2xBits16_inst23$coreir_commonlib_mux2x16_inst0$_join_out),
    .b(ADD_inst2_b),
    .O0(ADD_inst2_O0),
    .O1(ADD_inst2_O1),
    .O2(ADD_inst2_O2),
    .O3(ADD_inst2_O3),
    .O4(ADD_inst2_O4),
    .O5(ADD_inst2_O5),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
wire [4:0] Cond_inst0_code;
assign Cond_inst0_code = {inst[4],inst[3],inst[2],inst[1],inst[0]};
Cond Cond_inst0 (
    .code(Cond_inst0_code),
    .alu(LTE_inst0_O1),
    .Z(LTE_inst0_O2),
    .N(LTE_inst0_O3),
    .C(LTE_inst0_O4),
    .V(LTE_inst0_O5),
    .O(Cond_inst0_O),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
wire [4:0] Cond_inst1_code;
assign Cond_inst1_code = {inst[9],inst[8],inst[7],inst[6],inst[5]};
Cond Cond_inst1 (
    .code(Cond_inst1_code),
    .alu(GTE_inst0_O1),
    .Z(GTE_inst0_O2),
    .N(GTE_inst0_O3),
    .C(GTE_inst0_O4),
    .V(GTE_inst0_O5),
    .O(Cond_inst1_O),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
wire [4:0] Cond_inst2_code;
assign Cond_inst2_code = {inst[14],inst[13],inst[12],inst[11],inst[10]};
Cond Cond_inst2 (
    .code(Cond_inst2_code),
    .alu(SUB_inst0_O1),
    .Z(SUB_inst0_O2),
    .N(SUB_inst0_O3),
    .C(SUB_inst0_O4),
    .V(SUB_inst0_O5),
    .O(Cond_inst2_O),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
GTE GTE_inst0 (
    .signed_(inst[70]),
    .a(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
    .b(Mux2xBits16_inst9$coreir_commonlib_mux2x16_inst0$_join_out),
    .O0(GTE_inst0_O0),
    .O1(GTE_inst0_O1),
    .O2(GTE_inst0_O2),
    .O3(GTE_inst0_O3),
    .O4(GTE_inst0_O4),
    .O5(GTE_inst0_O5),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
wire [15:0] LTE_inst0_a;
assign LTE_inst0_a = {inputs[15],inputs[14],inputs[13],inputs[12],inputs[11],inputs[10],inputs[9],inputs[8],inputs[7],inputs[6],inputs[5],inputs[4],inputs[3],inputs[2],inputs[1],inputs[0]};
LTE LTE_inst0 (
    .signed_(inst[69]),
    .a(LTE_inst0_a),
    .b(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out),
    .O0(LTE_inst0_O0),
    .O1(LTE_inst0_O1),
    .O2(LTE_inst0_O2),
    .O3(LTE_inst0_O3),
    .O4(LTE_inst0_O4),
    .O5(LTE_inst0_O5),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
wire [7:0] LUT_inst0_lut;
assign LUT_inst0_lut = {inst[80],inst[79],inst[78],inst[77],inst[76],inst[75],inst[74],inst[73]};
LUT LUT_inst0 (
    .lut(LUT_inst0_lut),
    .bit0(inputs[64]),
    .bit1(inputs[65]),
    .bit2(inputs[66]),
    .O(LUT_inst0_O),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
MUL MUL_inst0 (
    .instr(inst[16:15]),
    .signed_(inst[72]),
    .a(Mux2xBits16_inst17$coreir_commonlib_mux2x16_inst0$_join_out),
    .b(Mux2xBits16_inst19$coreir_commonlib_mux2x16_inst0$_join_out),
    .O(MUL_inst0_O),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Cond_inst2_O),
    .in1(Cond_inst2_O),
    .sel(magma_Bits_3_eq_inst0_out),
    .out(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(Cond_inst1_O),
    .sel(magma_Bits_3_eq_inst1_out),
    .out(Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(inst[49]),
    .sel(magma_Bits_3_eq_inst2_out),
    .out(Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(Cond_inst0_O),
    .sel(magma_Bits_3_eq_inst3_out),
    .out(Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(LUT_inst0_O),
    .sel(magma_Bits_3_eq_inst4_out),
    .out(Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(ADD_inst0_O0),
    .in1(ADD_inst0_O0),
    .sel(magma_Bits_1_eq_inst0_out),
    .out(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_in1 = {inputs[47],inputs[46],inputs[45],inputs[44],inputs[43],inputs[42],inputs[41],inputs[40],inputs[39],inputs[38],inputs[37],inputs[36],inputs[35],inputs[34],inputs[33],inputs[32]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_1_eq_inst1_out),
    .out(Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst10$coreir_commonlib_mux2x16_inst0$_join_in0;
assign Mux2xBits16_inst10$coreir_commonlib_mux2x16_inst0$_join_in0 = {inputs[31],inputs[30],inputs[29],inputs[28],inputs[27],inputs[26],inputs[25],inputs[24],inputs[23],inputs[22],inputs[21],inputs[20],inputs[19],inputs[18],inputs[17],inputs[16]};
wire [15:0] Mux2xBits16_inst10$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst10$coreir_commonlib_mux2x16_inst0$_join_in1 = {inputs[31],inputs[30],inputs[29],inputs[28],inputs[27],inputs[26],inputs[25],inputs[24],inputs[23],inputs[22],inputs[21],inputs[20],inputs[19],inputs[18],inputs[17],inputs[16]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst10$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst10$coreir_commonlib_mux2x16_inst0$_join_in0),
    .in1(Mux2xBits16_inst10$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_1_eq_inst10_out),
    .out(Mux2xBits16_inst10$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst11$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst11$coreir_commonlib_mux2x16_inst0$_join_in1 = {inst[48],inst[47],inst[46],inst[45],inst[44],inst[43],inst[42],inst[41],inst[40],inst[39],inst[38],inst[37],inst[36],inst[35],inst[34],inst[33]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst11$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst10$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(Mux2xBits16_inst11$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_1_eq_inst11_out),
    .out(Mux2xBits16_inst11$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join_in0;
assign Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join_in0 = {inst[32],inst[31],inst[30],inst[29],inst[28],inst[27],inst[26],inst[25],inst[24],inst[23],inst[22],inst[21],inst[20],inst[19],inst[18],inst[17]};
wire [15:0] Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join_in1 = {inst[32],inst[31],inst[30],inst[29],inst[28],inst[27],inst[26],inst[25],inst[24],inst[23],inst[22],inst[21],inst[20],inst[19],inst[18],inst[17]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join_in0),
    .in1(Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_1_eq_inst12_out),
    .out(Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst13$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst13$coreir_commonlib_mux2x16_inst0$_join_in1 = {inputs[31],inputs[30],inputs[29],inputs[28],inputs[27],inputs[26],inputs[25],inputs[24],inputs[23],inputs[22],inputs[21],inputs[20],inputs[19],inputs[18],inputs[17],inputs[16]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst13$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(Mux2xBits16_inst13$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_1_eq_inst13_out),
    .out(Mux2xBits16_inst13$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst14$coreir_commonlib_mux2x16_inst0$_join_in0;
assign Mux2xBits16_inst14$coreir_commonlib_mux2x16_inst0$_join_in0 = {inst[32],inst[31],inst[30],inst[29],inst[28],inst[27],inst[26],inst[25],inst[24],inst[23],inst[22],inst[21],inst[20],inst[19],inst[18],inst[17]};
wire [15:0] Mux2xBits16_inst14$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst14$coreir_commonlib_mux2x16_inst0$_join_in1 = {inst[32],inst[31],inst[30],inst[29],inst[28],inst[27],inst[26],inst[25],inst[24],inst[23],inst[22],inst[21],inst[20],inst[19],inst[18],inst[17]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst14$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst14$coreir_commonlib_mux2x16_inst0$_join_in0),
    .in1(Mux2xBits16_inst14$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_1_eq_inst14_out),
    .out(Mux2xBits16_inst14$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst15$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst15$coreir_commonlib_mux2x16_inst0$_join_in1 = {inputs[31],inputs[30],inputs[29],inputs[28],inputs[27],inputs[26],inputs[25],inputs[24],inputs[23],inputs[22],inputs[21],inputs[20],inputs[19],inputs[18],inputs[17],inputs[16]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst15$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst14$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(Mux2xBits16_inst15$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_1_eq_inst15_out),
    .out(Mux2xBits16_inst15$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst16$coreir_commonlib_mux2x16_inst0$_join_in0;
assign Mux2xBits16_inst16$coreir_commonlib_mux2x16_inst0$_join_in0 = {inputs[15],inputs[14],inputs[13],inputs[12],inputs[11],inputs[10],inputs[9],inputs[8],inputs[7],inputs[6],inputs[5],inputs[4],inputs[3],inputs[2],inputs[1],inputs[0]};
wire [15:0] Mux2xBits16_inst16$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst16$coreir_commonlib_mux2x16_inst0$_join_in1 = {inputs[15],inputs[14],inputs[13],inputs[12],inputs[11],inputs[10],inputs[9],inputs[8],inputs[7],inputs[6],inputs[5],inputs[4],inputs[3],inputs[2],inputs[1],inputs[0]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst16$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst16$coreir_commonlib_mux2x16_inst0$_join_in0),
    .in1(Mux2xBits16_inst16$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_1_eq_inst16_out),
    .out(Mux2xBits16_inst16$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst17$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst16$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(LTE_inst0_O0),
    .sel(magma_Bits_1_eq_inst17_out),
    .out(Mux2xBits16_inst17$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst18$coreir_commonlib_mux2x16_inst0$_join_in0;
assign Mux2xBits16_inst18$coreir_commonlib_mux2x16_inst0$_join_in0 = {inst[32],inst[31],inst[30],inst[29],inst[28],inst[27],inst[26],inst[25],inst[24],inst[23],inst[22],inst[21],inst[20],inst[19],inst[18],inst[17]};
wire [15:0] Mux2xBits16_inst18$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst18$coreir_commonlib_mux2x16_inst0$_join_in1 = {inst[32],inst[31],inst[30],inst[29],inst[28],inst[27],inst[26],inst[25],inst[24],inst[23],inst[22],inst[21],inst[20],inst[19],inst[18],inst[17]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst18$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst18$coreir_commonlib_mux2x16_inst0$_join_in0),
    .in1(Mux2xBits16_inst18$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_1_eq_inst18_out),
    .out(Mux2xBits16_inst18$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst19$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst19$coreir_commonlib_mux2x16_inst0$_join_in1 = {inputs[63],inputs[62],inputs[61],inputs[60],inputs[59],inputs[58],inputs[57],inputs[56],inputs[55],inputs[54],inputs[53],inputs[52],inputs[51],inputs[50],inputs[49],inputs[48]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst19$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst18$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(Mux2xBits16_inst19$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_1_eq_inst19_out),
    .out(Mux2xBits16_inst19$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_in0;
assign Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_in0 = {inputs[31],inputs[30],inputs[29],inputs[28],inputs[27],inputs[26],inputs[25],inputs[24],inputs[23],inputs[22],inputs[21],inputs[20],inputs[19],inputs[18],inputs[17],inputs[16]};
wire [15:0] Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_in1 = {inputs[31],inputs[30],inputs[29],inputs[28],inputs[27],inputs[26],inputs[25],inputs[24],inputs[23],inputs[22],inputs[21],inputs[20],inputs[19],inputs[18],inputs[17],inputs[16]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_in0),
    .in1(Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_1_eq_inst2_out),
    .out(Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst20$coreir_commonlib_mux2x16_inst0$_join_in0;
assign Mux2xBits16_inst20$coreir_commonlib_mux2x16_inst0$_join_in0 = {inst[32],inst[31],inst[30],inst[29],inst[28],inst[27],inst[26],inst[25],inst[24],inst[23],inst[22],inst[21],inst[20],inst[19],inst[18],inst[17]};
wire [15:0] Mux2xBits16_inst20$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst20$coreir_commonlib_mux2x16_inst0$_join_in1 = {inst[32],inst[31],inst[30],inst[29],inst[28],inst[27],inst[26],inst[25],inst[24],inst[23],inst[22],inst[21],inst[20],inst[19],inst[18],inst[17]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst20$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst20$coreir_commonlib_mux2x16_inst0$_join_in0),
    .in1(Mux2xBits16_inst20$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_2_eq_inst0_out),
    .out(Mux2xBits16_inst20$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst21$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst20$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(MUL_inst0_O),
    .sel(magma_Bits_2_eq_inst1_out),
    .out(Mux2xBits16_inst21$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst22$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst21$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(ADD_inst1_O0),
    .sel(magma_Bits_2_eq_inst2_out),
    .out(Mux2xBits16_inst22$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst23$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst23$coreir_commonlib_mux2x16_inst0$_join_in1 = {inputs[63],inputs[62],inputs[61],inputs[60],inputs[59],inputs[58],inputs[57],inputs[56],inputs[55],inputs[54],inputs[53],inputs[52],inputs[51],inputs[50],inputs[49],inputs[48]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst23$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst22$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(Mux2xBits16_inst23$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_2_eq_inst3_out),
    .out(Mux2xBits16_inst23$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst24$coreir_commonlib_mux2x16_inst0$_join (
    .in0(SUB_inst0_O0),
    .in1(SUB_inst0_O0),
    .sel(magma_Bits_4_eq_inst0_out),
    .out(Mux2xBits16_inst24$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst25$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst24$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(GTE_inst0_O0),
    .sel(magma_Bits_4_eq_inst1_out),
    .out(Mux2xBits16_inst25$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst26$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst25$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(MUL_inst0_O),
    .sel(magma_Bits_4_eq_inst2_out),
    .out(Mux2xBits16_inst26$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst27$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst27$coreir_commonlib_mux2x16_inst0$_join_in1 = {inst[48],inst[47],inst[46],inst[45],inst[44],inst[43],inst[42],inst[41],inst[40],inst[39],inst[38],inst[37],inst[36],inst[35],inst[34],inst[33]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst27$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst26$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(Mux2xBits16_inst27$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_4_eq_inst3_out),
    .out(Mux2xBits16_inst27$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst28$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst27$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(Mux_inst0$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
    .sel(magma_Bits_4_eq_inst4_out),
    .out(Mux2xBits16_inst28$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst29$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst28$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(LTE_inst0_O0),
    .sel(magma_Bits_4_eq_inst5_out),
    .out(Mux2xBits16_inst29$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_in1 = {inst[48],inst[47],inst[46],inst[45],inst[44],inst[43],inst[42],inst[41],inst[40],inst[39],inst[38],inst[37],inst[36],inst[35],inst[34],inst[33]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_1_eq_inst3_out),
    .out(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst30$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst29$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(ABSD_inst0_O0),
    .sel(magma_Bits_4_eq_inst6_out),
    .out(Mux2xBits16_inst30$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst31$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst30$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(ADD_inst2_O0),
    .sel(magma_Bits_4_eq_inst7_out),
    .out(Mux2xBits16_inst31$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst32$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst31$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(SHR_inst0_O0),
    .sel(magma_Bits_4_eq_inst8_out),
    .out(Mux2xBits16_inst32$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_in0;
assign Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_in0 = {inst[32],inst[31],inst[30],inst[29],inst[28],inst[27],inst[26],inst[25],inst[24],inst[23],inst[22],inst[21],inst[20],inst[19],inst[18],inst[17]};
wire [15:0] Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_in1 = {inst[32],inst[31],inst[30],inst[29],inst[28],inst[27],inst[26],inst[25],inst[24],inst[23],inst[22],inst[21],inst[20],inst[19],inst[18],inst[17]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_in0),
    .in1(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_1_eq_inst4_out),
    .out(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join_in1 = {inputs[31],inputs[30],inputs[29],inputs[28],inputs[27],inputs[26],inputs[25],inputs[24],inputs[23],inputs[22],inputs[21],inputs[20],inputs[19],inputs[18],inputs[17],inputs[16]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_1_eq_inst5_out),
    .out(Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst6$coreir_commonlib_mux2x16_inst0$_join_in0;
assign Mux2xBits16_inst6$coreir_commonlib_mux2x16_inst0$_join_in0 = {inputs[15],inputs[14],inputs[13],inputs[12],inputs[11],inputs[10],inputs[9],inputs[8],inputs[7],inputs[6],inputs[5],inputs[4],inputs[3],inputs[2],inputs[1],inputs[0]};
wire [15:0] Mux2xBits16_inst6$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst6$coreir_commonlib_mux2x16_inst0$_join_in1 = {inputs[15],inputs[14],inputs[13],inputs[12],inputs[11],inputs[10],inputs[9],inputs[8],inputs[7],inputs[6],inputs[5],inputs[4],inputs[3],inputs[2],inputs[1],inputs[0]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst6$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst6$coreir_commonlib_mux2x16_inst0$_join_in0),
    .in1(Mux2xBits16_inst6$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_1_eq_inst6_out),
    .out(Mux2xBits16_inst6$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_in1 = {inst[48],inst[47],inst[46],inst[45],inst[44],inst[43],inst[42],inst[41],inst[40],inst[39],inst[38],inst[37],inst[36],inst[35],inst[34],inst[33]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst6$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_1_eq_inst7_out),
    .out(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst8$coreir_commonlib_mux2x16_inst0$_join_in0;
assign Mux2xBits16_inst8$coreir_commonlib_mux2x16_inst0$_join_in0 = {inst[32],inst[31],inst[30],inst[29],inst[28],inst[27],inst[26],inst[25],inst[24],inst[23],inst[22],inst[21],inst[20],inst[19],inst[18],inst[17]};
wire [15:0] Mux2xBits16_inst8$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst8$coreir_commonlib_mux2x16_inst0$_join_in1 = {inst[32],inst[31],inst[30],inst[29],inst[28],inst[27],inst[26],inst[25],inst[24],inst[23],inst[22],inst[21],inst[20],inst[19],inst[18],inst[17]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst8$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst8$coreir_commonlib_mux2x16_inst0$_join_in0),
    .in1(Mux2xBits16_inst8$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_1_eq_inst8_out),
    .out(Mux2xBits16_inst8$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux2xBits16_inst9$coreir_commonlib_mux2x16_inst0$_join_in1;
assign Mux2xBits16_inst9$coreir_commonlib_mux2x16_inst0$_join_in1 = {inputs[31],inputs[30],inputs[29],inputs[28],inputs[27],inputs[26],inputs[25],inputs[24],inputs[23],inputs[22],inputs[21],inputs[20],inputs[19],inputs[18],inputs[17],inputs[16]};
coreir_mux #(
    .width(16)
) Mux2xBits16_inst9$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst8$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(Mux2xBits16_inst9$coreir_commonlib_mux2x16_inst0$_join_in1),
    .sel(magma_Bits_1_eq_inst9_out),
    .out(Mux2xBits16_inst9$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] Mux_inst0$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_in0;
assign Mux_inst0$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_in0 = {inputs[15],inputs[14],inputs[13],inputs[12],inputs[11],inputs[10],inputs[9],inputs[8],inputs[7],inputs[6],inputs[5],inputs[4],inputs[3],inputs[2],inputs[1],inputs[0]};
coreir_mux #(
    .width(16)
) Mux_inst0$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux_inst0$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_in0),
    .in1(Mux2xBits16_inst15$coreir_commonlib_mux2x16_inst0$_join_out),
    .sel(inputs[64]),
    .out(Mux_inst0$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
wire [15:0] SHR_inst0_a;
assign SHR_inst0_a = {inputs[15],inputs[14],inputs[13],inputs[12],inputs[11],inputs[10],inputs[9],inputs[8],inputs[7],inputs[6],inputs[5],inputs[4],inputs[3],inputs[2],inputs[1],inputs[0]};
SHR SHR_inst0 (
    .signed_(inst[71]),
    .a(SHR_inst0_a),
    .b(Mux2xBits16_inst13$coreir_commonlib_mux2x16_inst0$_join_out),
    .O0(SHR_inst0_O0),
    .O1(SHR_inst0_O1),
    .O2(SHR_inst0_O2),
    .O3(SHR_inst0_O3),
    .O4(SHR_inst0_O4),
    .O5(SHR_inst0_O5),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
wire [15:0] SUB_inst0_a;
assign SUB_inst0_a = {inputs[15],inputs[14],inputs[13],inputs[12],inputs[11],inputs[10],inputs[9],inputs[8],inputs[7],inputs[6],inputs[5],inputs[4],inputs[3],inputs[2],inputs[1],inputs[0]};
SUB SUB_inst0 (
    .a(SUB_inst0_a),
    .b(Mux2xBits16_inst11$coreir_commonlib_mux2x16_inst0$_join_out),
    .O0(SUB_inst0_O0),
    .O1(SUB_inst0_O1),
    .O2(SUB_inst0_O2),
    .O3(SUB_inst0_O3),
    .O4(SUB_inst0_O4),
    .O5(SUB_inst0_O5),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
coreir_const #(
    .value(1'h0),
    .width(1)
) const_0_1 (
    .out(const_0_1_out)
);
coreir_const #(
    .value(2'h0),
    .width(2)
) const_0_2 (
    .out(const_0_2_out)
);
coreir_const #(
    .value(3'h0),
    .width(3)
) const_0_3 (
    .out(const_0_3_out)
);
coreir_const #(
    .value(4'h0),
    .width(4)
) const_0_4 (
    .out(const_0_4_out)
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_const #(
    .value(2'h1),
    .width(2)
) const_1_2 (
    .out(const_1_2_out)
);
coreir_const #(
    .value(3'h1),
    .width(3)
) const_1_3 (
    .out(const_1_3_out)
);
coreir_const #(
    .value(4'h1),
    .width(4)
) const_1_4 (
    .out(const_1_4_out)
);
coreir_const #(
    .value(2'h2),
    .width(2)
) const_2_2 (
    .out(const_2_2_out)
);
coreir_const #(
    .value(3'h2),
    .width(3)
) const_2_3 (
    .out(const_2_3_out)
);
coreir_const #(
    .value(4'h2),
    .width(4)
) const_2_4 (
    .out(const_2_4_out)
);
coreir_const #(
    .value(2'h3),
    .width(2)
) const_3_2 (
    .out(const_3_2_out)
);
coreir_const #(
    .value(3'h3),
    .width(3)
) const_3_3 (
    .out(const_3_3_out)
);
coreir_const #(
    .value(4'h3),
    .width(4)
) const_3_4 (
    .out(const_3_4_out)
);
coreir_const #(
    .value(3'h4),
    .width(3)
) const_4_3 (
    .out(const_4_3_out)
);
coreir_const #(
    .value(4'h4),
    .width(4)
) const_4_4 (
    .out(const_4_4_out)
);
coreir_const #(
    .value(4'h5),
    .width(4)
) const_5_4 (
    .out(const_5_4_out)
);
coreir_const #(
    .value(4'h6),
    .width(4)
) const_6_4 (
    .out(const_6_4_out)
);
coreir_const #(
    .value(4'h7),
    .width(4)
) const_7_4 (
    .out(const_7_4_out)
);
coreir_const #(
    .value(4'h8),
    .width(4)
) const_8_4 (
    .out(const_8_4_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst0 (
    .in0(const_0_1_out),
    .in1(inst[54]),
    .out(magma_Bits_1_eq_inst0_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst1 (
    .in0(const_1_1_out),
    .in1(inst[54]),
    .out(magma_Bits_1_eq_inst1_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst10 (
    .in0(const_0_1_out),
    .in1(inst[58]),
    .out(magma_Bits_1_eq_inst10_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst11 (
    .in0(const_1_1_out),
    .in1(inst[58]),
    .out(magma_Bits_1_eq_inst11_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst12 (
    .in0(const_0_1_out),
    .in1(inst[59]),
    .out(magma_Bits_1_eq_inst12_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst13 (
    .in0(const_1_1_out),
    .in1(inst[59]),
    .out(magma_Bits_1_eq_inst13_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst14 (
    .in0(const_0_1_out),
    .in1(inst[60]),
    .out(magma_Bits_1_eq_inst14_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst15 (
    .in0(const_1_1_out),
    .in1(inst[60]),
    .out(magma_Bits_1_eq_inst15_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst16 (
    .in0(const_0_1_out),
    .in1(inst[51]),
    .out(magma_Bits_1_eq_inst16_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst17 (
    .in0(const_1_1_out),
    .in1(inst[51]),
    .out(magma_Bits_1_eq_inst17_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst18 (
    .in0(const_0_1_out),
    .in1(inst[61]),
    .out(magma_Bits_1_eq_inst18_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst19 (
    .in0(const_1_1_out),
    .in1(inst[61]),
    .out(magma_Bits_1_eq_inst19_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst2 (
    .in0(const_0_1_out),
    .in1(inst[55]),
    .out(magma_Bits_1_eq_inst2_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst3 (
    .in0(const_1_1_out),
    .in1(inst[55]),
    .out(magma_Bits_1_eq_inst3_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst4 (
    .in0(const_0_1_out),
    .in1(inst[56]),
    .out(magma_Bits_1_eq_inst4_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst5 (
    .in0(const_1_1_out),
    .in1(inst[56]),
    .out(magma_Bits_1_eq_inst5_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst6 (
    .in0(const_0_1_out),
    .in1(inst[50]),
    .out(magma_Bits_1_eq_inst6_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst7 (
    .in0(const_1_1_out),
    .in1(inst[50]),
    .out(magma_Bits_1_eq_inst7_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst8 (
    .in0(const_0_1_out),
    .in1(inst[57]),
    .out(magma_Bits_1_eq_inst8_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst9 (
    .in0(const_1_1_out),
    .in1(inst[57]),
    .out(magma_Bits_1_eq_inst9_out)
);
wire [1:0] magma_Bits_2_eq_inst0_in1;
assign magma_Bits_2_eq_inst0_in1 = {inst[53],inst[52]};
coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst0 (
    .in0(const_0_2_out),
    .in1(magma_Bits_2_eq_inst0_in1),
    .out(magma_Bits_2_eq_inst0_out)
);
wire [1:0] magma_Bits_2_eq_inst1_in1;
assign magma_Bits_2_eq_inst1_in1 = {inst[53],inst[52]};
coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst1 (
    .in0(const_1_2_out),
    .in1(magma_Bits_2_eq_inst1_in1),
    .out(magma_Bits_2_eq_inst1_out)
);
wire [1:0] magma_Bits_2_eq_inst2_in1;
assign magma_Bits_2_eq_inst2_in1 = {inst[53],inst[52]};
coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst2 (
    .in0(const_2_2_out),
    .in1(magma_Bits_2_eq_inst2_in1),
    .out(magma_Bits_2_eq_inst2_out)
);
wire [1:0] magma_Bits_2_eq_inst3_in1;
assign magma_Bits_2_eq_inst3_in1 = {inst[53],inst[52]};
coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst3 (
    .in0(const_3_2_out),
    .in1(magma_Bits_2_eq_inst3_in1),
    .out(magma_Bits_2_eq_inst3_out)
);
wire [2:0] magma_Bits_3_eq_inst0_in1;
assign magma_Bits_3_eq_inst0_in1 = {inst[68],inst[67],inst[66]};
coreir_eq #(
    .width(3)
) magma_Bits_3_eq_inst0 (
    .in0(const_0_3_out),
    .in1(magma_Bits_3_eq_inst0_in1),
    .out(magma_Bits_3_eq_inst0_out)
);
wire [2:0] magma_Bits_3_eq_inst1_in1;
assign magma_Bits_3_eq_inst1_in1 = {inst[68],inst[67],inst[66]};
coreir_eq #(
    .width(3)
) magma_Bits_3_eq_inst1 (
    .in0(const_1_3_out),
    .in1(magma_Bits_3_eq_inst1_in1),
    .out(magma_Bits_3_eq_inst1_out)
);
wire [2:0] magma_Bits_3_eq_inst2_in1;
assign magma_Bits_3_eq_inst2_in1 = {inst[68],inst[67],inst[66]};
coreir_eq #(
    .width(3)
) magma_Bits_3_eq_inst2 (
    .in0(const_2_3_out),
    .in1(magma_Bits_3_eq_inst2_in1),
    .out(magma_Bits_3_eq_inst2_out)
);
wire [2:0] magma_Bits_3_eq_inst3_in1;
assign magma_Bits_3_eq_inst3_in1 = {inst[68],inst[67],inst[66]};
coreir_eq #(
    .width(3)
) magma_Bits_3_eq_inst3 (
    .in0(const_3_3_out),
    .in1(magma_Bits_3_eq_inst3_in1),
    .out(magma_Bits_3_eq_inst3_out)
);
wire [2:0] magma_Bits_3_eq_inst4_in1;
assign magma_Bits_3_eq_inst4_in1 = {inst[68],inst[67],inst[66]};
coreir_eq #(
    .width(3)
) magma_Bits_3_eq_inst4 (
    .in0(const_4_3_out),
    .in1(magma_Bits_3_eq_inst4_in1),
    .out(magma_Bits_3_eq_inst4_out)
);
wire [3:0] magma_Bits_4_eq_inst0_in1;
assign magma_Bits_4_eq_inst0_in1 = {inst[65],inst[64],inst[63],inst[62]};
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst0 (
    .in0(const_0_4_out),
    .in1(magma_Bits_4_eq_inst0_in1),
    .out(magma_Bits_4_eq_inst0_out)
);
wire [3:0] magma_Bits_4_eq_inst1_in1;
assign magma_Bits_4_eq_inst1_in1 = {inst[65],inst[64],inst[63],inst[62]};
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst1 (
    .in0(const_1_4_out),
    .in1(magma_Bits_4_eq_inst1_in1),
    .out(magma_Bits_4_eq_inst1_out)
);
wire [3:0] magma_Bits_4_eq_inst2_in1;
assign magma_Bits_4_eq_inst2_in1 = {inst[65],inst[64],inst[63],inst[62]};
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst2 (
    .in0(const_2_4_out),
    .in1(magma_Bits_4_eq_inst2_in1),
    .out(magma_Bits_4_eq_inst2_out)
);
wire [3:0] magma_Bits_4_eq_inst3_in1;
assign magma_Bits_4_eq_inst3_in1 = {inst[65],inst[64],inst[63],inst[62]};
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst3 (
    .in0(const_3_4_out),
    .in1(magma_Bits_4_eq_inst3_in1),
    .out(magma_Bits_4_eq_inst3_out)
);
wire [3:0] magma_Bits_4_eq_inst4_in1;
assign magma_Bits_4_eq_inst4_in1 = {inst[65],inst[64],inst[63],inst[62]};
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst4 (
    .in0(const_4_4_out),
    .in1(magma_Bits_4_eq_inst4_in1),
    .out(magma_Bits_4_eq_inst4_out)
);
wire [3:0] magma_Bits_4_eq_inst5_in1;
assign magma_Bits_4_eq_inst5_in1 = {inst[65],inst[64],inst[63],inst[62]};
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst5 (
    .in0(const_5_4_out),
    .in1(magma_Bits_4_eq_inst5_in1),
    .out(magma_Bits_4_eq_inst5_out)
);
wire [3:0] magma_Bits_4_eq_inst6_in1;
assign magma_Bits_4_eq_inst6_in1 = {inst[65],inst[64],inst[63],inst[62]};
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst6 (
    .in0(const_6_4_out),
    .in1(magma_Bits_4_eq_inst6_in1),
    .out(magma_Bits_4_eq_inst6_out)
);
wire [3:0] magma_Bits_4_eq_inst7_in1;
assign magma_Bits_4_eq_inst7_in1 = {inst[65],inst[64],inst[63],inst[62]};
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst7 (
    .in0(const_7_4_out),
    .in1(magma_Bits_4_eq_inst7_in1),
    .out(magma_Bits_4_eq_inst7_out)
);
wire [3:0] magma_Bits_4_eq_inst8_in1;
assign magma_Bits_4_eq_inst8_in1 = {inst[65],inst[64],inst[63],inst[62]};
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst8 (
    .in0(const_8_4_out),
    .in1(magma_Bits_4_eq_inst8_in1),
    .out(magma_Bits_4_eq_inst8_out)
);
assign O = {Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out[0],Mux2xBits16_inst32$coreir_commonlib_mux2x16_inst0$_join_out};
endmodule

module WrappedPE (
    input [80:0] inst,
    input [15:0] inputs0,
    input [15:0] inputs1,
    input [15:0] inputs2,
    input [15:0] inputs3,
    input inputs4,
    input inputs5,
    input inputs6,
    input clk_en,
    output [15:0] O0,
    output O1,
    input CLK,
    input ASYNCRESET
);
wire [16:0] PE_inst0$PE_gen_inst0_O;
wire [80:0] PE_inst0_inst_in;
wire [66:0] PE_inst0$PE_gen_inst0_inputs;
assign PE_inst0$PE_gen_inst0_inputs = {inputs6,inputs5,inputs4,inputs3,inputs2,inputs1,inputs0};
PE_gen PE_inst0$PE_gen_inst0 (
    .inst(PE_inst0_inst_in),
    .inputs(PE_inst0$PE_gen_inst0_inputs),
    .clk_en(clk_en),
    .O(PE_inst0$PE_gen_inst0_O),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
wire [80:0] PE_inst0_inst_out;
assign PE_inst0_inst_out = {inst[80:73],inst[72:69],inst[68:66],inst[65:62],inst[61:54],inst[53:50],inst[49:17],inst[16:15],inst[14:0]};
mantle_wire__typeBitIn81 PE_inst0_inst (
    .in(PE_inst0_inst_in),
    .out(PE_inst0_inst_out)
);
assign O0 = {PE_inst0$PE_gen_inst0_O[15],PE_inst0$PE_gen_inst0_O[14],PE_inst0$PE_gen_inst0_O[13],PE_inst0$PE_gen_inst0_O[12],PE_inst0$PE_gen_inst0_O[11],PE_inst0$PE_gen_inst0_O[10],PE_inst0$PE_gen_inst0_O[9],PE_inst0$PE_gen_inst0_O[8],PE_inst0$PE_gen_inst0_O[7],PE_inst0$PE_gen_inst0_O[6],PE_inst0$PE_gen_inst0_O[5],PE_inst0$PE_gen_inst0_O[4],PE_inst0$PE_gen_inst0_O[3],PE_inst0$PE_gen_inst0_O[2],PE_inst0$PE_gen_inst0_O[1],PE_inst0$PE_gen_inst0_O[0]};
assign O1 = PE_inst0$PE_gen_inst0_O[16];
endmodule

module PE_unq1 (
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    input [15:0] inputs0,
    input [15:0] inputs1,
    input [15:0] inputs2,
    input [15:0] inputs3,
    input [0:0] inputs4,
    input [0:0] inputs5,
    input [0:0] inputs6,
    output [15:0] pe_outputs_0,
    output [0:0] pe_outputs_1,
    output [31:0] read_config_data,
    input reset,
    input [0:0] stall
);
wire [0:0] Invert1_inst0_out;
wire [31:0] MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0_out;
wire [15:0] WrappedPE_inst0_O0;
wire WrappedPE_inst0_O1;
wire [31:0] config_reg_0_O;
wire [31:0] config_reg_1_O;
wire [31:0] config_reg_2_O;
wire [31:0] inst_0_inst0_O;
wire [31:0] inst_1_inst0_O;
wire [31:0] inst_2_inst0_O;
wire [7:0] self_config_config_addr_out;
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(stall),
    .out(Invert1_inst0_out)
);
commonlib_muxn__N3__width32 MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0 (
    .in_data_0(config_reg_0_O),
    .in_data_1(config_reg_1_O),
    .in_data_2(config_reg_2_O),
    .in_sel(self_config_config_addr_out[1:0]),
    .out(MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0_out)
);
wire [80:0] WrappedPE_inst0_inst;
assign WrappedPE_inst0_inst = {inst_2_inst0_O[16:0],inst_1_inst0_O,inst_0_inst0_O};
WrappedPE WrappedPE_inst0 (
    .inst(WrappedPE_inst0_inst),
    .inputs0(inputs0),
    .inputs1(inputs1),
    .inputs2(inputs2),
    .inputs3(inputs3),
    .inputs4(inputs4[0]),
    .inputs5(inputs5[0]),
    .inputs6(inputs6[0]),
    .clk_en(Invert1_inst0_out[0]),
    .O0(WrappedPE_inst0_O0),
    .O1(WrappedPE_inst0_O1),
    .CLK(clk),
    .ASYNCRESET(reset)
);
wire [7:0] config_reg_0_config_addr;
assign config_reg_0_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2],self_config_config_addr_out[1:0]};
ConfigRegister_32_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_reg_0_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_1_config_addr;
assign config_reg_1_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2],self_config_config_addr_out[1:0]};
ConfigRegister_32_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_reg_1_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_2_config_addr;
assign config_reg_2_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2],self_config_config_addr_out[1:0]};
ConfigRegister_32_8_32_2 config_reg_2 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_2_O),
    .config_addr(config_reg_2_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
inst_0 inst_0_inst0 (
    .I(config_reg_0_O),
    .O(inst_0_inst0_O)
);
inst_1 inst_1_inst0 (
    .I(config_reg_1_O),
    .O(inst_1_inst0_O)
);
inst_2 inst_2_inst0 (
    .I(config_reg_2_O),
    .O(inst_2_inst0_O)
);
mantle_wire__typeBit8 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
assign pe_outputs_0 = WrappedPE_inst0_O0;
assign pe_outputs_1 = WrappedPE_inst0_O1;
assign read_config_data = MuxWrapper_3_32_inst0$Mux3xBits32_inst0$coreir_commonlib_mux3x32_inst0_out;
endmodule

module Tile_PE (
    input [0:0] SB_T0_EAST_SB_IN_B1,
    input [15:0] SB_T0_EAST_SB_IN_B16,
    output [0:0] SB_T0_EAST_SB_OUT_B1,
    output [15:0] SB_T0_EAST_SB_OUT_B16,
    input [0:0] SB_T0_NORTH_SB_IN_B1,
    input [15:0] SB_T0_NORTH_SB_IN_B16,
    output [0:0] SB_T0_NORTH_SB_OUT_B1,
    output [15:0] SB_T0_NORTH_SB_OUT_B16,
    input [0:0] SB_T0_SOUTH_SB_IN_B1,
    input [15:0] SB_T0_SOUTH_SB_IN_B16,
    output [0:0] SB_T0_SOUTH_SB_OUT_B1,
    output [15:0] SB_T0_SOUTH_SB_OUT_B16,
    input [0:0] SB_T0_WEST_SB_IN_B1,
    input [15:0] SB_T0_WEST_SB_IN_B16,
    output [0:0] SB_T0_WEST_SB_OUT_B1,
    output [15:0] SB_T0_WEST_SB_OUT_B16,
    input [0:0] SB_T1_EAST_SB_IN_B1,
    input [15:0] SB_T1_EAST_SB_IN_B16,
    output [0:0] SB_T1_EAST_SB_OUT_B1,
    output [15:0] SB_T1_EAST_SB_OUT_B16,
    input [0:0] SB_T1_NORTH_SB_IN_B1,
    input [15:0] SB_T1_NORTH_SB_IN_B16,
    output [0:0] SB_T1_NORTH_SB_OUT_B1,
    output [15:0] SB_T1_NORTH_SB_OUT_B16,
    input [0:0] SB_T1_SOUTH_SB_IN_B1,
    input [15:0] SB_T1_SOUTH_SB_IN_B16,
    output [0:0] SB_T1_SOUTH_SB_OUT_B1,
    output [15:0] SB_T1_SOUTH_SB_OUT_B16,
    input [0:0] SB_T1_WEST_SB_IN_B1,
    input [15:0] SB_T1_WEST_SB_IN_B16,
    output [0:0] SB_T1_WEST_SB_OUT_B1,
    output [15:0] SB_T1_WEST_SB_OUT_B16,
    input [0:0] SB_T2_EAST_SB_IN_B1,
    input [15:0] SB_T2_EAST_SB_IN_B16,
    output [0:0] SB_T2_EAST_SB_OUT_B1,
    output [15:0] SB_T2_EAST_SB_OUT_B16,
    input [0:0] SB_T2_NORTH_SB_IN_B1,
    input [15:0] SB_T2_NORTH_SB_IN_B16,
    output [0:0] SB_T2_NORTH_SB_OUT_B1,
    output [15:0] SB_T2_NORTH_SB_OUT_B16,
    input [0:0] SB_T2_SOUTH_SB_IN_B1,
    input [15:0] SB_T2_SOUTH_SB_IN_B16,
    output [0:0] SB_T2_SOUTH_SB_OUT_B1,
    output [15:0] SB_T2_SOUTH_SB_OUT_B16,
    input [0:0] SB_T2_WEST_SB_IN_B1,
    input [15:0] SB_T2_WEST_SB_IN_B16,
    output [0:0] SB_T2_WEST_SB_OUT_B1,
    output [15:0] SB_T2_WEST_SB_OUT_B16,
    input [0:0] SB_T3_EAST_SB_IN_B1,
    input [15:0] SB_T3_EAST_SB_IN_B16,
    output [0:0] SB_T3_EAST_SB_OUT_B1,
    output [15:0] SB_T3_EAST_SB_OUT_B16,
    input [0:0] SB_T3_NORTH_SB_IN_B1,
    input [15:0] SB_T3_NORTH_SB_IN_B16,
    output [0:0] SB_T3_NORTH_SB_OUT_B1,
    output [15:0] SB_T3_NORTH_SB_OUT_B16,
    input [0:0] SB_T3_SOUTH_SB_IN_B1,
    input [15:0] SB_T3_SOUTH_SB_IN_B16,
    output [0:0] SB_T3_SOUTH_SB_OUT_B1,
    output [15:0] SB_T3_SOUTH_SB_OUT_B16,
    input [0:0] SB_T3_WEST_SB_IN_B1,
    input [15:0] SB_T3_WEST_SB_IN_B16,
    output [0:0] SB_T3_WEST_SB_OUT_B1,
    output [15:0] SB_T3_WEST_SB_OUT_B16,
    input [0:0] SB_T4_EAST_SB_IN_B1,
    input [15:0] SB_T4_EAST_SB_IN_B16,
    output [0:0] SB_T4_EAST_SB_OUT_B1,
    output [15:0] SB_T4_EAST_SB_OUT_B16,
    input [0:0] SB_T4_NORTH_SB_IN_B1,
    input [15:0] SB_T4_NORTH_SB_IN_B16,
    output [0:0] SB_T4_NORTH_SB_OUT_B1,
    output [15:0] SB_T4_NORTH_SB_OUT_B16,
    input [0:0] SB_T4_SOUTH_SB_IN_B1,
    input [15:0] SB_T4_SOUTH_SB_IN_B16,
    output [0:0] SB_T4_SOUTH_SB_OUT_B1,
    output [15:0] SB_T4_SOUTH_SB_OUT_B16,
    input [0:0] SB_T4_WEST_SB_IN_B1,
    input [15:0] SB_T4_WEST_SB_IN_B16,
    output [0:0] SB_T4_WEST_SB_OUT_B1,
    output [15:0] SB_T4_WEST_SB_OUT_B16,
    input clk,
    output clk_out,
    input clk_pass_through,
    output clk_pass_through_out_bot,
    output clk_pass_through_out_right,
    input [31:0] config_config_addr,
    input [31:0] config_config_data,
    output [31:0] config_out_config_addr,
    output [31:0] config_out_config_data,
    output [0:0] config_out_read,
    output [0:0] config_out_write,
    input [0:0] config_read,
    input [0:0] config_write,
    input [0:0] flush,
    output [0:0] flush_out,
    output [8:0] hi,
    output [7:0] lo,
    output [31:0] read_config_data,
    input [31:0] read_config_data_in,
    input reset,
    output reset_out,
    input [0:0] stall,
    output [0:0] stall_out,
    input [15:0] tile_id
);
wire [15:0] CB_data_in_pond_O;
wire [31:0] CB_data_in_pond_read_config_data;
wire [0:0] CB_flush_O;
wire [31:0] CB_flush_read_config_data;
wire [15:0] CB_inputs0_O;
wire [31:0] CB_inputs0_read_config_data;
wire [15:0] CB_inputs1_O;
wire [31:0] CB_inputs1_read_config_data;
wire [15:0] CB_inputs2_O;
wire [31:0] CB_inputs2_read_config_data;
wire [15:0] CB_inputs3_O;
wire [31:0] CB_inputs3_read_config_data;
wire [0:0] CB_inputs4_O;
wire [31:0] CB_inputs4_read_config_data;
wire [0:0] CB_inputs5_O;
wire [31:0] CB_inputs5_read_config_data;
wire [0:0] CB_inputs6_O;
wire [31:0] CB_inputs6_read_config_data;
wire DECODE_FEATURE_0_O;
wire DECODE_FEATURE_1_O;
wire DECODE_FEATURE_10_O;
wire DECODE_FEATURE_11_O;
wire DECODE_FEATURE_12_O;
wire DECODE_FEATURE_13_O;
wire DECODE_FEATURE_14_O;
wire DECODE_FEATURE_2_O;
wire DECODE_FEATURE_3_O;
wire DECODE_FEATURE_4_O;
wire DECODE_FEATURE_5_O;
wire DECODE_FEATURE_6_O;
wire DECODE_FEATURE_7_O;
wire DECODE_FEATURE_8_O;
wire DECODE_FEATURE_9_O;
wire FEATURE_AND_0_out;
wire FEATURE_AND_1_out;
wire FEATURE_AND_10_out;
wire FEATURE_AND_11_out;
wire FEATURE_AND_12_out;
wire FEATURE_AND_13_out;
wire FEATURE_AND_14_out;
wire FEATURE_AND_2_out;
wire FEATURE_AND_3_out;
wire FEATURE_AND_4_out;
wire FEATURE_AND_5_out;
wire FEATURE_AND_6_out;
wire FEATURE_AND_7_out;
wire FEATURE_AND_8_out;
wire FEATURE_AND_9_out;
wire [15:0] PE_inst0_pe_outputs_0;
wire [0:0] PE_inst0_pe_outputs_1;
wire [31:0] PE_inst0_read_config_data;
wire [15:0] PondCore_inst0_data_out_pond;
wire [31:0] PondCore_inst0_read_config_data;
wire [31:0] PondCore_inst0_read_config_data_1;
wire [0:0] PondCore_inst0_valid_out_pond;
wire [0:0] PowerDomainConfigReg_inst0_ps_en_out;
wire [31:0] PowerDomainConfigReg_inst0_read_config_data;
wire [31:0] PowerDomainOR_O;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T0_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T0_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T0_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T0_WEST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T1_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T1_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T1_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T1_WEST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T2_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T2_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T2_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T2_WEST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T3_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T3_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T3_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T3_WEST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T4_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T4_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T4_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T4_WEST_SB_OUT_B16;
wire [31:0] SB_ID0_5TRACKS_B16_PE_read_config_data;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1;
wire [31:0] SB_ID0_5TRACKS_B1_PE_read_config_data;
wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T3_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T3_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T3_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T3_WEST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T4_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T4_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T4_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T4_WEST_SB_IN_B16_O;
wire and_inst0_out;
wire and_inst1_out;
wire [7:0] const_0_8_out;
wire [8:0] const_511_9_out;
wire coreir_eq_16_inst0_out;
wire coreir_wrapOutClock_inst0_out;
wire coreir_wrapOutClock_inst1_out;
wire [31:0] read_data_mux_O;
wire [7:0] CB_data_in_pond_config_config_addr;
assign CB_data_in_pond_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
CB_data_in_pond CB_data_in_pond (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .O(CB_data_in_pond_O),
    .clk(clk),
    .config_config_addr(CB_data_in_pond_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_3_out),
    .read_config_data(CB_data_in_pond_read_config_data),
    .reset(reset)
);
wire [7:0] CB_flush_config_config_addr;
assign CB_flush_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
CB_flush CB_flush (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .O(CB_flush_O),
    .clk(clk),
    .config_config_addr(CB_flush_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_4_out),
    .read_config_data(CB_flush_read_config_data),
    .reset(reset)
);
wire [7:0] CB_inputs0_config_config_addr;
assign CB_inputs0_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
CB_inputs0 CB_inputs0 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .O(CB_inputs0_O),
    .clk(clk),
    .config_config_addr(CB_inputs0_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_5_out),
    .read_config_data(CB_inputs0_read_config_data),
    .reset(reset)
);
wire [7:0] CB_inputs1_config_config_addr;
assign CB_inputs1_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
CB_inputs1 CB_inputs1 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .O(CB_inputs1_O),
    .clk(clk),
    .config_config_addr(CB_inputs1_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_6_out),
    .read_config_data(CB_inputs1_read_config_data),
    .reset(reset)
);
wire [7:0] CB_inputs2_config_config_addr;
assign CB_inputs2_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
CB_inputs2 CB_inputs2 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .O(CB_inputs2_O),
    .clk(clk),
    .config_config_addr(CB_inputs2_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_7_out),
    .read_config_data(CB_inputs2_read_config_data),
    .reset(reset)
);
wire [7:0] CB_inputs3_config_config_addr;
assign CB_inputs3_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
CB_inputs3 CB_inputs3 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .O(CB_inputs3_O),
    .clk(clk),
    .config_config_addr(CB_inputs3_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_8_out),
    .read_config_data(CB_inputs3_read_config_data),
    .reset(reset)
);
wire [7:0] CB_inputs4_config_config_addr;
assign CB_inputs4_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
CB_inputs4 CB_inputs4 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .O(CB_inputs4_O),
    .clk(clk),
    .config_config_addr(CB_inputs4_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_9_out),
    .read_config_data(CB_inputs4_read_config_data),
    .reset(reset)
);
wire [7:0] CB_inputs5_config_config_addr;
assign CB_inputs5_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
CB_inputs5 CB_inputs5 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .O(CB_inputs5_O),
    .clk(clk),
    .config_config_addr(CB_inputs5_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_10_out),
    .read_config_data(CB_inputs5_read_config_data),
    .reset(reset)
);
wire [7:0] CB_inputs6_config_config_addr;
assign CB_inputs6_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
CB_inputs6 CB_inputs6 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .O(CB_inputs6_O),
    .clk(clk),
    .config_config_addr(CB_inputs6_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_11_out),
    .read_config_data(CB_inputs6_read_config_data),
    .reset(reset)
);
wire [7:0] DECODE_FEATURE_0_I;
assign DECODE_FEATURE_0_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode08 DECODE_FEATURE_0 (
    .I(DECODE_FEATURE_0_I),
    .O(DECODE_FEATURE_0_O)
);
wire [7:0] DECODE_FEATURE_1_I;
assign DECODE_FEATURE_1_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode18 DECODE_FEATURE_1 (
    .I(DECODE_FEATURE_1_I),
    .O(DECODE_FEATURE_1_O)
);
wire [7:0] DECODE_FEATURE_10_I;
assign DECODE_FEATURE_10_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode108 DECODE_FEATURE_10 (
    .I(DECODE_FEATURE_10_I),
    .O(DECODE_FEATURE_10_O)
);
wire [7:0] DECODE_FEATURE_11_I;
assign DECODE_FEATURE_11_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode118 DECODE_FEATURE_11 (
    .I(DECODE_FEATURE_11_I),
    .O(DECODE_FEATURE_11_O)
);
wire [7:0] DECODE_FEATURE_12_I;
assign DECODE_FEATURE_12_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode128 DECODE_FEATURE_12 (
    .I(DECODE_FEATURE_12_I),
    .O(DECODE_FEATURE_12_O)
);
wire [7:0] DECODE_FEATURE_13_I;
assign DECODE_FEATURE_13_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode138 DECODE_FEATURE_13 (
    .I(DECODE_FEATURE_13_I),
    .O(DECODE_FEATURE_13_O)
);
wire [7:0] DECODE_FEATURE_14_I;
assign DECODE_FEATURE_14_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode148 DECODE_FEATURE_14 (
    .I(DECODE_FEATURE_14_I),
    .O(DECODE_FEATURE_14_O)
);
wire [7:0] DECODE_FEATURE_2_I;
assign DECODE_FEATURE_2_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode28 DECODE_FEATURE_2 (
    .I(DECODE_FEATURE_2_I),
    .O(DECODE_FEATURE_2_O)
);
wire [7:0] DECODE_FEATURE_3_I;
assign DECODE_FEATURE_3_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode38 DECODE_FEATURE_3 (
    .I(DECODE_FEATURE_3_I),
    .O(DECODE_FEATURE_3_O)
);
wire [7:0] DECODE_FEATURE_4_I;
assign DECODE_FEATURE_4_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode48 DECODE_FEATURE_4 (
    .I(DECODE_FEATURE_4_I),
    .O(DECODE_FEATURE_4_O)
);
wire [7:0] DECODE_FEATURE_5_I;
assign DECODE_FEATURE_5_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode58 DECODE_FEATURE_5 (
    .I(DECODE_FEATURE_5_I),
    .O(DECODE_FEATURE_5_O)
);
wire [7:0] DECODE_FEATURE_6_I;
assign DECODE_FEATURE_6_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode68 DECODE_FEATURE_6 (
    .I(DECODE_FEATURE_6_I),
    .O(DECODE_FEATURE_6_O)
);
wire [7:0] DECODE_FEATURE_7_I;
assign DECODE_FEATURE_7_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode78 DECODE_FEATURE_7 (
    .I(DECODE_FEATURE_7_I),
    .O(DECODE_FEATURE_7_O)
);
wire [7:0] DECODE_FEATURE_8_I;
assign DECODE_FEATURE_8_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode88 DECODE_FEATURE_8 (
    .I(DECODE_FEATURE_8_I),
    .O(DECODE_FEATURE_8_O)
);
wire [7:0] DECODE_FEATURE_9_I;
assign DECODE_FEATURE_9_I = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
Decode98 DECODE_FEATURE_9 (
    .I(DECODE_FEATURE_9_I),
    .O(DECODE_FEATURE_9_O)
);
corebit_and FEATURE_AND_0 (
    .in0(DECODE_FEATURE_0_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_0_out)
);
corebit_and FEATURE_AND_1 (
    .in0(DECODE_FEATURE_1_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_1_out)
);
corebit_and FEATURE_AND_10 (
    .in0(DECODE_FEATURE_10_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_10_out)
);
corebit_and FEATURE_AND_11 (
    .in0(DECODE_FEATURE_11_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_11_out)
);
corebit_and FEATURE_AND_12 (
    .in0(DECODE_FEATURE_12_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_12_out)
);
corebit_and FEATURE_AND_13 (
    .in0(DECODE_FEATURE_13_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_13_out)
);
corebit_and FEATURE_AND_14 (
    .in0(DECODE_FEATURE_14_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_14_out)
);
corebit_and FEATURE_AND_2 (
    .in0(DECODE_FEATURE_2_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_2_out)
);
corebit_and FEATURE_AND_3 (
    .in0(DECODE_FEATURE_3_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_3_out)
);
corebit_and FEATURE_AND_4 (
    .in0(DECODE_FEATURE_4_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_4_out)
);
corebit_and FEATURE_AND_5 (
    .in0(DECODE_FEATURE_5_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_5_out)
);
corebit_and FEATURE_AND_6 (
    .in0(DECODE_FEATURE_6_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_6_out)
);
corebit_and FEATURE_AND_7 (
    .in0(DECODE_FEATURE_7_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_7_out)
);
corebit_and FEATURE_AND_8 (
    .in0(DECODE_FEATURE_8_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_8_out)
);
corebit_and FEATURE_AND_9 (
    .in0(DECODE_FEATURE_9_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_9_out)
);
wire [7:0] PE_inst0_config_config_addr;
assign PE_inst0_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
PE_unq1 PE_inst0 (
    .clk(clk),
    .config_config_addr(PE_inst0_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_0_out),
    .inputs0(CB_inputs0_O),
    .inputs1(CB_inputs1_O),
    .inputs2(CB_inputs2_O),
    .inputs3(CB_inputs3_O),
    .inputs4(CB_inputs4_O),
    .inputs5(CB_inputs5_O),
    .inputs6(CB_inputs6_O),
    .pe_outputs_0(PE_inst0_pe_outputs_0),
    .pe_outputs_1(PE_inst0_pe_outputs_1),
    .read_config_data(PE_inst0_read_config_data),
    .reset(reset),
    .stall(stall)
);
wire [7:0] PondCore_inst0_config_1_config_addr;
assign PondCore_inst0_config_1_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
wire [7:0] PondCore_inst0_config_config_addr;
assign PondCore_inst0_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
PondCore PondCore_inst0 (
    .clk(clk),
    .config_1_config_addr(PondCore_inst0_config_1_config_addr),
    .config_1_config_data(config_config_data),
    .config_1_read(config_read),
    .config_1_write(FEATURE_AND_2_out),
    .config_config_addr(PondCore_inst0_config_config_addr),
    .config_config_data(config_config_data),
    .config_en_0(DECODE_FEATURE_2_O),
    .config_read(config_read),
    .config_write(FEATURE_AND_1_out),
    .data_in_pond(CB_data_in_pond_O),
    .data_out_pond(PondCore_inst0_data_out_pond),
    .flush(CB_flush_O),
    .flush_core(flush),
    .read_config_data(PondCore_inst0_read_config_data),
    .read_config_data_1(PondCore_inst0_read_config_data_1),
    .reset(reset),
    .stall(stall),
    .valid_out_pond(PondCore_inst0_valid_out_pond)
);
wire [7:0] PowerDomainConfigReg_inst0_config_config_addr;
assign PowerDomainConfigReg_inst0_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
PowerDomainConfigReg PowerDomainConfigReg_inst0 (
    .clk(clk),
    .config_config_addr(PowerDomainConfigReg_inst0_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_14_out),
    .ps_en_out(PowerDomainConfigReg_inst0_ps_en_out),
    .read_config_data(PowerDomainConfigReg_inst0_read_config_data),
    .reset(reset)
);
PowerDomainOR PowerDomainOR (
    .I0(read_data_mux_O),
    .I1(read_config_data_in),
    .O(PowerDomainOR_O),
    .I_not(PowerDomainConfigReg_inst0_ps_en_out)
);
wire [7:0] SB_ID0_5TRACKS_B16_PE_config_config_addr;
assign SB_ID0_5TRACKS_B16_PE_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
SB_ID0_5TRACKS_B16_PE SB_ID0_5TRACKS_B16_PE (
    .SB_T0_EAST_SB_IN_B16(SB_T0_EAST_SB_IN_B16),
    .SB_T0_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B16(SB_T0_NORTH_SB_IN_B16),
    .SB_T0_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B16(SB_T0_SOUTH_SB_IN_B16),
    .SB_T0_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B16(SB_T0_WEST_SB_IN_B16),
    .SB_T0_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B16(SB_T1_EAST_SB_IN_B16),
    .SB_T1_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B16(SB_T1_NORTH_SB_IN_B16),
    .SB_T1_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B16(SB_T1_SOUTH_SB_IN_B16),
    .SB_T1_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B16(SB_T1_WEST_SB_IN_B16),
    .SB_T1_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B16(SB_T2_EAST_SB_IN_B16),
    .SB_T2_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B16(SB_T2_NORTH_SB_IN_B16),
    .SB_T2_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B16(SB_T2_SOUTH_SB_IN_B16),
    .SB_T2_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B16(SB_T2_WEST_SB_IN_B16),
    .SB_T2_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B16(SB_T3_EAST_SB_IN_B16),
    .SB_T3_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B16(SB_T3_NORTH_SB_IN_B16),
    .SB_T3_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B16(SB_T3_SOUTH_SB_IN_B16),
    .SB_T3_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B16(SB_T3_WEST_SB_IN_B16),
    .SB_T3_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B16(SB_T4_EAST_SB_IN_B16),
    .SB_T4_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B16(SB_T4_NORTH_SB_IN_B16),
    .SB_T4_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B16(SB_T4_SOUTH_SB_IN_B16),
    .SB_T4_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B16(SB_T4_WEST_SB_IN_B16),
    .SB_T4_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .config_config_addr(SB_ID0_5TRACKS_B16_PE_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_13_out),
    .data_out_pond(PondCore_inst0_data_out_pond),
    .pe_outputs_0(PE_inst0_pe_outputs_0),
    .read_config_data(SB_ID0_5TRACKS_B16_PE_read_config_data),
    .reset(reset),
    .stall(stall)
);
wire [7:0] SB_ID0_5TRACKS_B1_PE_config_config_addr;
assign SB_ID0_5TRACKS_B1_PE_config_config_addr = {config_config_addr[31],config_config_addr[30],config_config_addr[29],config_config_addr[28],config_config_addr[27],config_config_addr[26],config_config_addr[25],config_config_addr[24]};
SB_ID0_5TRACKS_B1_PE SB_ID0_5TRACKS_B1_PE (
    .SB_T0_EAST_SB_IN_B1(SB_T0_EAST_SB_IN_B1),
    .SB_T0_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B1(SB_T0_NORTH_SB_IN_B1),
    .SB_T0_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B1(SB_T0_SOUTH_SB_IN_B1),
    .SB_T0_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B1(SB_T0_WEST_SB_IN_B1),
    .SB_T0_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B1(SB_T1_EAST_SB_IN_B1),
    .SB_T1_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B1(SB_T1_NORTH_SB_IN_B1),
    .SB_T1_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B1(SB_T1_SOUTH_SB_IN_B1),
    .SB_T1_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B1(SB_T1_WEST_SB_IN_B1),
    .SB_T1_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B1(SB_T2_EAST_SB_IN_B1),
    .SB_T2_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B1(SB_T2_NORTH_SB_IN_B1),
    .SB_T2_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B1(SB_T2_SOUTH_SB_IN_B1),
    .SB_T2_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B1(SB_T2_WEST_SB_IN_B1),
    .SB_T2_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B1(SB_T3_EAST_SB_IN_B1),
    .SB_T3_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B1(SB_T3_NORTH_SB_IN_B1),
    .SB_T3_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B1(SB_T3_SOUTH_SB_IN_B1),
    .SB_T3_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B1(SB_T3_WEST_SB_IN_B1),
    .SB_T3_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B1(SB_T4_EAST_SB_IN_B1),
    .SB_T4_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B1(SB_T4_NORTH_SB_IN_B1),
    .SB_T4_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B1(SB_T4_SOUTH_SB_IN_B1),
    .SB_T4_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B1(SB_T4_WEST_SB_IN_B1),
    .SB_T4_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1),
    .clk(clk),
    .config_config_addr(SB_ID0_5TRACKS_B1_PE_config_config_addr),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_12_out),
    .pe_outputs_1(PE_inst0_pe_outputs_1),
    .read_config_data(SB_ID0_5TRACKS_B1_PE_read_config_data),
    .reset(reset),
    .stall(stall),
    .valid_out_pond(PondCore_inst0_valid_out_pond)
);
MuxWrapper_1_1 WIRE_SB_T0_EAST_SB_IN_B1 (
    .I(SB_T0_EAST_SB_IN_B1),
    .O(WIRE_SB_T0_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T0_EAST_SB_IN_B16 (
    .I(SB_T0_EAST_SB_IN_B16),
    .O(WIRE_SB_T0_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T0_NORTH_SB_IN_B1 (
    .I(SB_T0_NORTH_SB_IN_B1),
    .O(WIRE_SB_T0_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T0_NORTH_SB_IN_B16 (
    .I(SB_T0_NORTH_SB_IN_B16),
    .O(WIRE_SB_T0_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T0_SOUTH_SB_IN_B1 (
    .I(SB_T0_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T0_SOUTH_SB_IN_B16 (
    .I(SB_T0_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T0_WEST_SB_IN_B1 (
    .I(SB_T0_WEST_SB_IN_B1),
    .O(WIRE_SB_T0_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T0_WEST_SB_IN_B16 (
    .I(SB_T0_WEST_SB_IN_B16),
    .O(WIRE_SB_T0_WEST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T1_EAST_SB_IN_B1 (
    .I(SB_T1_EAST_SB_IN_B1),
    .O(WIRE_SB_T1_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T1_EAST_SB_IN_B16 (
    .I(SB_T1_EAST_SB_IN_B16),
    .O(WIRE_SB_T1_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T1_NORTH_SB_IN_B1 (
    .I(SB_T1_NORTH_SB_IN_B1),
    .O(WIRE_SB_T1_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T1_NORTH_SB_IN_B16 (
    .I(SB_T1_NORTH_SB_IN_B16),
    .O(WIRE_SB_T1_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T1_SOUTH_SB_IN_B1 (
    .I(SB_T1_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T1_SOUTH_SB_IN_B16 (
    .I(SB_T1_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T1_WEST_SB_IN_B1 (
    .I(SB_T1_WEST_SB_IN_B1),
    .O(WIRE_SB_T1_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T1_WEST_SB_IN_B16 (
    .I(SB_T1_WEST_SB_IN_B16),
    .O(WIRE_SB_T1_WEST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T2_EAST_SB_IN_B1 (
    .I(SB_T2_EAST_SB_IN_B1),
    .O(WIRE_SB_T2_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T2_EAST_SB_IN_B16 (
    .I(SB_T2_EAST_SB_IN_B16),
    .O(WIRE_SB_T2_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T2_NORTH_SB_IN_B1 (
    .I(SB_T2_NORTH_SB_IN_B1),
    .O(WIRE_SB_T2_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T2_NORTH_SB_IN_B16 (
    .I(SB_T2_NORTH_SB_IN_B16),
    .O(WIRE_SB_T2_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T2_SOUTH_SB_IN_B1 (
    .I(SB_T2_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T2_SOUTH_SB_IN_B16 (
    .I(SB_T2_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T2_WEST_SB_IN_B1 (
    .I(SB_T2_WEST_SB_IN_B1),
    .O(WIRE_SB_T2_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T2_WEST_SB_IN_B16 (
    .I(SB_T2_WEST_SB_IN_B16),
    .O(WIRE_SB_T2_WEST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T3_EAST_SB_IN_B1 (
    .I(SB_T3_EAST_SB_IN_B1),
    .O(WIRE_SB_T3_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T3_EAST_SB_IN_B16 (
    .I(SB_T3_EAST_SB_IN_B16),
    .O(WIRE_SB_T3_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T3_NORTH_SB_IN_B1 (
    .I(SB_T3_NORTH_SB_IN_B1),
    .O(WIRE_SB_T3_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T3_NORTH_SB_IN_B16 (
    .I(SB_T3_NORTH_SB_IN_B16),
    .O(WIRE_SB_T3_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T3_SOUTH_SB_IN_B1 (
    .I(SB_T3_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T3_SOUTH_SB_IN_B16 (
    .I(SB_T3_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T3_WEST_SB_IN_B1 (
    .I(SB_T3_WEST_SB_IN_B1),
    .O(WIRE_SB_T3_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T3_WEST_SB_IN_B16 (
    .I(SB_T3_WEST_SB_IN_B16),
    .O(WIRE_SB_T3_WEST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T4_EAST_SB_IN_B1 (
    .I(SB_T4_EAST_SB_IN_B1),
    .O(WIRE_SB_T4_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T4_EAST_SB_IN_B16 (
    .I(SB_T4_EAST_SB_IN_B16),
    .O(WIRE_SB_T4_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T4_NORTH_SB_IN_B1 (
    .I(SB_T4_NORTH_SB_IN_B1),
    .O(WIRE_SB_T4_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T4_NORTH_SB_IN_B16 (
    .I(SB_T4_NORTH_SB_IN_B16),
    .O(WIRE_SB_T4_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T4_SOUTH_SB_IN_B1 (
    .I(SB_T4_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T4_SOUTH_SB_IN_B16 (
    .I(SB_T4_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T4_WEST_SB_IN_B1 (
    .I(SB_T4_WEST_SB_IN_B1),
    .O(WIRE_SB_T4_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T4_WEST_SB_IN_B16 (
    .I(SB_T4_WEST_SB_IN_B16),
    .O(WIRE_SB_T4_WEST_SB_IN_B16_O)
);
corebit_and and_inst0 (
    .in0(coreir_eq_16_inst0_out),
    .in1(config_read[0]),
    .out(and_inst0_out)
);
corebit_and and_inst1 (
    .in0(coreir_eq_16_inst0_out),
    .in1(config_write[0]),
    .out(and_inst1_out)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
coreir_const #(
    .value(9'h1ff),
    .width(9)
) const_511_9 (
    .out(const_511_9_out)
);
wire [15:0] coreir_eq_16_inst0_in1;
assign coreir_eq_16_inst0_in1 = {config_config_addr[15],config_config_addr[14],config_config_addr[13],config_config_addr[12],config_config_addr[11],config_config_addr[10],config_config_addr[9],config_config_addr[8],config_config_addr[7],config_config_addr[6],config_config_addr[5],config_config_addr[4],config_config_addr[3],config_config_addr[2],config_config_addr[1],config_config_addr[0]};
coreir_eq #(
    .width(16)
) coreir_eq_16_inst0 (
    .in0(tile_id),
    .in1(coreir_eq_16_inst0_in1),
    .out(coreir_eq_16_inst0_out)
);
coreir_wrap coreir_wrapOutClock_inst0 (
    .in(clk_pass_through),
    .out(coreir_wrapOutClock_inst0_out)
);
coreir_wrap coreir_wrapOutClock_inst1 (
    .in(clk_pass_through),
    .out(coreir_wrapOutClock_inst1_out)
);
wire [7:0] read_data_mux_S;
assign read_data_mux_S = {config_config_addr[23],config_config_addr[22],config_config_addr[21],config_config_addr[20],config_config_addr[19],config_config_addr[18],config_config_addr[17],config_config_addr[16]};
MuxWithDefaultWrapper_15_32_8_0 read_data_mux (
    .EN(and_inst0_out),
    .I_0(PE_inst0_read_config_data),
    .I_1(PondCore_inst0_read_config_data),
    .I_10(CB_inputs5_read_config_data),
    .I_11(CB_inputs6_read_config_data),
    .I_12(SB_ID0_5TRACKS_B1_PE_read_config_data),
    .I_13(SB_ID0_5TRACKS_B16_PE_read_config_data),
    .I_14(PowerDomainConfigReg_inst0_read_config_data),
    .I_2(PondCore_inst0_read_config_data_1),
    .I_3(CB_data_in_pond_read_config_data),
    .I_4(CB_flush_read_config_data),
    .I_5(CB_inputs0_read_config_data),
    .I_6(CB_inputs1_read_config_data),
    .I_7(CB_inputs2_read_config_data),
    .I_8(CB_inputs3_read_config_data),
    .I_9(CB_inputs4_read_config_data),
    .O(read_data_mux_O),
    .S(read_data_mux_S)
);
assign SB_T0_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1;
assign SB_T0_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T0_EAST_SB_OUT_B16;
assign SB_T0_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1;
assign SB_T0_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T0_NORTH_SB_OUT_B16;
assign SB_T0_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1;
assign SB_T0_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T0_SOUTH_SB_OUT_B16;
assign SB_T0_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1;
assign SB_T0_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T0_WEST_SB_OUT_B16;
assign SB_T1_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1;
assign SB_T1_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T1_EAST_SB_OUT_B16;
assign SB_T1_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1;
assign SB_T1_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T1_NORTH_SB_OUT_B16;
assign SB_T1_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1;
assign SB_T1_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T1_SOUTH_SB_OUT_B16;
assign SB_T1_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1;
assign SB_T1_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T1_WEST_SB_OUT_B16;
assign SB_T2_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1;
assign SB_T2_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T2_EAST_SB_OUT_B16;
assign SB_T2_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1;
assign SB_T2_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T2_NORTH_SB_OUT_B16;
assign SB_T2_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1;
assign SB_T2_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T2_SOUTH_SB_OUT_B16;
assign SB_T2_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1;
assign SB_T2_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T2_WEST_SB_OUT_B16;
assign SB_T3_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1;
assign SB_T3_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T3_EAST_SB_OUT_B16;
assign SB_T3_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1;
assign SB_T3_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T3_NORTH_SB_OUT_B16;
assign SB_T3_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1;
assign SB_T3_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T3_SOUTH_SB_OUT_B16;
assign SB_T3_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1;
assign SB_T3_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T3_WEST_SB_OUT_B16;
assign SB_T4_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1;
assign SB_T4_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T4_EAST_SB_OUT_B16;
assign SB_T4_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1;
assign SB_T4_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T4_NORTH_SB_OUT_B16;
assign SB_T4_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1;
assign SB_T4_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T4_SOUTH_SB_OUT_B16;
assign SB_T4_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1;
assign SB_T4_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T4_WEST_SB_OUT_B16;
assign clk_out = coreir_wrapOutClock_inst0_out;
assign clk_pass_through_out_bot = clk_pass_through;
assign clk_pass_through_out_right = coreir_wrapOutClock_inst1_out;
assign config_out_config_addr = config_config_addr;
assign config_out_config_data = config_config_data;
assign config_out_read = config_read;
assign config_out_write = config_write;
assign flush_out = flush;
assign hi = const_511_9_out;
assign lo = const_0_8_out;
assign read_config_data = PowerDomainOR_O;
assign reset_out = reset;
assign stall_out = stall;
endmodule

module Interconnect (
    input clk,
    input [31:0] config_0_config_addr,
    input [31:0] config_0_config_data,
    input [0:0] config_0_read,
    input [0:0] config_0_write,
    input [31:0] config_1_config_addr,
    input [31:0] config_1_config_data,
    input [0:0] config_1_read,
    input [0:0] config_1_write,
    input [31:0] config_2_config_addr,
    input [31:0] config_2_config_data,
    input [0:0] config_2_read,
    input [0:0] config_2_write,
    input [31:0] config_3_config_addr,
    input [31:0] config_3_config_data,
    input [0:0] config_3_read,
    input [0:0] config_3_write,
    input [0:0] flush,
    input [15:0] glb2io_16_X00_Y00,
    input [15:0] glb2io_16_X01_Y00,
    input [15:0] glb2io_16_X02_Y00,
    input [15:0] glb2io_16_X03_Y00,
    input [0:0] glb2io_1_X00_Y00,
    input [0:0] glb2io_1_X01_Y00,
    input [0:0] glb2io_1_X02_Y00,
    input [0:0] glb2io_1_X03_Y00,
    output [15:0] io2glb_16_X00_Y00,
    output [15:0] io2glb_16_X01_Y00,
    output [15:0] io2glb_16_X02_Y00,
    output [15:0] io2glb_16_X03_Y00,
    output [0:0] io2glb_1_X00_Y00,
    output [0:0] io2glb_1_X01_Y00,
    output [0:0] io2glb_1_X02_Y00,
    output [0:0] io2glb_1_X03_Y00,
    output [31:0] read_config_data,
    input reset,
    input [3:0] stall
);
wire [0:0] Tile_X00_Y00_io2glb_1;
wire [0:0] Tile_X00_Y00_io2f_1;
wire [15:0] Tile_X00_Y00_io2glb_16;
wire [15:0] Tile_X00_Y00_io2f_16;
wire [8:0] Tile_X00_Y00_hi;
wire [7:0] Tile_X00_Y00_lo;
wire [0:0] Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y01_clk_out;
wire Tile_X00_Y01_clk_pass_through_out_bot;
wire Tile_X00_Y01_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y01_config_out_config_addr;
wire [31:0] Tile_X00_Y01_config_out_config_data;
wire [0:0] Tile_X00_Y01_config_out_read;
wire [0:0] Tile_X00_Y01_config_out_write;
wire [0:0] Tile_X00_Y01_flush_out;
wire [8:0] Tile_X00_Y01_hi;
wire [7:0] Tile_X00_Y01_lo;
wire [31:0] Tile_X00_Y01_read_config_data;
wire Tile_X00_Y01_reset_out;
wire [0:0] Tile_X00_Y01_stall_out;
wire [0:0] Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y02_clk_out;
wire Tile_X00_Y02_clk_pass_through_out_bot;
wire Tile_X00_Y02_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y02_config_out_config_addr;
wire [31:0] Tile_X00_Y02_config_out_config_data;
wire [0:0] Tile_X00_Y02_config_out_read;
wire [0:0] Tile_X00_Y02_config_out_write;
wire [0:0] Tile_X00_Y02_flush_out;
wire [8:0] Tile_X00_Y02_hi;
wire [7:0] Tile_X00_Y02_lo;
wire [31:0] Tile_X00_Y02_read_config_data;
wire Tile_X00_Y02_reset_out;
wire [0:0] Tile_X00_Y02_stall_out;
wire [0:0] Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y03_clk_out;
wire Tile_X00_Y03_clk_pass_through_out_bot;
wire Tile_X00_Y03_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y03_config_out_config_addr;
wire [31:0] Tile_X00_Y03_config_out_config_data;
wire [0:0] Tile_X00_Y03_config_out_read;
wire [0:0] Tile_X00_Y03_config_out_write;
wire [0:0] Tile_X00_Y03_flush_out;
wire [8:0] Tile_X00_Y03_hi;
wire [7:0] Tile_X00_Y03_lo;
wire [31:0] Tile_X00_Y03_read_config_data;
wire Tile_X00_Y03_reset_out;
wire [0:0] Tile_X00_Y03_stall_out;
wire [0:0] Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y04_clk_out;
wire Tile_X00_Y04_clk_pass_through_out_bot;
wire Tile_X00_Y04_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y04_config_out_config_addr;
wire [31:0] Tile_X00_Y04_config_out_config_data;
wire [0:0] Tile_X00_Y04_config_out_read;
wire [0:0] Tile_X00_Y04_config_out_write;
wire [0:0] Tile_X00_Y04_flush_out;
wire [8:0] Tile_X00_Y04_hi;
wire [7:0] Tile_X00_Y04_lo;
wire [31:0] Tile_X00_Y04_read_config_data;
wire Tile_X00_Y04_reset_out;
wire [0:0] Tile_X00_Y04_stall_out;
wire [0:0] Tile_X01_Y00_io2glb_1;
wire [0:0] Tile_X01_Y00_io2f_1;
wire [15:0] Tile_X01_Y00_io2glb_16;
wire [15:0] Tile_X01_Y00_io2f_16;
wire [8:0] Tile_X01_Y00_hi;
wire [7:0] Tile_X01_Y00_lo;
wire [0:0] Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y01_clk_out;
wire Tile_X01_Y01_clk_pass_through_out_bot;
wire Tile_X01_Y01_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y01_config_out_config_addr;
wire [31:0] Tile_X01_Y01_config_out_config_data;
wire [0:0] Tile_X01_Y01_config_out_read;
wire [0:0] Tile_X01_Y01_config_out_write;
wire [0:0] Tile_X01_Y01_flush_out;
wire [8:0] Tile_X01_Y01_hi;
wire [7:0] Tile_X01_Y01_lo;
wire [31:0] Tile_X01_Y01_read_config_data;
wire Tile_X01_Y01_reset_out;
wire [0:0] Tile_X01_Y01_stall_out;
wire [0:0] Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y02_clk_out;
wire Tile_X01_Y02_clk_pass_through_out_bot;
wire Tile_X01_Y02_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y02_config_out_config_addr;
wire [31:0] Tile_X01_Y02_config_out_config_data;
wire [0:0] Tile_X01_Y02_config_out_read;
wire [0:0] Tile_X01_Y02_config_out_write;
wire [0:0] Tile_X01_Y02_flush_out;
wire [8:0] Tile_X01_Y02_hi;
wire [7:0] Tile_X01_Y02_lo;
wire [31:0] Tile_X01_Y02_read_config_data;
wire Tile_X01_Y02_reset_out;
wire [0:0] Tile_X01_Y02_stall_out;
wire [0:0] Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y03_clk_out;
wire Tile_X01_Y03_clk_pass_through_out_bot;
wire Tile_X01_Y03_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y03_config_out_config_addr;
wire [31:0] Tile_X01_Y03_config_out_config_data;
wire [0:0] Tile_X01_Y03_config_out_read;
wire [0:0] Tile_X01_Y03_config_out_write;
wire [0:0] Tile_X01_Y03_flush_out;
wire [8:0] Tile_X01_Y03_hi;
wire [7:0] Tile_X01_Y03_lo;
wire [31:0] Tile_X01_Y03_read_config_data;
wire Tile_X01_Y03_reset_out;
wire [0:0] Tile_X01_Y03_stall_out;
wire [0:0] Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y04_clk_out;
wire Tile_X01_Y04_clk_pass_through_out_bot;
wire Tile_X01_Y04_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y04_config_out_config_addr;
wire [31:0] Tile_X01_Y04_config_out_config_data;
wire [0:0] Tile_X01_Y04_config_out_read;
wire [0:0] Tile_X01_Y04_config_out_write;
wire [0:0] Tile_X01_Y04_flush_out;
wire [8:0] Tile_X01_Y04_hi;
wire [7:0] Tile_X01_Y04_lo;
wire [31:0] Tile_X01_Y04_read_config_data;
wire Tile_X01_Y04_reset_out;
wire [0:0] Tile_X01_Y04_stall_out;
wire [0:0] Tile_X02_Y00_io2glb_1;
wire [0:0] Tile_X02_Y00_io2f_1;
wire [15:0] Tile_X02_Y00_io2glb_16;
wire [15:0] Tile_X02_Y00_io2f_16;
wire [8:0] Tile_X02_Y00_hi;
wire [7:0] Tile_X02_Y00_lo;
wire [0:0] Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y01_clk_out;
wire Tile_X02_Y01_clk_pass_through_out_bot;
wire Tile_X02_Y01_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y01_config_out_config_addr;
wire [31:0] Tile_X02_Y01_config_out_config_data;
wire [0:0] Tile_X02_Y01_config_out_read;
wire [0:0] Tile_X02_Y01_config_out_write;
wire [0:0] Tile_X02_Y01_flush_out;
wire [8:0] Tile_X02_Y01_hi;
wire [7:0] Tile_X02_Y01_lo;
wire [31:0] Tile_X02_Y01_read_config_data;
wire Tile_X02_Y01_reset_out;
wire [0:0] Tile_X02_Y01_stall_out;
wire [0:0] Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y02_clk_out;
wire Tile_X02_Y02_clk_pass_through_out_bot;
wire Tile_X02_Y02_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y02_config_out_config_addr;
wire [31:0] Tile_X02_Y02_config_out_config_data;
wire [0:0] Tile_X02_Y02_config_out_read;
wire [0:0] Tile_X02_Y02_config_out_write;
wire [0:0] Tile_X02_Y02_flush_out;
wire [8:0] Tile_X02_Y02_hi;
wire [7:0] Tile_X02_Y02_lo;
wire [31:0] Tile_X02_Y02_read_config_data;
wire Tile_X02_Y02_reset_out;
wire [0:0] Tile_X02_Y02_stall_out;
wire [0:0] Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y03_clk_out;
wire Tile_X02_Y03_clk_pass_through_out_bot;
wire Tile_X02_Y03_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y03_config_out_config_addr;
wire [31:0] Tile_X02_Y03_config_out_config_data;
wire [0:0] Tile_X02_Y03_config_out_read;
wire [0:0] Tile_X02_Y03_config_out_write;
wire [0:0] Tile_X02_Y03_flush_out;
wire [8:0] Tile_X02_Y03_hi;
wire [7:0] Tile_X02_Y03_lo;
wire [31:0] Tile_X02_Y03_read_config_data;
wire Tile_X02_Y03_reset_out;
wire [0:0] Tile_X02_Y03_stall_out;
wire [0:0] Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y04_clk_out;
wire Tile_X02_Y04_clk_pass_through_out_bot;
wire Tile_X02_Y04_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y04_config_out_config_addr;
wire [31:0] Tile_X02_Y04_config_out_config_data;
wire [0:0] Tile_X02_Y04_config_out_read;
wire [0:0] Tile_X02_Y04_config_out_write;
wire [0:0] Tile_X02_Y04_flush_out;
wire [8:0] Tile_X02_Y04_hi;
wire [7:0] Tile_X02_Y04_lo;
wire [31:0] Tile_X02_Y04_read_config_data;
wire Tile_X02_Y04_reset_out;
wire [0:0] Tile_X02_Y04_stall_out;
wire [0:0] Tile_X03_Y00_io2glb_1;
wire [0:0] Tile_X03_Y00_io2f_1;
wire [15:0] Tile_X03_Y00_io2glb_16;
wire [15:0] Tile_X03_Y00_io2f_16;
wire [8:0] Tile_X03_Y00_hi;
wire [7:0] Tile_X03_Y00_lo;
wire [0:0] Tile_X03_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y01_clk_out;
wire [31:0] Tile_X03_Y01_config_out_config_addr;
wire [31:0] Tile_X03_Y01_config_out_config_data;
wire [0:0] Tile_X03_Y01_config_out_read;
wire [0:0] Tile_X03_Y01_config_out_write;
wire [0:0] Tile_X03_Y01_flush_out;
wire [8:0] Tile_X03_Y01_hi;
wire [7:0] Tile_X03_Y01_lo;
wire [31:0] Tile_X03_Y01_read_config_data;
wire Tile_X03_Y01_reset_out;
wire [0:0] Tile_X03_Y01_stall_out;
wire [0:0] Tile_X03_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y02_clk_out;
wire [31:0] Tile_X03_Y02_config_out_config_addr;
wire [31:0] Tile_X03_Y02_config_out_config_data;
wire [0:0] Tile_X03_Y02_config_out_read;
wire [0:0] Tile_X03_Y02_config_out_write;
wire [0:0] Tile_X03_Y02_flush_out;
wire [8:0] Tile_X03_Y02_hi;
wire [7:0] Tile_X03_Y02_lo;
wire [31:0] Tile_X03_Y02_read_config_data;
wire Tile_X03_Y02_reset_out;
wire [0:0] Tile_X03_Y02_stall_out;
wire [0:0] Tile_X03_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y03_clk_out;
wire [31:0] Tile_X03_Y03_config_out_config_addr;
wire [31:0] Tile_X03_Y03_config_out_config_data;
wire [0:0] Tile_X03_Y03_config_out_read;
wire [0:0] Tile_X03_Y03_config_out_write;
wire [0:0] Tile_X03_Y03_flush_out;
wire [8:0] Tile_X03_Y03_hi;
wire [7:0] Tile_X03_Y03_lo;
wire [31:0] Tile_X03_Y03_read_config_data;
wire Tile_X03_Y03_reset_out;
wire [0:0] Tile_X03_Y03_stall_out;
wire [0:0] Tile_X03_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y04_clk_out;
wire [31:0] Tile_X03_Y04_config_out_config_addr;
wire [31:0] Tile_X03_Y04_config_out_config_data;
wire [0:0] Tile_X03_Y04_config_out_read;
wire [0:0] Tile_X03_Y04_config_out_write;
wire [0:0] Tile_X03_Y04_flush_out;
wire [8:0] Tile_X03_Y04_hi;
wire [7:0] Tile_X03_Y04_lo;
wire [31:0] Tile_X03_Y04_read_config_data;
wire Tile_X03_Y04_reset_out;
wire [0:0] Tile_X03_Y04_stall_out;
wire [0:0] const_0_1_out;
wire [15:0] const_0_16_out;
wire [31:0] const_0_32_out;
wire coreir_wrapInClock_inst0_out;
wire coreir_wrapInClock_inst1_out;
wire coreir_wrapInClock_inst2_out;
wire [31:0] read_config_data_or_final_O;
wire [3:0] self_stall_out;
wire [15:0] Tile_X00_Y00_tile_id;
assign Tile_X00_Y00_tile_id = {Tile_X00_Y00_lo[7],Tile_X00_Y00_lo[7],Tile_X00_Y00_lo[6],Tile_X00_Y00_lo[6],Tile_X00_Y00_lo[5],Tile_X00_Y00_lo[5],Tile_X00_Y00_lo[4],Tile_X00_Y00_lo[4],Tile_X00_Y00_lo[3],Tile_X00_Y00_lo[3],Tile_X00_Y00_lo[2],Tile_X00_Y00_lo[2],Tile_X00_Y00_lo[1],Tile_X00_Y00_lo[1],Tile_X00_Y00_lo[0],Tile_X00_Y00_lo[0]};
Tile_io_core Tile_X00_Y00 (
    .tile_id(Tile_X00_Y00_tile_id),
    .glb2io_1(glb2io_1_X00_Y00),
    .f2io_1(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X00_Y00_io2glb_1),
    .io2f_1(Tile_X00_Y00_io2f_1),
    .glb2io_16(glb2io_16_X00_Y00),
    .f2io_16(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X00_Y00_io2glb_16),
    .io2f_16(Tile_X00_Y00_io2f_16),
    .hi(Tile_X00_Y00_hi),
    .lo(Tile_X00_Y00_lo)
);
wire [15:0] Tile_X00_Y01_tile_id;
assign Tile_X00_Y01_tile_id = {Tile_X00_Y01_lo[7],Tile_X00_Y01_lo[7],Tile_X00_Y01_lo[6],Tile_X00_Y01_lo[6],Tile_X00_Y01_lo[5],Tile_X00_Y01_lo[5],Tile_X00_Y01_lo[4],Tile_X00_Y01_lo[4],Tile_X00_Y01_lo[3],Tile_X00_Y01_lo[3],Tile_X00_Y01_lo[2],Tile_X00_Y01_lo[2],Tile_X00_Y01_lo[1],Tile_X00_Y01_lo[1],Tile_X00_Y01_lo[0],Tile_X00_Y01_hi[0]};
Tile_PE Tile_X00_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .clk_out(Tile_X00_Y01_clk_out),
    .clk_pass_through(coreir_wrapInClock_inst0_out),
    .clk_pass_through_out_bot(Tile_X00_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y01_clk_pass_through_out_right),
    .config_config_addr(config_0_config_addr),
    .config_config_data(config_0_config_data),
    .config_out_config_addr(Tile_X00_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y01_config_out_config_data),
    .config_out_read(Tile_X00_Y01_config_out_read),
    .config_out_write(Tile_X00_Y01_config_out_write),
    .config_read(config_0_read),
    .config_write(config_0_write),
    .flush(flush),
    .flush_out(Tile_X00_Y01_flush_out),
    .hi(Tile_X00_Y01_hi),
    .lo(Tile_X00_Y01_lo),
    .read_config_data(Tile_X00_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X00_Y01_reset_out),
    .stall(self_stall_out[0:0]),
    .stall_out(Tile_X00_Y01_stall_out),
    .tile_id(Tile_X00_Y01_tile_id)
);
wire [15:0] Tile_X00_Y02_tile_id;
assign Tile_X00_Y02_tile_id = {Tile_X00_Y02_lo[7],Tile_X00_Y02_lo[7],Tile_X00_Y02_lo[6],Tile_X00_Y02_lo[6],Tile_X00_Y02_lo[5],Tile_X00_Y02_lo[5],Tile_X00_Y02_lo[4],Tile_X00_Y02_lo[4],Tile_X00_Y02_lo[3],Tile_X00_Y02_lo[3],Tile_X00_Y02_lo[2],Tile_X00_Y02_lo[2],Tile_X00_Y02_lo[1],Tile_X00_Y02_lo[1],Tile_X00_Y02_hi[1],Tile_X00_Y02_lo[0]};
Tile_PE Tile_X00_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y01_clk_out),
    .clk_out(Tile_X00_Y02_clk_out),
    .clk_pass_through(Tile_X00_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y02_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y01_config_out_config_addr),
    .config_config_data(Tile_X00_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y02_config_out_config_data),
    .config_out_read(Tile_X00_Y02_config_out_read),
    .config_out_write(Tile_X00_Y02_config_out_write),
    .config_read(Tile_X00_Y01_config_out_read),
    .config_write(Tile_X00_Y01_config_out_write),
    .flush(Tile_X00_Y01_flush_out),
    .flush_out(Tile_X00_Y02_flush_out),
    .hi(Tile_X00_Y02_hi),
    .lo(Tile_X00_Y02_lo),
    .read_config_data(Tile_X00_Y02_read_config_data),
    .read_config_data_in(Tile_X00_Y01_read_config_data),
    .reset(Tile_X00_Y01_reset_out),
    .reset_out(Tile_X00_Y02_reset_out),
    .stall(Tile_X00_Y01_stall_out),
    .stall_out(Tile_X00_Y02_stall_out),
    .tile_id(Tile_X00_Y02_tile_id)
);
wire [15:0] Tile_X00_Y03_tile_id;
assign Tile_X00_Y03_tile_id = {Tile_X00_Y03_lo[7],Tile_X00_Y03_lo[7],Tile_X00_Y03_lo[6],Tile_X00_Y03_lo[6],Tile_X00_Y03_lo[5],Tile_X00_Y03_lo[5],Tile_X00_Y03_lo[4],Tile_X00_Y03_lo[4],Tile_X00_Y03_lo[3],Tile_X00_Y03_lo[3],Tile_X00_Y03_lo[2],Tile_X00_Y03_lo[2],Tile_X00_Y03_lo[1],Tile_X00_Y03_lo[1],Tile_X00_Y03_hi[1],Tile_X00_Y03_hi[0]};
Tile_PE Tile_X00_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y02_clk_out),
    .clk_out(Tile_X00_Y03_clk_out),
    .clk_pass_through(Tile_X00_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y03_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y02_config_out_config_addr),
    .config_config_data(Tile_X00_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y03_config_out_config_data),
    .config_out_read(Tile_X00_Y03_config_out_read),
    .config_out_write(Tile_X00_Y03_config_out_write),
    .config_read(Tile_X00_Y02_config_out_read),
    .config_write(Tile_X00_Y02_config_out_write),
    .flush(Tile_X00_Y02_flush_out),
    .flush_out(Tile_X00_Y03_flush_out),
    .hi(Tile_X00_Y03_hi),
    .lo(Tile_X00_Y03_lo),
    .read_config_data(Tile_X00_Y03_read_config_data),
    .read_config_data_in(Tile_X00_Y02_read_config_data),
    .reset(Tile_X00_Y02_reset_out),
    .reset_out(Tile_X00_Y03_reset_out),
    .stall(Tile_X00_Y02_stall_out),
    .stall_out(Tile_X00_Y03_stall_out),
    .tile_id(Tile_X00_Y03_tile_id)
);
wire [15:0] Tile_X00_Y04_tile_id;
assign Tile_X00_Y04_tile_id = {Tile_X00_Y04_lo[7],Tile_X00_Y04_lo[7],Tile_X00_Y04_lo[6],Tile_X00_Y04_lo[6],Tile_X00_Y04_lo[5],Tile_X00_Y04_lo[5],Tile_X00_Y04_lo[4],Tile_X00_Y04_lo[4],Tile_X00_Y04_lo[3],Tile_X00_Y04_lo[3],Tile_X00_Y04_lo[2],Tile_X00_Y04_lo[2],Tile_X00_Y04_lo[1],Tile_X00_Y04_hi[1],Tile_X00_Y04_lo[0],Tile_X00_Y04_lo[0]};
Tile_PE Tile_X00_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y03_clk_out),
    .clk_out(Tile_X00_Y04_clk_out),
    .clk_pass_through(Tile_X00_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y04_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y03_config_out_config_addr),
    .config_config_data(Tile_X00_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y04_config_out_config_data),
    .config_out_read(Tile_X00_Y04_config_out_read),
    .config_out_write(Tile_X00_Y04_config_out_write),
    .config_read(Tile_X00_Y03_config_out_read),
    .config_write(Tile_X00_Y03_config_out_write),
    .flush(Tile_X00_Y03_flush_out),
    .flush_out(Tile_X00_Y04_flush_out),
    .hi(Tile_X00_Y04_hi),
    .lo(Tile_X00_Y04_lo),
    .read_config_data(Tile_X00_Y04_read_config_data),
    .read_config_data_in(Tile_X00_Y03_read_config_data),
    .reset(Tile_X00_Y03_reset_out),
    .reset_out(Tile_X00_Y04_reset_out),
    .stall(Tile_X00_Y03_stall_out),
    .stall_out(Tile_X00_Y04_stall_out),
    .tile_id(Tile_X00_Y04_tile_id)
);
wire [15:0] Tile_X01_Y00_tile_id;
assign Tile_X01_Y00_tile_id = {Tile_X01_Y00_lo[7],Tile_X01_Y00_lo[7],Tile_X01_Y00_lo[6],Tile_X01_Y00_lo[6],Tile_X01_Y00_lo[5],Tile_X01_Y00_lo[5],Tile_X01_Y00_lo[4],Tile_X01_Y00_hi[4],Tile_X01_Y00_lo[3],Tile_X01_Y00_lo[3],Tile_X01_Y00_lo[2],Tile_X01_Y00_lo[2],Tile_X01_Y00_lo[1],Tile_X01_Y00_lo[1],Tile_X01_Y00_lo[0],Tile_X01_Y00_lo[0]};
Tile_io_core Tile_X01_Y00 (
    .tile_id(Tile_X01_Y00_tile_id),
    .glb2io_1(glb2io_1_X01_Y00),
    .f2io_1(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X01_Y00_io2glb_1),
    .io2f_1(Tile_X01_Y00_io2f_1),
    .glb2io_16(glb2io_16_X01_Y00),
    .f2io_16(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X01_Y00_io2glb_16),
    .io2f_16(Tile_X01_Y00_io2f_16),
    .hi(Tile_X01_Y00_hi),
    .lo(Tile_X01_Y00_lo)
);
wire [15:0] Tile_X01_Y01_tile_id;
assign Tile_X01_Y01_tile_id = {Tile_X01_Y01_lo[7],Tile_X01_Y01_lo[7],Tile_X01_Y01_lo[6],Tile_X01_Y01_lo[6],Tile_X01_Y01_lo[5],Tile_X01_Y01_lo[5],Tile_X01_Y01_lo[4],Tile_X01_Y01_hi[4],Tile_X01_Y01_lo[3],Tile_X01_Y01_lo[3],Tile_X01_Y01_lo[2],Tile_X01_Y01_lo[2],Tile_X01_Y01_lo[1],Tile_X01_Y01_lo[1],Tile_X01_Y01_lo[0],Tile_X01_Y01_hi[0]};
Tile_PE Tile_X01_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .clk_out(Tile_X01_Y01_clk_out),
    .clk_pass_through(coreir_wrapInClock_inst1_out),
    .clk_pass_through_out_bot(Tile_X01_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y01_clk_pass_through_out_right),
    .config_config_addr(config_1_config_addr),
    .config_config_data(config_1_config_data),
    .config_out_config_addr(Tile_X01_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y01_config_out_config_data),
    .config_out_read(Tile_X01_Y01_config_out_read),
    .config_out_write(Tile_X01_Y01_config_out_write),
    .config_read(config_1_read),
    .config_write(config_1_write),
    .flush(flush),
    .flush_out(Tile_X01_Y01_flush_out),
    .hi(Tile_X01_Y01_hi),
    .lo(Tile_X01_Y01_lo),
    .read_config_data(Tile_X01_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X01_Y01_reset_out),
    .stall(self_stall_out[1:1]),
    .stall_out(Tile_X01_Y01_stall_out),
    .tile_id(Tile_X01_Y01_tile_id)
);
wire [15:0] Tile_X01_Y02_tile_id;
assign Tile_X01_Y02_tile_id = {Tile_X01_Y02_lo[7],Tile_X01_Y02_lo[7],Tile_X01_Y02_lo[6],Tile_X01_Y02_lo[6],Tile_X01_Y02_lo[5],Tile_X01_Y02_lo[5],Tile_X01_Y02_lo[4],Tile_X01_Y02_hi[4],Tile_X01_Y02_lo[3],Tile_X01_Y02_lo[3],Tile_X01_Y02_lo[2],Tile_X01_Y02_lo[2],Tile_X01_Y02_lo[1],Tile_X01_Y02_lo[1],Tile_X01_Y02_hi[1],Tile_X01_Y02_lo[0]};
Tile_PE Tile_X01_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y01_clk_out),
    .clk_out(Tile_X01_Y02_clk_out),
    .clk_pass_through(Tile_X01_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y02_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y01_config_out_config_addr),
    .config_config_data(Tile_X01_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y02_config_out_config_data),
    .config_out_read(Tile_X01_Y02_config_out_read),
    .config_out_write(Tile_X01_Y02_config_out_write),
    .config_read(Tile_X01_Y01_config_out_read),
    .config_write(Tile_X01_Y01_config_out_write),
    .flush(Tile_X01_Y01_flush_out),
    .flush_out(Tile_X01_Y02_flush_out),
    .hi(Tile_X01_Y02_hi),
    .lo(Tile_X01_Y02_lo),
    .read_config_data(Tile_X01_Y02_read_config_data),
    .read_config_data_in(Tile_X01_Y01_read_config_data),
    .reset(Tile_X01_Y01_reset_out),
    .reset_out(Tile_X01_Y02_reset_out),
    .stall(Tile_X01_Y01_stall_out),
    .stall_out(Tile_X01_Y02_stall_out),
    .tile_id(Tile_X01_Y02_tile_id)
);
wire [15:0] Tile_X01_Y03_tile_id;
assign Tile_X01_Y03_tile_id = {Tile_X01_Y03_lo[7],Tile_X01_Y03_lo[7],Tile_X01_Y03_lo[6],Tile_X01_Y03_lo[6],Tile_X01_Y03_lo[5],Tile_X01_Y03_lo[5],Tile_X01_Y03_lo[4],Tile_X01_Y03_hi[4],Tile_X01_Y03_lo[3],Tile_X01_Y03_lo[3],Tile_X01_Y03_lo[2],Tile_X01_Y03_lo[2],Tile_X01_Y03_lo[1],Tile_X01_Y03_lo[1],Tile_X01_Y03_hi[1],Tile_X01_Y03_hi[0]};
Tile_PE Tile_X01_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y02_clk_out),
    .clk_out(Tile_X01_Y03_clk_out),
    .clk_pass_through(Tile_X01_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y03_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y02_config_out_config_addr),
    .config_config_data(Tile_X01_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y03_config_out_config_data),
    .config_out_read(Tile_X01_Y03_config_out_read),
    .config_out_write(Tile_X01_Y03_config_out_write),
    .config_read(Tile_X01_Y02_config_out_read),
    .config_write(Tile_X01_Y02_config_out_write),
    .flush(Tile_X01_Y02_flush_out),
    .flush_out(Tile_X01_Y03_flush_out),
    .hi(Tile_X01_Y03_hi),
    .lo(Tile_X01_Y03_lo),
    .read_config_data(Tile_X01_Y03_read_config_data),
    .read_config_data_in(Tile_X01_Y02_read_config_data),
    .reset(Tile_X01_Y02_reset_out),
    .reset_out(Tile_X01_Y03_reset_out),
    .stall(Tile_X01_Y02_stall_out),
    .stall_out(Tile_X01_Y03_stall_out),
    .tile_id(Tile_X01_Y03_tile_id)
);
wire [15:0] Tile_X01_Y04_tile_id;
assign Tile_X01_Y04_tile_id = {Tile_X01_Y04_lo[7],Tile_X01_Y04_lo[7],Tile_X01_Y04_lo[6],Tile_X01_Y04_lo[6],Tile_X01_Y04_lo[5],Tile_X01_Y04_lo[5],Tile_X01_Y04_lo[4],Tile_X01_Y04_hi[4],Tile_X01_Y04_lo[3],Tile_X01_Y04_lo[3],Tile_X01_Y04_lo[2],Tile_X01_Y04_lo[2],Tile_X01_Y04_lo[1],Tile_X01_Y04_hi[1],Tile_X01_Y04_lo[0],Tile_X01_Y04_lo[0]};
Tile_PE Tile_X01_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y03_clk_out),
    .clk_out(Tile_X01_Y04_clk_out),
    .clk_pass_through(Tile_X01_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y04_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y03_config_out_config_addr),
    .config_config_data(Tile_X01_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y04_config_out_config_data),
    .config_out_read(Tile_X01_Y04_config_out_read),
    .config_out_write(Tile_X01_Y04_config_out_write),
    .config_read(Tile_X01_Y03_config_out_read),
    .config_write(Tile_X01_Y03_config_out_write),
    .flush(Tile_X01_Y03_flush_out),
    .flush_out(Tile_X01_Y04_flush_out),
    .hi(Tile_X01_Y04_hi),
    .lo(Tile_X01_Y04_lo),
    .read_config_data(Tile_X01_Y04_read_config_data),
    .read_config_data_in(Tile_X01_Y03_read_config_data),
    .reset(Tile_X01_Y03_reset_out),
    .reset_out(Tile_X01_Y04_reset_out),
    .stall(Tile_X01_Y03_stall_out),
    .stall_out(Tile_X01_Y04_stall_out),
    .tile_id(Tile_X01_Y04_tile_id)
);
wire [15:0] Tile_X02_Y00_tile_id;
assign Tile_X02_Y00_tile_id = {Tile_X02_Y00_lo[7],Tile_X02_Y00_lo[7],Tile_X02_Y00_lo[6],Tile_X02_Y00_lo[6],Tile_X02_Y00_lo[5],Tile_X02_Y00_lo[5],Tile_X02_Y00_hi[5],Tile_X02_Y00_lo[4],Tile_X02_Y00_lo[3],Tile_X02_Y00_lo[3],Tile_X02_Y00_lo[2],Tile_X02_Y00_lo[2],Tile_X02_Y00_lo[1],Tile_X02_Y00_lo[1],Tile_X02_Y00_lo[0],Tile_X02_Y00_lo[0]};
Tile_io_core Tile_X02_Y00 (
    .tile_id(Tile_X02_Y00_tile_id),
    .glb2io_1(glb2io_1_X02_Y00),
    .f2io_1(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X02_Y00_io2glb_1),
    .io2f_1(Tile_X02_Y00_io2f_1),
    .glb2io_16(glb2io_16_X02_Y00),
    .f2io_16(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X02_Y00_io2glb_16),
    .io2f_16(Tile_X02_Y00_io2f_16),
    .hi(Tile_X02_Y00_hi),
    .lo(Tile_X02_Y00_lo)
);
wire [15:0] Tile_X02_Y01_tile_id;
assign Tile_X02_Y01_tile_id = {Tile_X02_Y01_lo[7],Tile_X02_Y01_lo[7],Tile_X02_Y01_lo[6],Tile_X02_Y01_lo[6],Tile_X02_Y01_lo[5],Tile_X02_Y01_lo[5],Tile_X02_Y01_hi[5],Tile_X02_Y01_lo[4],Tile_X02_Y01_lo[3],Tile_X02_Y01_lo[3],Tile_X02_Y01_lo[2],Tile_X02_Y01_lo[2],Tile_X02_Y01_lo[1],Tile_X02_Y01_lo[1],Tile_X02_Y01_lo[0],Tile_X02_Y01_hi[0]};
Tile_PE Tile_X02_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .clk_out(Tile_X02_Y01_clk_out),
    .clk_pass_through(coreir_wrapInClock_inst2_out),
    .clk_pass_through_out_bot(Tile_X02_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y01_clk_pass_through_out_right),
    .config_config_addr(config_2_config_addr),
    .config_config_data(config_2_config_data),
    .config_out_config_addr(Tile_X02_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y01_config_out_config_data),
    .config_out_read(Tile_X02_Y01_config_out_read),
    .config_out_write(Tile_X02_Y01_config_out_write),
    .config_read(config_2_read),
    .config_write(config_2_write),
    .flush(flush),
    .flush_out(Tile_X02_Y01_flush_out),
    .hi(Tile_X02_Y01_hi),
    .lo(Tile_X02_Y01_lo),
    .read_config_data(Tile_X02_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X02_Y01_reset_out),
    .stall(self_stall_out[2:2]),
    .stall_out(Tile_X02_Y01_stall_out),
    .tile_id(Tile_X02_Y01_tile_id)
);
wire [15:0] Tile_X02_Y02_tile_id;
assign Tile_X02_Y02_tile_id = {Tile_X02_Y02_lo[7],Tile_X02_Y02_lo[7],Tile_X02_Y02_lo[6],Tile_X02_Y02_lo[6],Tile_X02_Y02_lo[5],Tile_X02_Y02_lo[5],Tile_X02_Y02_hi[5],Tile_X02_Y02_lo[4],Tile_X02_Y02_lo[3],Tile_X02_Y02_lo[3],Tile_X02_Y02_lo[2],Tile_X02_Y02_lo[2],Tile_X02_Y02_lo[1],Tile_X02_Y02_lo[1],Tile_X02_Y02_hi[1],Tile_X02_Y02_lo[0]};
Tile_PE Tile_X02_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y01_clk_out),
    .clk_out(Tile_X02_Y02_clk_out),
    .clk_pass_through(Tile_X02_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y02_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y01_config_out_config_addr),
    .config_config_data(Tile_X02_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y02_config_out_config_data),
    .config_out_read(Tile_X02_Y02_config_out_read),
    .config_out_write(Tile_X02_Y02_config_out_write),
    .config_read(Tile_X02_Y01_config_out_read),
    .config_write(Tile_X02_Y01_config_out_write),
    .flush(Tile_X02_Y01_flush_out),
    .flush_out(Tile_X02_Y02_flush_out),
    .hi(Tile_X02_Y02_hi),
    .lo(Tile_X02_Y02_lo),
    .read_config_data(Tile_X02_Y02_read_config_data),
    .read_config_data_in(Tile_X02_Y01_read_config_data),
    .reset(Tile_X02_Y01_reset_out),
    .reset_out(Tile_X02_Y02_reset_out),
    .stall(Tile_X02_Y01_stall_out),
    .stall_out(Tile_X02_Y02_stall_out),
    .tile_id(Tile_X02_Y02_tile_id)
);
wire [15:0] Tile_X02_Y03_tile_id;
assign Tile_X02_Y03_tile_id = {Tile_X02_Y03_lo[7],Tile_X02_Y03_lo[7],Tile_X02_Y03_lo[6],Tile_X02_Y03_lo[6],Tile_X02_Y03_lo[5],Tile_X02_Y03_lo[5],Tile_X02_Y03_hi[5],Tile_X02_Y03_lo[4],Tile_X02_Y03_lo[3],Tile_X02_Y03_lo[3],Tile_X02_Y03_lo[2],Tile_X02_Y03_lo[2],Tile_X02_Y03_lo[1],Tile_X02_Y03_lo[1],Tile_X02_Y03_hi[1],Tile_X02_Y03_hi[0]};
Tile_PE Tile_X02_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y02_clk_out),
    .clk_out(Tile_X02_Y03_clk_out),
    .clk_pass_through(Tile_X02_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y03_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y02_config_out_config_addr),
    .config_config_data(Tile_X02_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y03_config_out_config_data),
    .config_out_read(Tile_X02_Y03_config_out_read),
    .config_out_write(Tile_X02_Y03_config_out_write),
    .config_read(Tile_X02_Y02_config_out_read),
    .config_write(Tile_X02_Y02_config_out_write),
    .flush(Tile_X02_Y02_flush_out),
    .flush_out(Tile_X02_Y03_flush_out),
    .hi(Tile_X02_Y03_hi),
    .lo(Tile_X02_Y03_lo),
    .read_config_data(Tile_X02_Y03_read_config_data),
    .read_config_data_in(Tile_X02_Y02_read_config_data),
    .reset(Tile_X02_Y02_reset_out),
    .reset_out(Tile_X02_Y03_reset_out),
    .stall(Tile_X02_Y02_stall_out),
    .stall_out(Tile_X02_Y03_stall_out),
    .tile_id(Tile_X02_Y03_tile_id)
);
wire [15:0] Tile_X02_Y04_tile_id;
assign Tile_X02_Y04_tile_id = {Tile_X02_Y04_lo[7],Tile_X02_Y04_lo[7],Tile_X02_Y04_lo[6],Tile_X02_Y04_lo[6],Tile_X02_Y04_lo[5],Tile_X02_Y04_lo[5],Tile_X02_Y04_hi[5],Tile_X02_Y04_lo[4],Tile_X02_Y04_lo[3],Tile_X02_Y04_lo[3],Tile_X02_Y04_lo[2],Tile_X02_Y04_lo[2],Tile_X02_Y04_lo[1],Tile_X02_Y04_hi[1],Tile_X02_Y04_lo[0],Tile_X02_Y04_lo[0]};
Tile_PE Tile_X02_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y03_clk_out),
    .clk_out(Tile_X02_Y04_clk_out),
    .clk_pass_through(Tile_X02_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y04_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y03_config_out_config_addr),
    .config_config_data(Tile_X02_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y04_config_out_config_data),
    .config_out_read(Tile_X02_Y04_config_out_read),
    .config_out_write(Tile_X02_Y04_config_out_write),
    .config_read(Tile_X02_Y03_config_out_read),
    .config_write(Tile_X02_Y03_config_out_write),
    .flush(Tile_X02_Y03_flush_out),
    .flush_out(Tile_X02_Y04_flush_out),
    .hi(Tile_X02_Y04_hi),
    .lo(Tile_X02_Y04_lo),
    .read_config_data(Tile_X02_Y04_read_config_data),
    .read_config_data_in(Tile_X02_Y03_read_config_data),
    .reset(Tile_X02_Y03_reset_out),
    .reset_out(Tile_X02_Y04_reset_out),
    .stall(Tile_X02_Y03_stall_out),
    .stall_out(Tile_X02_Y04_stall_out),
    .tile_id(Tile_X02_Y04_tile_id)
);
wire [15:0] Tile_X03_Y00_tile_id;
assign Tile_X03_Y00_tile_id = {Tile_X03_Y00_lo[7],Tile_X03_Y00_lo[7],Tile_X03_Y00_lo[6],Tile_X03_Y00_lo[6],Tile_X03_Y00_lo[5],Tile_X03_Y00_lo[5],Tile_X03_Y00_hi[5],Tile_X03_Y00_hi[4],Tile_X03_Y00_lo[3],Tile_X03_Y00_lo[3],Tile_X03_Y00_lo[2],Tile_X03_Y00_lo[2],Tile_X03_Y00_lo[1],Tile_X03_Y00_lo[1],Tile_X03_Y00_lo[0],Tile_X03_Y00_lo[0]};
Tile_io_core Tile_X03_Y00 (
    .tile_id(Tile_X03_Y00_tile_id),
    .glb2io_1(glb2io_1_X03_Y00),
    .f2io_1(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X03_Y00_io2glb_1),
    .io2f_1(Tile_X03_Y00_io2f_1),
    .glb2io_16(glb2io_16_X03_Y00),
    .f2io_16(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X03_Y00_io2glb_16),
    .io2f_16(Tile_X03_Y00_io2f_16),
    .hi(Tile_X03_Y00_hi),
    .lo(Tile_X03_Y00_lo)
);
wire [15:0] Tile_X03_Y01_tile_id;
assign Tile_X03_Y01_tile_id = {Tile_X03_Y01_lo[7],Tile_X03_Y01_lo[7],Tile_X03_Y01_lo[6],Tile_X03_Y01_lo[6],Tile_X03_Y01_lo[5],Tile_X03_Y01_lo[5],Tile_X03_Y01_hi[5],Tile_X03_Y01_hi[4],Tile_X03_Y01_lo[3],Tile_X03_Y01_lo[3],Tile_X03_Y01_lo[2],Tile_X03_Y01_lo[2],Tile_X03_Y01_lo[1],Tile_X03_Y01_lo[1],Tile_X03_Y01_lo[0],Tile_X03_Y01_hi[0]};
Tile_MemCore Tile_X03_Y01 (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y01_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y01_clk_out),
    .config_config_addr(config_3_config_addr),
    .config_config_data(config_3_config_data),
    .config_out_config_addr(Tile_X03_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y01_config_out_config_data),
    .config_out_read(Tile_X03_Y01_config_out_read),
    .config_out_write(Tile_X03_Y01_config_out_write),
    .config_read(config_3_read),
    .config_write(config_3_write),
    .flush(flush),
    .flush_out(Tile_X03_Y01_flush_out),
    .hi(Tile_X03_Y01_hi),
    .lo(Tile_X03_Y01_lo),
    .read_config_data(Tile_X03_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X03_Y01_reset_out),
    .stall(self_stall_out[3:3]),
    .stall_out(Tile_X03_Y01_stall_out),
    .tile_id(Tile_X03_Y01_tile_id)
);
wire [15:0] Tile_X03_Y02_tile_id;
assign Tile_X03_Y02_tile_id = {Tile_X03_Y02_lo[7],Tile_X03_Y02_lo[7],Tile_X03_Y02_lo[6],Tile_X03_Y02_lo[6],Tile_X03_Y02_lo[5],Tile_X03_Y02_lo[5],Tile_X03_Y02_hi[5],Tile_X03_Y02_hi[4],Tile_X03_Y02_lo[3],Tile_X03_Y02_lo[3],Tile_X03_Y02_lo[2],Tile_X03_Y02_lo[2],Tile_X03_Y02_lo[1],Tile_X03_Y02_lo[1],Tile_X03_Y02_hi[1],Tile_X03_Y02_lo[0]};
Tile_MemCore Tile_X03_Y02 (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y02_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y02_clk_out),
    .config_config_addr(Tile_X03_Y01_config_out_config_addr),
    .config_config_data(Tile_X03_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y02_config_out_config_data),
    .config_out_read(Tile_X03_Y02_config_out_read),
    .config_out_write(Tile_X03_Y02_config_out_write),
    .config_read(Tile_X03_Y01_config_out_read),
    .config_write(Tile_X03_Y01_config_out_write),
    .flush(Tile_X03_Y01_flush_out),
    .flush_out(Tile_X03_Y02_flush_out),
    .hi(Tile_X03_Y02_hi),
    .lo(Tile_X03_Y02_lo),
    .read_config_data(Tile_X03_Y02_read_config_data),
    .read_config_data_in(Tile_X03_Y01_read_config_data),
    .reset(Tile_X03_Y01_reset_out),
    .reset_out(Tile_X03_Y02_reset_out),
    .stall(Tile_X03_Y01_stall_out),
    .stall_out(Tile_X03_Y02_stall_out),
    .tile_id(Tile_X03_Y02_tile_id)
);
wire [15:0] Tile_X03_Y03_tile_id;
assign Tile_X03_Y03_tile_id = {Tile_X03_Y03_lo[7],Tile_X03_Y03_lo[7],Tile_X03_Y03_lo[6],Tile_X03_Y03_lo[6],Tile_X03_Y03_lo[5],Tile_X03_Y03_lo[5],Tile_X03_Y03_hi[5],Tile_X03_Y03_hi[4],Tile_X03_Y03_lo[3],Tile_X03_Y03_lo[3],Tile_X03_Y03_lo[2],Tile_X03_Y03_lo[2],Tile_X03_Y03_lo[1],Tile_X03_Y03_lo[1],Tile_X03_Y03_hi[1],Tile_X03_Y03_hi[0]};
Tile_MemCore Tile_X03_Y03 (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y03_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y03_clk_out),
    .config_config_addr(Tile_X03_Y02_config_out_config_addr),
    .config_config_data(Tile_X03_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y03_config_out_config_data),
    .config_out_read(Tile_X03_Y03_config_out_read),
    .config_out_write(Tile_X03_Y03_config_out_write),
    .config_read(Tile_X03_Y02_config_out_read),
    .config_write(Tile_X03_Y02_config_out_write),
    .flush(Tile_X03_Y02_flush_out),
    .flush_out(Tile_X03_Y03_flush_out),
    .hi(Tile_X03_Y03_hi),
    .lo(Tile_X03_Y03_lo),
    .read_config_data(Tile_X03_Y03_read_config_data),
    .read_config_data_in(Tile_X03_Y02_read_config_data),
    .reset(Tile_X03_Y02_reset_out),
    .reset_out(Tile_X03_Y03_reset_out),
    .stall(Tile_X03_Y02_stall_out),
    .stall_out(Tile_X03_Y03_stall_out),
    .tile_id(Tile_X03_Y03_tile_id)
);
wire [15:0] Tile_X03_Y04_tile_id;
assign Tile_X03_Y04_tile_id = {Tile_X03_Y04_lo[7],Tile_X03_Y04_lo[7],Tile_X03_Y04_lo[6],Tile_X03_Y04_lo[6],Tile_X03_Y04_lo[5],Tile_X03_Y04_lo[5],Tile_X03_Y04_hi[5],Tile_X03_Y04_hi[4],Tile_X03_Y04_lo[3],Tile_X03_Y04_lo[3],Tile_X03_Y04_lo[2],Tile_X03_Y04_lo[2],Tile_X03_Y04_lo[1],Tile_X03_Y04_hi[1],Tile_X03_Y04_lo[0],Tile_X03_Y04_lo[0]};
Tile_MemCore Tile_X03_Y04 (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y04_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y04_clk_out),
    .config_config_addr(Tile_X03_Y03_config_out_config_addr),
    .config_config_data(Tile_X03_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y04_config_out_config_data),
    .config_out_read(Tile_X03_Y04_config_out_read),
    .config_out_write(Tile_X03_Y04_config_out_write),
    .config_read(Tile_X03_Y03_config_out_read),
    .config_write(Tile_X03_Y03_config_out_write),
    .flush(Tile_X03_Y03_flush_out),
    .flush_out(Tile_X03_Y04_flush_out),
    .hi(Tile_X03_Y04_hi),
    .lo(Tile_X03_Y04_lo),
    .read_config_data(Tile_X03_Y04_read_config_data),
    .read_config_data_in(Tile_X03_Y03_read_config_data),
    .reset(Tile_X03_Y03_reset_out),
    .reset_out(Tile_X03_Y04_reset_out),
    .stall(Tile_X03_Y03_stall_out),
    .stall_out(Tile_X03_Y04_stall_out),
    .tile_id(Tile_X03_Y04_tile_id)
);
coreir_const #(
    .value(1'h0),
    .width(1)
) const_0_1 (
    .out(const_0_1_out)
);
coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
coreir_const #(
    .value(32'h00000000),
    .width(32)
) const_0_32 (
    .out(const_0_32_out)
);
coreir_wrap coreir_wrapInClock_inst0 (
    .in(clk),
    .out(coreir_wrapInClock_inst0_out)
);
coreir_wrap coreir_wrapInClock_inst1 (
    .in(clk),
    .out(coreir_wrapInClock_inst1_out)
);
coreir_wrap coreir_wrapInClock_inst2 (
    .in(clk),
    .out(coreir_wrapInClock_inst2_out)
);
Or4x32 read_config_data_or_final (
    .I0(Tile_X00_Y04_read_config_data),
    .I1(Tile_X01_Y04_read_config_data),
    .I2(Tile_X02_Y04_read_config_data),
    .I3(Tile_X03_Y04_read_config_data),
    .O(read_config_data_or_final_O)
);
mantle_wire__typeBit4 self_stall (
    .in(stall),
    .out(self_stall_out)
);
assign io2glb_16_X00_Y00 = Tile_X00_Y00_io2glb_16;
assign io2glb_16_X01_Y00 = Tile_X01_Y00_io2glb_16;
assign io2glb_16_X02_Y00 = Tile_X02_Y00_io2glb_16;
assign io2glb_16_X03_Y00 = Tile_X03_Y00_io2glb_16;
assign io2glb_1_X00_Y00 = Tile_X00_Y00_io2glb_1;
assign io2glb_1_X01_Y00 = Tile_X01_Y00_io2glb_1;
assign io2glb_1_X02_Y00 = Tile_X02_Y00_io2glb_1;
assign io2glb_1_X03_Y00 = Tile_X03_Y00_io2glb_1;
assign read_config_data = read_config_data_or_final_O;
endmodule

module Garnet (
    input [12:0] axi4_slave_araddr,
    output axi4_slave_arready,
    input axi4_slave_arvalid,
    input [12:0] axi4_slave_awaddr,
    output axi4_slave_awready,
    input axi4_slave_awvalid,
    input axi4_slave_bready,
    output [1:0] axi4_slave_bresp,
    output axi4_slave_bvalid,
    output [31:0] axi4_slave_rdata,
    input axi4_slave_rready,
    output [1:0] axi4_slave_rresp,
    output axi4_slave_rvalid,
    input [31:0] axi4_slave_wdata,
    output axi4_slave_wready,
    input axi4_slave_wvalid,
    output cgra_running_clk_out,
    input clk_in,
    output interrupt,
    input jtag_tck,
    input jtag_tdi,
    output jtag_tdo,
    input jtag_tms,
    input jtag_trst_n,
    input [18:0] proc_packet_rd_addr,
    output [63:0] proc_packet_rd_data,
    output proc_packet_rd_data_valid,
    input proc_packet_rd_en,
    input [18:0] proc_packet_wr_addr,
    input [63:0] proc_packet_wr_data,
    input proc_packet_wr_en,
    input [7:0] proc_packet_wr_strb,
    input reset_in
);
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_clk_out;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_reset_out;
wire [3:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_stall;
wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_clk_en_master;
wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_clk_en_bank_master;
wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_pcfg_broadcast_stall;
wire [0:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_flush_crossbar_sel;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_en;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_clk_en;
wire [11:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_addr;
wire [31:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_data;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_en;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_clk_en;
wire [11:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_addr;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_en;
wire [18:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_addr;
wire [31:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_data;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_rd_en;
wire [18:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_rd_addr;
wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_strm_g2f_start_pulse;
wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_strm_f2g_start_pulse;
wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_pc_start_pulse;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_read;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_write;
wire [31:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_addr;
wire [31:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_wr_data;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_awready;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_wready;
wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_bresp;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_bvalid;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_arready;
wire [31:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rdata;
wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rresp;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rvalid;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_interrupt;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_tdo;
wire [15:0] Interconnect_inst0_io2glb_16_X00_Y00;
wire [15:0] Interconnect_inst0_io2glb_16_X01_Y00;
wire [15:0] Interconnect_inst0_io2glb_16_X02_Y00;
wire [15:0] Interconnect_inst0_io2glb_16_X03_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X00_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X01_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X02_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X03_Y00;
wire [31:0] Interconnect_inst0_read_config_data;
wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_1_1;
wire [1:0] global_buffer_W_inst0_strm_f2g_interrupt_pulse;
wire [0:0] global_buffer_W_inst0_if_sram_cfg_rd_data_valid;
wire [0:0] global_buffer_W_inst0_strm_data_valid_g2f_1_1;
wire [0:0] global_buffer_W_inst0_strm_data_valid_g2f_0_0;
wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_0_0;
wire [0:0] global_buffer_W_inst0_strm_data_valid_g2f_0_1;
wire [15:0] global_buffer_W_inst0_strm_data_g2f_0_0;
wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_1_1;
wire [63:0] global_buffer_W_inst0_proc_rd_data;
wire [1:0] global_buffer_W_inst0_pcfg_g2f_interrupt_pulse;
wire [31:0] global_buffer_W_inst0_if_cfg_rd_data;
wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_1_1;
wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_0_1;
wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_1_1;
wire [0:0] global_buffer_W_inst0_strm_data_flush_g2f;
wire [15:0] global_buffer_W_inst0_strm_data_g2f_1_1;
wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_1_0;
wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_1_0;
wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_0_0;
wire [15:0] global_buffer_W_inst0_strm_data_g2f_0_1;
wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_0_1;
wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_0_1;
wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_1_0;
wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_0_1;
wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_1_0;
wire [0:0] global_buffer_W_inst0_strm_data_valid_g2f_1_0;
wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_0_0;
wire [15:0] global_buffer_W_inst0_strm_data_g2f_1_0;
wire [31:0] global_buffer_W_inst0_if_sram_cfg_rd_data;
wire [0:0] global_buffer_W_inst0_proc_rd_data_valid;
wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_0_0;
wire [0:0] global_buffer_W_inst0_if_cfg_rd_data_valid;
wire [1:0] global_buffer_W_inst0_strm_g2f_interrupt_pulse;
wire [3:0] global_buffer_W_inst0_cgra_stall;
global_controller GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0 (
    .clk_in(clk_in),
    .reset_in(reset_in),
    .clk_out(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_clk_out),
    .reset_out(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_reset_out),
    .cgra_stall(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_stall),
    .glb_clk_en_master(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_clk_en_master),
    .glb_clk_en_bank_master(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_clk_en_bank_master),
    .glb_pcfg_broadcast_stall(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_pcfg_broadcast_stall),
    .glb_flush_crossbar_sel(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_flush_crossbar_sel),
    .glb_cfg_wr_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_en),
    .glb_cfg_wr_clk_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_clk_en),
    .glb_cfg_wr_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_addr),
    .glb_cfg_wr_data(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_data),
    .glb_cfg_rd_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_en),
    .glb_cfg_rd_clk_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_clk_en),
    .glb_cfg_rd_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_addr),
    .glb_cfg_rd_data(global_buffer_W_inst0_if_cfg_rd_data),
    .glb_cfg_rd_data_valid(global_buffer_W_inst0_if_cfg_rd_data_valid[0]),
    .sram_cfg_wr_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_en),
    .sram_cfg_wr_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_addr),
    .sram_cfg_wr_data(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_data),
    .sram_cfg_rd_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_rd_en),
    .sram_cfg_rd_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_rd_addr),
    .sram_cfg_rd_data(global_buffer_W_inst0_if_sram_cfg_rd_data),
    .sram_cfg_rd_data_valid(global_buffer_W_inst0_if_sram_cfg_rd_data_valid[0]),
    .strm_g2f_start_pulse(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_strm_g2f_start_pulse),
    .strm_f2g_start_pulse(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_strm_f2g_start_pulse),
    .pc_start_pulse(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_pc_start_pulse),
    .strm_g2f_interrupt_pulse(global_buffer_W_inst0_strm_g2f_interrupt_pulse),
    .strm_f2g_interrupt_pulse(global_buffer_W_inst0_strm_f2g_interrupt_pulse),
    .pcfg_g2f_interrupt_pulse(global_buffer_W_inst0_pcfg_g2f_interrupt_pulse),
    .cgra_cfg_read(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_read),
    .cgra_cfg_write(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_write),
    .cgra_cfg_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_addr),
    .cgra_cfg_wr_data(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_wr_data),
    .cgra_cfg_rd_data(Interconnect_inst0_read_config_data),
    .axi_awaddr(axi4_slave_awaddr),
    .axi_awvalid(axi4_slave_awvalid),
    .axi_awready(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_awready),
    .axi_wdata(axi4_slave_wdata),
    .axi_wvalid(axi4_slave_wvalid),
    .axi_wready(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_wready),
    .axi_bready(axi4_slave_bready),
    .axi_bresp(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_bresp),
    .axi_bvalid(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_bvalid),
    .axi_araddr(axi4_slave_araddr),
    .axi_arvalid(axi4_slave_arvalid),
    .axi_arready(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_arready),
    .axi_rdata(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rdata),
    .axi_rresp(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rresp),
    .axi_rvalid(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rvalid),
    .axi_rready(axi4_slave_rready),
    .interrupt(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_interrupt),
    .tck(jtag_tck),
    .tdi(jtag_tdi),
    .tms(jtag_tms),
    .trst_n(jtag_trst_n),
    .tdo(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_tdo)
);
Interconnect Interconnect_inst0 (
    .clk(clk_in),
    .config_0_config_addr(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_0_0),
    .config_0_config_data(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_0_0),
    .config_0_read(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_0_0),
    .config_0_write(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_0_0),
    .config_1_config_addr(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_0_1),
    .config_1_config_data(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_0_1),
    .config_1_read(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_0_1),
    .config_1_write(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_0_1),
    .config_2_config_addr(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_1_0),
    .config_2_config_data(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_1_0),
    .config_2_read(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_1_0),
    .config_2_write(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_1_0),
    .config_3_config_addr(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_1_1),
    .config_3_config_data(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_1_1),
    .config_3_read(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_1_1),
    .config_3_write(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_1_1),
    .flush(global_buffer_W_inst0_strm_data_flush_g2f),
    .glb2io_16_X00_Y00(global_buffer_W_inst0_strm_data_g2f_0_0),
    .glb2io_16_X01_Y00(global_buffer_W_inst0_strm_data_g2f_0_1),
    .glb2io_16_X02_Y00(global_buffer_W_inst0_strm_data_g2f_1_0),
    .glb2io_16_X03_Y00(global_buffer_W_inst0_strm_data_g2f_1_1),
    .glb2io_1_X00_Y00(global_buffer_W_inst0_strm_data_valid_g2f_0_0),
    .glb2io_1_X01_Y00(global_buffer_W_inst0_strm_data_valid_g2f_0_1),
    .glb2io_1_X02_Y00(global_buffer_W_inst0_strm_data_valid_g2f_1_0),
    .glb2io_1_X03_Y00(global_buffer_W_inst0_strm_data_valid_g2f_1_1),
    .io2glb_16_X00_Y00(Interconnect_inst0_io2glb_16_X00_Y00),
    .io2glb_16_X01_Y00(Interconnect_inst0_io2glb_16_X01_Y00),
    .io2glb_16_X02_Y00(Interconnect_inst0_io2glb_16_X02_Y00),
    .io2glb_16_X03_Y00(Interconnect_inst0_io2glb_16_X03_Y00),
    .io2glb_1_X00_Y00(Interconnect_inst0_io2glb_1_X00_Y00),
    .io2glb_1_X01_Y00(Interconnect_inst0_io2glb_1_X01_Y00),
    .io2glb_1_X02_Y00(Interconnect_inst0_io2glb_1_X02_Y00),
    .io2glb_1_X03_Y00(Interconnect_inst0_io2glb_1_X03_Y00),
    .read_config_data(Interconnect_inst0_read_config_data),
    .reset(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_reset_out),
    .stall(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_stall)
);
global_buffer_W global_buffer_W_inst0 (
    .cgra_cfg_g2f_cfg_addr_1_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_1_1),
    .if_cfg_rd_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_en),
    .strm_f2g_interrupt_pulse(global_buffer_W_inst0_strm_f2g_interrupt_pulse),
    .proc_wr_addr(proc_packet_wr_addr),
    .if_cfg_rd_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_addr),
    .if_sram_cfg_rd_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_rd_addr),
    .if_sram_cfg_rd_data_valid(global_buffer_W_inst0_if_sram_cfg_rd_data_valid),
    .proc_rd_en(proc_packet_rd_en),
    .strm_data_valid_f2g_1_0(Interconnect_inst0_io2glb_1_X02_Y00),
    .if_sram_cfg_wr_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_addr),
    .pcfg_start_pulse(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_pc_start_pulse),
    .strm_data_valid_g2f_1_1(global_buffer_W_inst0_strm_data_valid_g2f_1_1),
    .clk(clk_in),
    .strm_data_valid_f2g_0_0(Interconnect_inst0_io2glb_1_X00_Y00),
    .strm_data_valid_g2f_0_0(global_buffer_W_inst0_strm_data_valid_g2f_0_0),
    .cgra_cfg_jtag_gc2glb_rd_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_read),
    .if_cfg_wr_clk_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_clk_en),
    .cgra_cfg_g2f_cfg_wr_en_0_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_0_0),
    .proc_rd_addr(proc_packet_rd_addr),
    .strm_data_f2g_1_0(Interconnect_inst0_io2glb_16_X02_Y00),
    .strm_data_valid_g2f_0_1(global_buffer_W_inst0_strm_data_valid_g2f_0_1),
    .if_cfg_wr_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_addr),
    .strm_data_g2f_0_0(global_buffer_W_inst0_strm_data_g2f_0_0),
    .proc_wr_en(proc_packet_wr_en),
    .pcfg_broadcast_stall(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_pcfg_broadcast_stall),
    .if_cfg_rd_clk_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_clk_en),
    .cgra_cfg_g2f_cfg_rd_en_1_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_1_1),
    .cgra_stall_in(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_stall),
    .proc_rd_data(global_buffer_W_inst0_proc_rd_data),
    .strm_data_valid_f2g_1_1(Interconnect_inst0_io2glb_1_X03_Y00),
    .pcfg_g2f_interrupt_pulse(global_buffer_W_inst0_pcfg_g2f_interrupt_pulse),
    .if_cfg_rd_data(global_buffer_W_inst0_if_cfg_rd_data),
    .reset(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_reset_out),
    .if_sram_cfg_wr_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_en),
    .cgra_cfg_jtag_gc2glb_wr_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_write),
    .if_sram_cfg_wr_data(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_data),
    .cgra_cfg_g2f_cfg_data_1_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_1_1),
    .cgra_cfg_g2f_cfg_rd_en_0_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_0_1),
    .cgra_cfg_g2f_cfg_wr_en_1_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_1_1),
    .strm_data_flush_g2f(global_buffer_W_inst0_strm_data_flush_g2f),
    .strm_data_f2g_0_0(Interconnect_inst0_io2glb_16_X00_Y00),
    .strm_data_g2f_1_1(global_buffer_W_inst0_strm_data_g2f_1_1),
    .strm_f2g_start_pulse(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_strm_f2g_start_pulse),
    .glb_clk_en_master(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_clk_en_master),
    .strm_data_f2g_0_1(Interconnect_inst0_io2glb_16_X01_Y00),
    .if_sram_cfg_rd_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_rd_en),
    .if_cfg_wr_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_en),
    .cgra_cfg_g2f_cfg_data_1_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_1_0),
    .cgra_cfg_g2f_cfg_addr_1_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_1_0),
    .cgra_cfg_g2f_cfg_rd_en_0_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_0_0),
    .strm_data_f2g_1_1(Interconnect_inst0_io2glb_16_X03_Y00),
    .strm_data_g2f_0_1(global_buffer_W_inst0_strm_data_g2f_0_1),
    .cgra_cfg_g2f_cfg_addr_0_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_0_1),
    .cgra_cfg_g2f_cfg_wr_en_0_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_0_1),
    .cgra_cfg_g2f_cfg_rd_en_1_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_1_0),
    .cgra_cfg_g2f_cfg_data_0_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_0_1),
    .cgra_cfg_g2f_cfg_wr_en_1_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_1_0),
    .cgra_cfg_jtag_gc2glb_data(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_wr_data),
    .strm_data_valid_g2f_1_0(global_buffer_W_inst0_strm_data_valid_g2f_1_0),
    .cgra_cfg_g2f_cfg_addr_0_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_0_0),
    .strm_data_g2f_1_0(global_buffer_W_inst0_strm_data_g2f_1_0),
    .if_cfg_wr_data(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_data),
    .strm_data_valid_f2g_0_1(Interconnect_inst0_io2glb_1_X01_Y00),
    .strm_g2f_start_pulse(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_strm_g2f_start_pulse),
    .flush_crossbar_sel(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_flush_crossbar_sel),
    .proc_wr_data(proc_packet_wr_data),
    .if_sram_cfg_rd_data(global_buffer_W_inst0_if_sram_cfg_rd_data),
    .proc_rd_data_valid(global_buffer_W_inst0_proc_rd_data_valid),
    .cgra_cfg_g2f_cfg_data_0_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_0_0),
    .glb_clk_en_bank_master(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_clk_en_bank_master),
    .if_cfg_rd_data_valid(global_buffer_W_inst0_if_cfg_rd_data_valid),
    .proc_wr_strb(proc_packet_wr_strb),
    .strm_g2f_interrupt_pulse(global_buffer_W_inst0_strm_g2f_interrupt_pulse),
    .cgra_cfg_jtag_gc2glb_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_addr),
    .cgra_stall(global_buffer_W_inst0_cgra_stall)
);
assign axi4_slave_arready = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_arready;
assign axi4_slave_awready = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_awready;
assign axi4_slave_bresp = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_bresp;
assign axi4_slave_bvalid = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_bvalid;
assign axi4_slave_rdata = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rdata;
assign axi4_slave_rresp = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rresp;
assign axi4_slave_rvalid = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rvalid;
assign axi4_slave_wready = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_wready;
assign cgra_running_clk_out = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_clk_out;
assign interrupt = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_interrupt;
assign jtag_tdo = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_tdo;
assign proc_packet_rd_data = global_buffer_W_inst0_proc_rd_data;
assign proc_packet_rd_data_valid = global_buffer_W_inst0_proc_rd_data_valid[0];
endmodule

