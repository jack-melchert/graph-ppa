// Module `global_controller` defined externally
module mux_aoi_ready_valid_const_21_17 ( 
	input logic  [16 : 0] I[20:0], 
	input logic  [4 : 0] S ,
	input logic ready_in,
	output logic ready_out,
	input logic [20:0]  valid_in,
	output logic valid_out,
	output logic  [31 : 0] out_sel,
	output logic [16 : 0] O); 
	logic  [16 : 0] O_int0;
	logic  [16 : 0] O_int1;
	logic  [16 : 0] O_int2;
	logic  [16 : 0] O_int3;
	logic  [16 : 0] O_int4;
	logic  [16 : 0] O_int5;
	logic  [16 : 0] O_int6;
	logic  [16 : 0] O_int7;
	logic  [16 : 0] O_int8;
	logic  [16 : 0] O_int9;
	logic  [16 : 0] O_int10;
	logic [10:0] valid_out_temp;

precoder_17_21 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_17_21 u_mux_logic ( 
	.I0 (I[0]),
	.I1 (I[1]),
	.I2 (I[2]),
	.I3 (I[3]),
	.I4 (I[4]),
	.I5 (I[5]),
	.I6 (I[6]),
	.I7 (I[7]),
	.I8 (I[8]),
	.I9 (I[9]),
	.I10 (I[10]),
	.I11 (I[11]),
	.I12 (I[12]),
	.I13 (I[13]),
	.I14 (I[14]),
	.I15 (I[15]),
	.I16 (I[16]),
	.I17 (I[17]),
	.I18 (I[18]),
	.I19 (I[19]),
	.I20 (I[20]),
	.out_sel(out_sel), 
	.valid_in(valid_in),
	.valid_out(valid_out_temp),
	.O0(O_int0), 
	.O1(O_int1), 
	.O2(O_int2), 
	.O3(O_int3), 
	.O4(O_int4), 
	.O5(O_int5), 
	.O6(O_int6), 
	.O7(O_int7), 
	.O8(O_int8), 
	.O9(O_int9), 
	.O10(O_int10)); 
	assign O = (  	O_int0 | 	O_int1 | 	O_int2 | 	O_int3 | 	O_int4 | 	O_int5 | 	O_int6 | 	O_int7 | 	O_int8 | 	O_int9 | 	O_int10 	); 
	assign ready_out = ready_in;
	assign valid_out = |valid_out_temp;

endmodule 

module precoder_17_21 (
	input logic  [4 : 0] S ,
	output logic  [31 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		5'd0    :   out_sel = 32'b00000000000000000000000000000001;
		5'd1    :   out_sel = 32'b00000000000000000000000000000010;
		5'd2    :   out_sel = 32'b00000000000000000000000000000100;
		5'd3    :   out_sel = 32'b00000000000000000000000000001000;
		5'd4    :   out_sel = 32'b00000000000000000000000000010000;
		5'd5    :   out_sel = 32'b00000000000000000000000000100000;
		5'd6    :   out_sel = 32'b00000000000000000000000001000000;
		5'd7    :   out_sel = 32'b00000000000000000000000010000000;
		5'd8    :   out_sel = 32'b00000000000000000000000100000000;
		5'd9    :   out_sel = 32'b00000000000000000000001000000000;
		5'd10    :   out_sel = 32'b00000000000000000000010000000000;
		5'd11    :   out_sel = 32'b00000000000000000000100000000000;
		5'd12    :   out_sel = 32'b00000000000000000001000000000000;
		5'd13    :   out_sel = 32'b00000000000000000010000000000000;
		5'd14    :   out_sel = 32'b00000000000000000100000000000000;
		5'd15    :   out_sel = 32'b00000000000000001000000000000000;
		5'd16    :   out_sel = 32'b00000000000000010000000000000000;
		5'd17    :   out_sel = 32'b00000000000000100000000000000000;
		5'd18    :   out_sel = 32'b00000000000001000000000000000000;
		5'd19    :   out_sel = 32'b00000000000010000000000000000000;
		5'd20    :   out_sel = 32'b00000000000100000000000000000000;
		5'd21    :   out_sel = 32'b00000000001000000000000000000000;
		default :   out_sel = 32'b0;
	endcase 
end 

endmodule 

module mux_logic_17_21 ( 
	input logic  [31 : 0] out_sel,
	input logic  [16 : 0] I0, 
	input logic  [16 : 0] I1, 
	input logic  [16 : 0] I2, 
	input logic  [16 : 0] I3, 
	input logic  [16 : 0] I4, 
	input logic  [16 : 0] I5, 
	input logic  [16 : 0] I6, 
	input logic  [16 : 0] I7, 
	input logic  [16 : 0] I8, 
	input logic  [16 : 0] I9, 
	input logic  [16 : 0] I10, 
	input logic  [16 : 0] I11, 
	input logic  [16 : 0] I12, 
	input logic  [16 : 0] I13, 
	input logic  [16 : 0] I14, 
	input logic  [16 : 0] I15, 
	input logic  [16 : 0] I16, 
	input logic  [16 : 0] I17, 
	input logic  [16 : 0] I18, 
	input logic  [16 : 0] I19, 
	input logic  [16 : 0] I20, 
	input logic [20:0] valid_in,
	output logic [10:0] valid_out,
	output logic  [16 : 0] O0, 
	output logic  [16 : 0] O1, 
	output logic  [16 : 0] O2, 
	output logic  [16 : 0] O3, 
	output logic  [16 : 0] O4, 
	output logic  [16 : 0] O5, 
	output logic  [16 : 0] O6, 
	output logic  [16 : 0] O7, 
	output logic  [16 : 0] O8, 
	output logic  [16 : 0] O9, 
	output logic  [16 : 0] O10); 
	AO_CELL inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	AO_CELL inst_1_0 ( 
	.A1(out_sel[2]), 
	.A2(I2[0]), 
	.B1(out_sel[3]), 
	.B2(I3[0]), 
	.Z(O1[0])); 
	AO_CELL inst_2_0 ( 
	.A1(out_sel[4]), 
	.A2(I4[0]), 
	.B1(out_sel[5]), 
	.B2(I5[0]), 
	.Z(O2[0])); 
	AO_CELL inst_3_0 ( 
	.A1(out_sel[6]), 
	.A2(I6[0]), 
	.B1(out_sel[7]), 
	.B2(I7[0]), 
	.Z(O3[0])); 
	AO_CELL inst_4_0 ( 
	.A1(out_sel[8]), 
	.A2(I8[0]), 
	.B1(out_sel[9]), 
	.B2(I9[0]), 
	.Z(O4[0])); 
	AO_CELL inst_5_0 ( 
	.A1(out_sel[10]), 
	.A2(I10[0]), 
	.B1(out_sel[11]), 
	.B2(I11[0]), 
	.Z(O5[0])); 
	AO_CELL inst_6_0 ( 
	.A1(out_sel[12]), 
	.A2(I12[0]), 
	.B1(out_sel[13]), 
	.B2(I13[0]), 
	.Z(O6[0])); 
	AO_CELL inst_7_0 ( 
	.A1(out_sel[14]), 
	.A2(I14[0]), 
	.B1(out_sel[15]), 
	.B2(I15[0]), 
	.Z(O7[0])); 
	AO_CELL inst_8_0 ( 
	.A1(out_sel[16]), 
	.A2(I16[0]), 
	.B1(out_sel[17]), 
	.B2(I17[0]), 
	.Z(O8[0])); 
	AO_CELL inst_9_0 ( 
	.A1(out_sel[18]), 
	.A2(I18[0]), 
	.B1(out_sel[19]), 
	.B2(I19[0]), 
	.Z(O9[0])); 
	AO_CELL inst_10_0 ( 
	.A1(out_sel[20]), 
	.A2(I20[0]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(O10[0])); 
	AO_CELL inst_0_1 ( 
	.A1(out_sel[0]), 
	.A2(I0[1]), 
	.B1(out_sel[1]), 
	.B2(I1[1]), 
	.Z(O0[1])); 
	AO_CELL inst_1_1 ( 
	.A1(out_sel[2]), 
	.A2(I2[1]), 
	.B1(out_sel[3]), 
	.B2(I3[1]), 
	.Z(O1[1])); 
	AO_CELL inst_2_1 ( 
	.A1(out_sel[4]), 
	.A2(I4[1]), 
	.B1(out_sel[5]), 
	.B2(I5[1]), 
	.Z(O2[1])); 
	AO_CELL inst_3_1 ( 
	.A1(out_sel[6]), 
	.A2(I6[1]), 
	.B1(out_sel[7]), 
	.B2(I7[1]), 
	.Z(O3[1])); 
	AO_CELL inst_4_1 ( 
	.A1(out_sel[8]), 
	.A2(I8[1]), 
	.B1(out_sel[9]), 
	.B2(I9[1]), 
	.Z(O4[1])); 
	AO_CELL inst_5_1 ( 
	.A1(out_sel[10]), 
	.A2(I10[1]), 
	.B1(out_sel[11]), 
	.B2(I11[1]), 
	.Z(O5[1])); 
	AO_CELL inst_6_1 ( 
	.A1(out_sel[12]), 
	.A2(I12[1]), 
	.B1(out_sel[13]), 
	.B2(I13[1]), 
	.Z(O6[1])); 
	AO_CELL inst_7_1 ( 
	.A1(out_sel[14]), 
	.A2(I14[1]), 
	.B1(out_sel[15]), 
	.B2(I15[1]), 
	.Z(O7[1])); 
	AO_CELL inst_8_1 ( 
	.A1(out_sel[16]), 
	.A2(I16[1]), 
	.B1(out_sel[17]), 
	.B2(I17[1]), 
	.Z(O8[1])); 
	AO_CELL inst_9_1 ( 
	.A1(out_sel[18]), 
	.A2(I18[1]), 
	.B1(out_sel[19]), 
	.B2(I19[1]), 
	.Z(O9[1])); 
	AO_CELL inst_10_1 ( 
	.A1(out_sel[20]), 
	.A2(I20[1]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(O10[1])); 
	AO_CELL inst_0_2 ( 
	.A1(out_sel[0]), 
	.A2(I0[2]), 
	.B1(out_sel[1]), 
	.B2(I1[2]), 
	.Z(O0[2])); 
	AO_CELL inst_1_2 ( 
	.A1(out_sel[2]), 
	.A2(I2[2]), 
	.B1(out_sel[3]), 
	.B2(I3[2]), 
	.Z(O1[2])); 
	AO_CELL inst_2_2 ( 
	.A1(out_sel[4]), 
	.A2(I4[2]), 
	.B1(out_sel[5]), 
	.B2(I5[2]), 
	.Z(O2[2])); 
	AO_CELL inst_3_2 ( 
	.A1(out_sel[6]), 
	.A2(I6[2]), 
	.B1(out_sel[7]), 
	.B2(I7[2]), 
	.Z(O3[2])); 
	AO_CELL inst_4_2 ( 
	.A1(out_sel[8]), 
	.A2(I8[2]), 
	.B1(out_sel[9]), 
	.B2(I9[2]), 
	.Z(O4[2])); 
	AO_CELL inst_5_2 ( 
	.A1(out_sel[10]), 
	.A2(I10[2]), 
	.B1(out_sel[11]), 
	.B2(I11[2]), 
	.Z(O5[2])); 
	AO_CELL inst_6_2 ( 
	.A1(out_sel[12]), 
	.A2(I12[2]), 
	.B1(out_sel[13]), 
	.B2(I13[2]), 
	.Z(O6[2])); 
	AO_CELL inst_7_2 ( 
	.A1(out_sel[14]), 
	.A2(I14[2]), 
	.B1(out_sel[15]), 
	.B2(I15[2]), 
	.Z(O7[2])); 
	AO_CELL inst_8_2 ( 
	.A1(out_sel[16]), 
	.A2(I16[2]), 
	.B1(out_sel[17]), 
	.B2(I17[2]), 
	.Z(O8[2])); 
	AO_CELL inst_9_2 ( 
	.A1(out_sel[18]), 
	.A2(I18[2]), 
	.B1(out_sel[19]), 
	.B2(I19[2]), 
	.Z(O9[2])); 
	AO_CELL inst_10_2 ( 
	.A1(out_sel[20]), 
	.A2(I20[2]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(O10[2])); 
	AO_CELL inst_0_3 ( 
	.A1(out_sel[0]), 
	.A2(I0[3]), 
	.B1(out_sel[1]), 
	.B2(I1[3]), 
	.Z(O0[3])); 
	AO_CELL inst_1_3 ( 
	.A1(out_sel[2]), 
	.A2(I2[3]), 
	.B1(out_sel[3]), 
	.B2(I3[3]), 
	.Z(O1[3])); 
	AO_CELL inst_2_3 ( 
	.A1(out_sel[4]), 
	.A2(I4[3]), 
	.B1(out_sel[5]), 
	.B2(I5[3]), 
	.Z(O2[3])); 
	AO_CELL inst_3_3 ( 
	.A1(out_sel[6]), 
	.A2(I6[3]), 
	.B1(out_sel[7]), 
	.B2(I7[3]), 
	.Z(O3[3])); 
	AO_CELL inst_4_3 ( 
	.A1(out_sel[8]), 
	.A2(I8[3]), 
	.B1(out_sel[9]), 
	.B2(I9[3]), 
	.Z(O4[3])); 
	AO_CELL inst_5_3 ( 
	.A1(out_sel[10]), 
	.A2(I10[3]), 
	.B1(out_sel[11]), 
	.B2(I11[3]), 
	.Z(O5[3])); 
	AO_CELL inst_6_3 ( 
	.A1(out_sel[12]), 
	.A2(I12[3]), 
	.B1(out_sel[13]), 
	.B2(I13[3]), 
	.Z(O6[3])); 
	AO_CELL inst_7_3 ( 
	.A1(out_sel[14]), 
	.A2(I14[3]), 
	.B1(out_sel[15]), 
	.B2(I15[3]), 
	.Z(O7[3])); 
	AO_CELL inst_8_3 ( 
	.A1(out_sel[16]), 
	.A2(I16[3]), 
	.B1(out_sel[17]), 
	.B2(I17[3]), 
	.Z(O8[3])); 
	AO_CELL inst_9_3 ( 
	.A1(out_sel[18]), 
	.A2(I18[3]), 
	.B1(out_sel[19]), 
	.B2(I19[3]), 
	.Z(O9[3])); 
	AO_CELL inst_10_3 ( 
	.A1(out_sel[20]), 
	.A2(I20[3]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(O10[3])); 
	AO_CELL inst_0_4 ( 
	.A1(out_sel[0]), 
	.A2(I0[4]), 
	.B1(out_sel[1]), 
	.B2(I1[4]), 
	.Z(O0[4])); 
	AO_CELL inst_1_4 ( 
	.A1(out_sel[2]), 
	.A2(I2[4]), 
	.B1(out_sel[3]), 
	.B2(I3[4]), 
	.Z(O1[4])); 
	AO_CELL inst_2_4 ( 
	.A1(out_sel[4]), 
	.A2(I4[4]), 
	.B1(out_sel[5]), 
	.B2(I5[4]), 
	.Z(O2[4])); 
	AO_CELL inst_3_4 ( 
	.A1(out_sel[6]), 
	.A2(I6[4]), 
	.B1(out_sel[7]), 
	.B2(I7[4]), 
	.Z(O3[4])); 
	AO_CELL inst_4_4 ( 
	.A1(out_sel[8]), 
	.A2(I8[4]), 
	.B1(out_sel[9]), 
	.B2(I9[4]), 
	.Z(O4[4])); 
	AO_CELL inst_5_4 ( 
	.A1(out_sel[10]), 
	.A2(I10[4]), 
	.B1(out_sel[11]), 
	.B2(I11[4]), 
	.Z(O5[4])); 
	AO_CELL inst_6_4 ( 
	.A1(out_sel[12]), 
	.A2(I12[4]), 
	.B1(out_sel[13]), 
	.B2(I13[4]), 
	.Z(O6[4])); 
	AO_CELL inst_7_4 ( 
	.A1(out_sel[14]), 
	.A2(I14[4]), 
	.B1(out_sel[15]), 
	.B2(I15[4]), 
	.Z(O7[4])); 
	AO_CELL inst_8_4 ( 
	.A1(out_sel[16]), 
	.A2(I16[4]), 
	.B1(out_sel[17]), 
	.B2(I17[4]), 
	.Z(O8[4])); 
	AO_CELL inst_9_4 ( 
	.A1(out_sel[18]), 
	.A2(I18[4]), 
	.B1(out_sel[19]), 
	.B2(I19[4]), 
	.Z(O9[4])); 
	AO_CELL inst_10_4 ( 
	.A1(out_sel[20]), 
	.A2(I20[4]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(O10[4])); 
	AO_CELL inst_0_5 ( 
	.A1(out_sel[0]), 
	.A2(I0[5]), 
	.B1(out_sel[1]), 
	.B2(I1[5]), 
	.Z(O0[5])); 
	AO_CELL inst_1_5 ( 
	.A1(out_sel[2]), 
	.A2(I2[5]), 
	.B1(out_sel[3]), 
	.B2(I3[5]), 
	.Z(O1[5])); 
	AO_CELL inst_2_5 ( 
	.A1(out_sel[4]), 
	.A2(I4[5]), 
	.B1(out_sel[5]), 
	.B2(I5[5]), 
	.Z(O2[5])); 
	AO_CELL inst_3_5 ( 
	.A1(out_sel[6]), 
	.A2(I6[5]), 
	.B1(out_sel[7]), 
	.B2(I7[5]), 
	.Z(O3[5])); 
	AO_CELL inst_4_5 ( 
	.A1(out_sel[8]), 
	.A2(I8[5]), 
	.B1(out_sel[9]), 
	.B2(I9[5]), 
	.Z(O4[5])); 
	AO_CELL inst_5_5 ( 
	.A1(out_sel[10]), 
	.A2(I10[5]), 
	.B1(out_sel[11]), 
	.B2(I11[5]), 
	.Z(O5[5])); 
	AO_CELL inst_6_5 ( 
	.A1(out_sel[12]), 
	.A2(I12[5]), 
	.B1(out_sel[13]), 
	.B2(I13[5]), 
	.Z(O6[5])); 
	AO_CELL inst_7_5 ( 
	.A1(out_sel[14]), 
	.A2(I14[5]), 
	.B1(out_sel[15]), 
	.B2(I15[5]), 
	.Z(O7[5])); 
	AO_CELL inst_8_5 ( 
	.A1(out_sel[16]), 
	.A2(I16[5]), 
	.B1(out_sel[17]), 
	.B2(I17[5]), 
	.Z(O8[5])); 
	AO_CELL inst_9_5 ( 
	.A1(out_sel[18]), 
	.A2(I18[5]), 
	.B1(out_sel[19]), 
	.B2(I19[5]), 
	.Z(O9[5])); 
	AO_CELL inst_10_5 ( 
	.A1(out_sel[20]), 
	.A2(I20[5]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(O10[5])); 
	AO_CELL inst_0_6 ( 
	.A1(out_sel[0]), 
	.A2(I0[6]), 
	.B1(out_sel[1]), 
	.B2(I1[6]), 
	.Z(O0[6])); 
	AO_CELL inst_1_6 ( 
	.A1(out_sel[2]), 
	.A2(I2[6]), 
	.B1(out_sel[3]), 
	.B2(I3[6]), 
	.Z(O1[6])); 
	AO_CELL inst_2_6 ( 
	.A1(out_sel[4]), 
	.A2(I4[6]), 
	.B1(out_sel[5]), 
	.B2(I5[6]), 
	.Z(O2[6])); 
	AO_CELL inst_3_6 ( 
	.A1(out_sel[6]), 
	.A2(I6[6]), 
	.B1(out_sel[7]), 
	.B2(I7[6]), 
	.Z(O3[6])); 
	AO_CELL inst_4_6 ( 
	.A1(out_sel[8]), 
	.A2(I8[6]), 
	.B1(out_sel[9]), 
	.B2(I9[6]), 
	.Z(O4[6])); 
	AO_CELL inst_5_6 ( 
	.A1(out_sel[10]), 
	.A2(I10[6]), 
	.B1(out_sel[11]), 
	.B2(I11[6]), 
	.Z(O5[6])); 
	AO_CELL inst_6_6 ( 
	.A1(out_sel[12]), 
	.A2(I12[6]), 
	.B1(out_sel[13]), 
	.B2(I13[6]), 
	.Z(O6[6])); 
	AO_CELL inst_7_6 ( 
	.A1(out_sel[14]), 
	.A2(I14[6]), 
	.B1(out_sel[15]), 
	.B2(I15[6]), 
	.Z(O7[6])); 
	AO_CELL inst_8_6 ( 
	.A1(out_sel[16]), 
	.A2(I16[6]), 
	.B1(out_sel[17]), 
	.B2(I17[6]), 
	.Z(O8[6])); 
	AO_CELL inst_9_6 ( 
	.A1(out_sel[18]), 
	.A2(I18[6]), 
	.B1(out_sel[19]), 
	.B2(I19[6]), 
	.Z(O9[6])); 
	AO_CELL inst_10_6 ( 
	.A1(out_sel[20]), 
	.A2(I20[6]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(O10[6])); 
	AO_CELL inst_0_7 ( 
	.A1(out_sel[0]), 
	.A2(I0[7]), 
	.B1(out_sel[1]), 
	.B2(I1[7]), 
	.Z(O0[7])); 
	AO_CELL inst_1_7 ( 
	.A1(out_sel[2]), 
	.A2(I2[7]), 
	.B1(out_sel[3]), 
	.B2(I3[7]), 
	.Z(O1[7])); 
	AO_CELL inst_2_7 ( 
	.A1(out_sel[4]), 
	.A2(I4[7]), 
	.B1(out_sel[5]), 
	.B2(I5[7]), 
	.Z(O2[7])); 
	AO_CELL inst_3_7 ( 
	.A1(out_sel[6]), 
	.A2(I6[7]), 
	.B1(out_sel[7]), 
	.B2(I7[7]), 
	.Z(O3[7])); 
	AO_CELL inst_4_7 ( 
	.A1(out_sel[8]), 
	.A2(I8[7]), 
	.B1(out_sel[9]), 
	.B2(I9[7]), 
	.Z(O4[7])); 
	AO_CELL inst_5_7 ( 
	.A1(out_sel[10]), 
	.A2(I10[7]), 
	.B1(out_sel[11]), 
	.B2(I11[7]), 
	.Z(O5[7])); 
	AO_CELL inst_6_7 ( 
	.A1(out_sel[12]), 
	.A2(I12[7]), 
	.B1(out_sel[13]), 
	.B2(I13[7]), 
	.Z(O6[7])); 
	AO_CELL inst_7_7 ( 
	.A1(out_sel[14]), 
	.A2(I14[7]), 
	.B1(out_sel[15]), 
	.B2(I15[7]), 
	.Z(O7[7])); 
	AO_CELL inst_8_7 ( 
	.A1(out_sel[16]), 
	.A2(I16[7]), 
	.B1(out_sel[17]), 
	.B2(I17[7]), 
	.Z(O8[7])); 
	AO_CELL inst_9_7 ( 
	.A1(out_sel[18]), 
	.A2(I18[7]), 
	.B1(out_sel[19]), 
	.B2(I19[7]), 
	.Z(O9[7])); 
	AO_CELL inst_10_7 ( 
	.A1(out_sel[20]), 
	.A2(I20[7]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(O10[7])); 
	AO_CELL inst_0_8 ( 
	.A1(out_sel[0]), 
	.A2(I0[8]), 
	.B1(out_sel[1]), 
	.B2(I1[8]), 
	.Z(O0[8])); 
	AO_CELL inst_1_8 ( 
	.A1(out_sel[2]), 
	.A2(I2[8]), 
	.B1(out_sel[3]), 
	.B2(I3[8]), 
	.Z(O1[8])); 
	AO_CELL inst_2_8 ( 
	.A1(out_sel[4]), 
	.A2(I4[8]), 
	.B1(out_sel[5]), 
	.B2(I5[8]), 
	.Z(O2[8])); 
	AO_CELL inst_3_8 ( 
	.A1(out_sel[6]), 
	.A2(I6[8]), 
	.B1(out_sel[7]), 
	.B2(I7[8]), 
	.Z(O3[8])); 
	AO_CELL inst_4_8 ( 
	.A1(out_sel[8]), 
	.A2(I8[8]), 
	.B1(out_sel[9]), 
	.B2(I9[8]), 
	.Z(O4[8])); 
	AO_CELL inst_5_8 ( 
	.A1(out_sel[10]), 
	.A2(I10[8]), 
	.B1(out_sel[11]), 
	.B2(I11[8]), 
	.Z(O5[8])); 
	AO_CELL inst_6_8 ( 
	.A1(out_sel[12]), 
	.A2(I12[8]), 
	.B1(out_sel[13]), 
	.B2(I13[8]), 
	.Z(O6[8])); 
	AO_CELL inst_7_8 ( 
	.A1(out_sel[14]), 
	.A2(I14[8]), 
	.B1(out_sel[15]), 
	.B2(I15[8]), 
	.Z(O7[8])); 
	AO_CELL inst_8_8 ( 
	.A1(out_sel[16]), 
	.A2(I16[8]), 
	.B1(out_sel[17]), 
	.B2(I17[8]), 
	.Z(O8[8])); 
	AO_CELL inst_9_8 ( 
	.A1(out_sel[18]), 
	.A2(I18[8]), 
	.B1(out_sel[19]), 
	.B2(I19[8]), 
	.Z(O9[8])); 
	AO_CELL inst_10_8 ( 
	.A1(out_sel[20]), 
	.A2(I20[8]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(O10[8])); 
	AO_CELL inst_0_9 ( 
	.A1(out_sel[0]), 
	.A2(I0[9]), 
	.B1(out_sel[1]), 
	.B2(I1[9]), 
	.Z(O0[9])); 
	AO_CELL inst_1_9 ( 
	.A1(out_sel[2]), 
	.A2(I2[9]), 
	.B1(out_sel[3]), 
	.B2(I3[9]), 
	.Z(O1[9])); 
	AO_CELL inst_2_9 ( 
	.A1(out_sel[4]), 
	.A2(I4[9]), 
	.B1(out_sel[5]), 
	.B2(I5[9]), 
	.Z(O2[9])); 
	AO_CELL inst_3_9 ( 
	.A1(out_sel[6]), 
	.A2(I6[9]), 
	.B1(out_sel[7]), 
	.B2(I7[9]), 
	.Z(O3[9])); 
	AO_CELL inst_4_9 ( 
	.A1(out_sel[8]), 
	.A2(I8[9]), 
	.B1(out_sel[9]), 
	.B2(I9[9]), 
	.Z(O4[9])); 
	AO_CELL inst_5_9 ( 
	.A1(out_sel[10]), 
	.A2(I10[9]), 
	.B1(out_sel[11]), 
	.B2(I11[9]), 
	.Z(O5[9])); 
	AO_CELL inst_6_9 ( 
	.A1(out_sel[12]), 
	.A2(I12[9]), 
	.B1(out_sel[13]), 
	.B2(I13[9]), 
	.Z(O6[9])); 
	AO_CELL inst_7_9 ( 
	.A1(out_sel[14]), 
	.A2(I14[9]), 
	.B1(out_sel[15]), 
	.B2(I15[9]), 
	.Z(O7[9])); 
	AO_CELL inst_8_9 ( 
	.A1(out_sel[16]), 
	.A2(I16[9]), 
	.B1(out_sel[17]), 
	.B2(I17[9]), 
	.Z(O8[9])); 
	AO_CELL inst_9_9 ( 
	.A1(out_sel[18]), 
	.A2(I18[9]), 
	.B1(out_sel[19]), 
	.B2(I19[9]), 
	.Z(O9[9])); 
	AO_CELL inst_10_9 ( 
	.A1(out_sel[20]), 
	.A2(I20[9]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(O10[9])); 
	AO_CELL inst_0_10 ( 
	.A1(out_sel[0]), 
	.A2(I0[10]), 
	.B1(out_sel[1]), 
	.B2(I1[10]), 
	.Z(O0[10])); 
	AO_CELL inst_1_10 ( 
	.A1(out_sel[2]), 
	.A2(I2[10]), 
	.B1(out_sel[3]), 
	.B2(I3[10]), 
	.Z(O1[10])); 
	AO_CELL inst_2_10 ( 
	.A1(out_sel[4]), 
	.A2(I4[10]), 
	.B1(out_sel[5]), 
	.B2(I5[10]), 
	.Z(O2[10])); 
	AO_CELL inst_3_10 ( 
	.A1(out_sel[6]), 
	.A2(I6[10]), 
	.B1(out_sel[7]), 
	.B2(I7[10]), 
	.Z(O3[10])); 
	AO_CELL inst_4_10 ( 
	.A1(out_sel[8]), 
	.A2(I8[10]), 
	.B1(out_sel[9]), 
	.B2(I9[10]), 
	.Z(O4[10])); 
	AO_CELL inst_5_10 ( 
	.A1(out_sel[10]), 
	.A2(I10[10]), 
	.B1(out_sel[11]), 
	.B2(I11[10]), 
	.Z(O5[10])); 
	AO_CELL inst_6_10 ( 
	.A1(out_sel[12]), 
	.A2(I12[10]), 
	.B1(out_sel[13]), 
	.B2(I13[10]), 
	.Z(O6[10])); 
	AO_CELL inst_7_10 ( 
	.A1(out_sel[14]), 
	.A2(I14[10]), 
	.B1(out_sel[15]), 
	.B2(I15[10]), 
	.Z(O7[10])); 
	AO_CELL inst_8_10 ( 
	.A1(out_sel[16]), 
	.A2(I16[10]), 
	.B1(out_sel[17]), 
	.B2(I17[10]), 
	.Z(O8[10])); 
	AO_CELL inst_9_10 ( 
	.A1(out_sel[18]), 
	.A2(I18[10]), 
	.B1(out_sel[19]), 
	.B2(I19[10]), 
	.Z(O9[10])); 
	AO_CELL inst_10_10 ( 
	.A1(out_sel[20]), 
	.A2(I20[10]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(O10[10])); 
	AO_CELL inst_0_11 ( 
	.A1(out_sel[0]), 
	.A2(I0[11]), 
	.B1(out_sel[1]), 
	.B2(I1[11]), 
	.Z(O0[11])); 
	AO_CELL inst_1_11 ( 
	.A1(out_sel[2]), 
	.A2(I2[11]), 
	.B1(out_sel[3]), 
	.B2(I3[11]), 
	.Z(O1[11])); 
	AO_CELL inst_2_11 ( 
	.A1(out_sel[4]), 
	.A2(I4[11]), 
	.B1(out_sel[5]), 
	.B2(I5[11]), 
	.Z(O2[11])); 
	AO_CELL inst_3_11 ( 
	.A1(out_sel[6]), 
	.A2(I6[11]), 
	.B1(out_sel[7]), 
	.B2(I7[11]), 
	.Z(O3[11])); 
	AO_CELL inst_4_11 ( 
	.A1(out_sel[8]), 
	.A2(I8[11]), 
	.B1(out_sel[9]), 
	.B2(I9[11]), 
	.Z(O4[11])); 
	AO_CELL inst_5_11 ( 
	.A1(out_sel[10]), 
	.A2(I10[11]), 
	.B1(out_sel[11]), 
	.B2(I11[11]), 
	.Z(O5[11])); 
	AO_CELL inst_6_11 ( 
	.A1(out_sel[12]), 
	.A2(I12[11]), 
	.B1(out_sel[13]), 
	.B2(I13[11]), 
	.Z(O6[11])); 
	AO_CELL inst_7_11 ( 
	.A1(out_sel[14]), 
	.A2(I14[11]), 
	.B1(out_sel[15]), 
	.B2(I15[11]), 
	.Z(O7[11])); 
	AO_CELL inst_8_11 ( 
	.A1(out_sel[16]), 
	.A2(I16[11]), 
	.B1(out_sel[17]), 
	.B2(I17[11]), 
	.Z(O8[11])); 
	AO_CELL inst_9_11 ( 
	.A1(out_sel[18]), 
	.A2(I18[11]), 
	.B1(out_sel[19]), 
	.B2(I19[11]), 
	.Z(O9[11])); 
	AO_CELL inst_10_11 ( 
	.A1(out_sel[20]), 
	.A2(I20[11]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(O10[11])); 
	AO_CELL inst_0_12 ( 
	.A1(out_sel[0]), 
	.A2(I0[12]), 
	.B1(out_sel[1]), 
	.B2(I1[12]), 
	.Z(O0[12])); 
	AO_CELL inst_1_12 ( 
	.A1(out_sel[2]), 
	.A2(I2[12]), 
	.B1(out_sel[3]), 
	.B2(I3[12]), 
	.Z(O1[12])); 
	AO_CELL inst_2_12 ( 
	.A1(out_sel[4]), 
	.A2(I4[12]), 
	.B1(out_sel[5]), 
	.B2(I5[12]), 
	.Z(O2[12])); 
	AO_CELL inst_3_12 ( 
	.A1(out_sel[6]), 
	.A2(I6[12]), 
	.B1(out_sel[7]), 
	.B2(I7[12]), 
	.Z(O3[12])); 
	AO_CELL inst_4_12 ( 
	.A1(out_sel[8]), 
	.A2(I8[12]), 
	.B1(out_sel[9]), 
	.B2(I9[12]), 
	.Z(O4[12])); 
	AO_CELL inst_5_12 ( 
	.A1(out_sel[10]), 
	.A2(I10[12]), 
	.B1(out_sel[11]), 
	.B2(I11[12]), 
	.Z(O5[12])); 
	AO_CELL inst_6_12 ( 
	.A1(out_sel[12]), 
	.A2(I12[12]), 
	.B1(out_sel[13]), 
	.B2(I13[12]), 
	.Z(O6[12])); 
	AO_CELL inst_7_12 ( 
	.A1(out_sel[14]), 
	.A2(I14[12]), 
	.B1(out_sel[15]), 
	.B2(I15[12]), 
	.Z(O7[12])); 
	AO_CELL inst_8_12 ( 
	.A1(out_sel[16]), 
	.A2(I16[12]), 
	.B1(out_sel[17]), 
	.B2(I17[12]), 
	.Z(O8[12])); 
	AO_CELL inst_9_12 ( 
	.A1(out_sel[18]), 
	.A2(I18[12]), 
	.B1(out_sel[19]), 
	.B2(I19[12]), 
	.Z(O9[12])); 
	AO_CELL inst_10_12 ( 
	.A1(out_sel[20]), 
	.A2(I20[12]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(O10[12])); 
	AO_CELL inst_0_13 ( 
	.A1(out_sel[0]), 
	.A2(I0[13]), 
	.B1(out_sel[1]), 
	.B2(I1[13]), 
	.Z(O0[13])); 
	AO_CELL inst_1_13 ( 
	.A1(out_sel[2]), 
	.A2(I2[13]), 
	.B1(out_sel[3]), 
	.B2(I3[13]), 
	.Z(O1[13])); 
	AO_CELL inst_2_13 ( 
	.A1(out_sel[4]), 
	.A2(I4[13]), 
	.B1(out_sel[5]), 
	.B2(I5[13]), 
	.Z(O2[13])); 
	AO_CELL inst_3_13 ( 
	.A1(out_sel[6]), 
	.A2(I6[13]), 
	.B1(out_sel[7]), 
	.B2(I7[13]), 
	.Z(O3[13])); 
	AO_CELL inst_4_13 ( 
	.A1(out_sel[8]), 
	.A2(I8[13]), 
	.B1(out_sel[9]), 
	.B2(I9[13]), 
	.Z(O4[13])); 
	AO_CELL inst_5_13 ( 
	.A1(out_sel[10]), 
	.A2(I10[13]), 
	.B1(out_sel[11]), 
	.B2(I11[13]), 
	.Z(O5[13])); 
	AO_CELL inst_6_13 ( 
	.A1(out_sel[12]), 
	.A2(I12[13]), 
	.B1(out_sel[13]), 
	.B2(I13[13]), 
	.Z(O6[13])); 
	AO_CELL inst_7_13 ( 
	.A1(out_sel[14]), 
	.A2(I14[13]), 
	.B1(out_sel[15]), 
	.B2(I15[13]), 
	.Z(O7[13])); 
	AO_CELL inst_8_13 ( 
	.A1(out_sel[16]), 
	.A2(I16[13]), 
	.B1(out_sel[17]), 
	.B2(I17[13]), 
	.Z(O8[13])); 
	AO_CELL inst_9_13 ( 
	.A1(out_sel[18]), 
	.A2(I18[13]), 
	.B1(out_sel[19]), 
	.B2(I19[13]), 
	.Z(O9[13])); 
	AO_CELL inst_10_13 ( 
	.A1(out_sel[20]), 
	.A2(I20[13]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(O10[13])); 
	AO_CELL inst_0_14 ( 
	.A1(out_sel[0]), 
	.A2(I0[14]), 
	.B1(out_sel[1]), 
	.B2(I1[14]), 
	.Z(O0[14])); 
	AO_CELL inst_1_14 ( 
	.A1(out_sel[2]), 
	.A2(I2[14]), 
	.B1(out_sel[3]), 
	.B2(I3[14]), 
	.Z(O1[14])); 
	AO_CELL inst_2_14 ( 
	.A1(out_sel[4]), 
	.A2(I4[14]), 
	.B1(out_sel[5]), 
	.B2(I5[14]), 
	.Z(O2[14])); 
	AO_CELL inst_3_14 ( 
	.A1(out_sel[6]), 
	.A2(I6[14]), 
	.B1(out_sel[7]), 
	.B2(I7[14]), 
	.Z(O3[14])); 
	AO_CELL inst_4_14 ( 
	.A1(out_sel[8]), 
	.A2(I8[14]), 
	.B1(out_sel[9]), 
	.B2(I9[14]), 
	.Z(O4[14])); 
	AO_CELL inst_5_14 ( 
	.A1(out_sel[10]), 
	.A2(I10[14]), 
	.B1(out_sel[11]), 
	.B2(I11[14]), 
	.Z(O5[14])); 
	AO_CELL inst_6_14 ( 
	.A1(out_sel[12]), 
	.A2(I12[14]), 
	.B1(out_sel[13]), 
	.B2(I13[14]), 
	.Z(O6[14])); 
	AO_CELL inst_7_14 ( 
	.A1(out_sel[14]), 
	.A2(I14[14]), 
	.B1(out_sel[15]), 
	.B2(I15[14]), 
	.Z(O7[14])); 
	AO_CELL inst_8_14 ( 
	.A1(out_sel[16]), 
	.A2(I16[14]), 
	.B1(out_sel[17]), 
	.B2(I17[14]), 
	.Z(O8[14])); 
	AO_CELL inst_9_14 ( 
	.A1(out_sel[18]), 
	.A2(I18[14]), 
	.B1(out_sel[19]), 
	.B2(I19[14]), 
	.Z(O9[14])); 
	AO_CELL inst_10_14 ( 
	.A1(out_sel[20]), 
	.A2(I20[14]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(O10[14])); 
	AO_CELL inst_0_15 ( 
	.A1(out_sel[0]), 
	.A2(I0[15]), 
	.B1(out_sel[1]), 
	.B2(I1[15]), 
	.Z(O0[15])); 
	AO_CELL inst_1_15 ( 
	.A1(out_sel[2]), 
	.A2(I2[15]), 
	.B1(out_sel[3]), 
	.B2(I3[15]), 
	.Z(O1[15])); 
	AO_CELL inst_2_15 ( 
	.A1(out_sel[4]), 
	.A2(I4[15]), 
	.B1(out_sel[5]), 
	.B2(I5[15]), 
	.Z(O2[15])); 
	AO_CELL inst_3_15 ( 
	.A1(out_sel[6]), 
	.A2(I6[15]), 
	.B1(out_sel[7]), 
	.B2(I7[15]), 
	.Z(O3[15])); 
	AO_CELL inst_4_15 ( 
	.A1(out_sel[8]), 
	.A2(I8[15]), 
	.B1(out_sel[9]), 
	.B2(I9[15]), 
	.Z(O4[15])); 
	AO_CELL inst_5_15 ( 
	.A1(out_sel[10]), 
	.A2(I10[15]), 
	.B1(out_sel[11]), 
	.B2(I11[15]), 
	.Z(O5[15])); 
	AO_CELL inst_6_15 ( 
	.A1(out_sel[12]), 
	.A2(I12[15]), 
	.B1(out_sel[13]), 
	.B2(I13[15]), 
	.Z(O6[15])); 
	AO_CELL inst_7_15 ( 
	.A1(out_sel[14]), 
	.A2(I14[15]), 
	.B1(out_sel[15]), 
	.B2(I15[15]), 
	.Z(O7[15])); 
	AO_CELL inst_8_15 ( 
	.A1(out_sel[16]), 
	.A2(I16[15]), 
	.B1(out_sel[17]), 
	.B2(I17[15]), 
	.Z(O8[15])); 
	AO_CELL inst_9_15 ( 
	.A1(out_sel[18]), 
	.A2(I18[15]), 
	.B1(out_sel[19]), 
	.B2(I19[15]), 
	.Z(O9[15])); 
	AO_CELL inst_10_15 ( 
	.A1(out_sel[20]), 
	.A2(I20[15]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(O10[15])); 
	AO_CELL inst_0_16 ( 
	.A1(out_sel[0]), 
	.A2(I0[16]), 
	.B1(out_sel[1]), 
	.B2(I1[16]), 
	.Z(O0[16])); 
	AO_CELL inst_1_16 ( 
	.A1(out_sel[2]), 
	.A2(I2[16]), 
	.B1(out_sel[3]), 
	.B2(I3[16]), 
	.Z(O1[16])); 
	AO_CELL inst_2_16 ( 
	.A1(out_sel[4]), 
	.A2(I4[16]), 
	.B1(out_sel[5]), 
	.B2(I5[16]), 
	.Z(O2[16])); 
	AO_CELL inst_3_16 ( 
	.A1(out_sel[6]), 
	.A2(I6[16]), 
	.B1(out_sel[7]), 
	.B2(I7[16]), 
	.Z(O3[16])); 
	AO_CELL inst_4_16 ( 
	.A1(out_sel[8]), 
	.A2(I8[16]), 
	.B1(out_sel[9]), 
	.B2(I9[16]), 
	.Z(O4[16])); 
	AO_CELL inst_5_16 ( 
	.A1(out_sel[10]), 
	.A2(I10[16]), 
	.B1(out_sel[11]), 
	.B2(I11[16]), 
	.Z(O5[16])); 
	AO_CELL inst_6_16 ( 
	.A1(out_sel[12]), 
	.A2(I12[16]), 
	.B1(out_sel[13]), 
	.B2(I13[16]), 
	.Z(O6[16])); 
	AO_CELL inst_7_16 ( 
	.A1(out_sel[14]), 
	.A2(I14[16]), 
	.B1(out_sel[15]), 
	.B2(I15[16]), 
	.Z(O7[16])); 
	AO_CELL inst_8_16 ( 
	.A1(out_sel[16]), 
	.A2(I16[16]), 
	.B1(out_sel[17]), 
	.B2(I17[16]), 
	.Z(O8[16])); 
	AO_CELL inst_9_16 ( 
	.A1(out_sel[18]), 
	.A2(I18[16]), 
	.B1(out_sel[19]), 
	.B2(I19[16]), 
	.Z(O9[16])); 
	AO_CELL inst_10_16 ( 
	.A1(out_sel[20]), 
	.A2(I20[16]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(O10[16])); 
	AO_CELL inst_0_valid ( 
	.A1(out_sel[0]), 
	.A2(valid_in[0]), 
	.B1(out_sel[1]), 
	.B2(valid_in[1]), 
	.Z(valid_out[0])); 
	AO_CELL inst_1_valid ( 
	.A1(out_sel[2]), 
	.A2(valid_in[2]), 
	.B1(out_sel[3]), 
	.B2(valid_in[3]), 
	.Z(valid_out[1])); 
	AO_CELL inst_2_valid ( 
	.A1(out_sel[4]), 
	.A2(valid_in[4]), 
	.B1(out_sel[5]), 
	.B2(valid_in[5]), 
	.Z(valid_out[2])); 
	AO_CELL inst_3_valid ( 
	.A1(out_sel[6]), 
	.A2(valid_in[6]), 
	.B1(out_sel[7]), 
	.B2(valid_in[7]), 
	.Z(valid_out[3])); 
	AO_CELL inst_4_valid ( 
	.A1(out_sel[8]), 
	.A2(valid_in[8]), 
	.B1(out_sel[9]), 
	.B2(valid_in[9]), 
	.Z(valid_out[4])); 
	AO_CELL inst_5_valid ( 
	.A1(out_sel[10]), 
	.A2(valid_in[10]), 
	.B1(out_sel[11]), 
	.B2(valid_in[11]), 
	.Z(valid_out[5])); 
	AO_CELL inst_6_valid ( 
	.A1(out_sel[12]), 
	.A2(valid_in[12]), 
	.B1(out_sel[13]), 
	.B2(valid_in[13]), 
	.Z(valid_out[6])); 
	AO_CELL inst_7_valid ( 
	.A1(out_sel[14]), 
	.A2(valid_in[14]), 
	.B1(out_sel[15]), 
	.B2(valid_in[15]), 
	.Z(valid_out[7])); 
	AO_CELL inst_8_valid ( 
	.A1(out_sel[16]), 
	.A2(valid_in[16]), 
	.B1(out_sel[17]), 
	.B2(valid_in[17]), 
	.Z(valid_out[8])); 
	AO_CELL inst_9_valid ( 
	.A1(out_sel[18]), 
	.A2(valid_in[18]), 
	.B1(out_sel[19]), 
	.B2(valid_in[19]), 
	.Z(valid_out[9])); 
	AO_CELL inst_10_valid ( 
	.A1(out_sel[20]), 
	.A2(valid_in[20]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(valid_out[10])); 
endmodule 

module mux_aoi_ready_valid_const_21_1 ( 
	input logic  [0 : 0] I[20:0], 
	input logic  [4 : 0] S ,
	input logic ready_in,
	output logic ready_out,
	input logic [20:0]  valid_in,
	output logic valid_out,
	output logic  [31 : 0] out_sel,
	output logic [0 : 0] O); 
	logic  [0 : 0] O_int0;
	logic  [0 : 0] O_int1;
	logic  [0 : 0] O_int2;
	logic  [0 : 0] O_int3;
	logic  [0 : 0] O_int4;
	logic  [0 : 0] O_int5;
	logic  [0 : 0] O_int6;
	logic  [0 : 0] O_int7;
	logic  [0 : 0] O_int8;
	logic  [0 : 0] O_int9;
	logic  [0 : 0] O_int10;
	logic [10:0] valid_out_temp;

precoder_1_21 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_1_21 u_mux_logic ( 
	.I0 (I[0]),
	.I1 (I[1]),
	.I2 (I[2]),
	.I3 (I[3]),
	.I4 (I[4]),
	.I5 (I[5]),
	.I6 (I[6]),
	.I7 (I[7]),
	.I8 (I[8]),
	.I9 (I[9]),
	.I10 (I[10]),
	.I11 (I[11]),
	.I12 (I[12]),
	.I13 (I[13]),
	.I14 (I[14]),
	.I15 (I[15]),
	.I16 (I[16]),
	.I17 (I[17]),
	.I18 (I[18]),
	.I19 (I[19]),
	.I20 (I[20]),
	.out_sel(out_sel), 
	.valid_in(valid_in),
	.valid_out(valid_out_temp),
	.O0(O_int0), 
	.O1(O_int1), 
	.O2(O_int2), 
	.O3(O_int3), 
	.O4(O_int4), 
	.O5(O_int5), 
	.O6(O_int6), 
	.O7(O_int7), 
	.O8(O_int8), 
	.O9(O_int9), 
	.O10(O_int10)); 
	assign O = (  	O_int0 | 	O_int1 | 	O_int2 | 	O_int3 | 	O_int4 | 	O_int5 | 	O_int6 | 	O_int7 | 	O_int8 | 	O_int9 | 	O_int10 	); 
	assign ready_out = ready_in;
	assign valid_out = |valid_out_temp;

endmodule 

module precoder_1_21 (
	input logic  [4 : 0] S ,
	output logic  [31 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		5'd0    :   out_sel = 32'b00000000000000000000000000000001;
		5'd1    :   out_sel = 32'b00000000000000000000000000000010;
		5'd2    :   out_sel = 32'b00000000000000000000000000000100;
		5'd3    :   out_sel = 32'b00000000000000000000000000001000;
		5'd4    :   out_sel = 32'b00000000000000000000000000010000;
		5'd5    :   out_sel = 32'b00000000000000000000000000100000;
		5'd6    :   out_sel = 32'b00000000000000000000000001000000;
		5'd7    :   out_sel = 32'b00000000000000000000000010000000;
		5'd8    :   out_sel = 32'b00000000000000000000000100000000;
		5'd9    :   out_sel = 32'b00000000000000000000001000000000;
		5'd10    :   out_sel = 32'b00000000000000000000010000000000;
		5'd11    :   out_sel = 32'b00000000000000000000100000000000;
		5'd12    :   out_sel = 32'b00000000000000000001000000000000;
		5'd13    :   out_sel = 32'b00000000000000000010000000000000;
		5'd14    :   out_sel = 32'b00000000000000000100000000000000;
		5'd15    :   out_sel = 32'b00000000000000001000000000000000;
		5'd16    :   out_sel = 32'b00000000000000010000000000000000;
		5'd17    :   out_sel = 32'b00000000000000100000000000000000;
		5'd18    :   out_sel = 32'b00000000000001000000000000000000;
		5'd19    :   out_sel = 32'b00000000000010000000000000000000;
		5'd20    :   out_sel = 32'b00000000000100000000000000000000;
		5'd21    :   out_sel = 32'b00000000001000000000000000000000;
		default :   out_sel = 32'b0;
	endcase 
end 

endmodule 

module mux_logic_1_21 ( 
	input logic  [31 : 0] out_sel,
	input logic  [0 : 0] I0, 
	input logic  [0 : 0] I1, 
	input logic  [0 : 0] I2, 
	input logic  [0 : 0] I3, 
	input logic  [0 : 0] I4, 
	input logic  [0 : 0] I5, 
	input logic  [0 : 0] I6, 
	input logic  [0 : 0] I7, 
	input logic  [0 : 0] I8, 
	input logic  [0 : 0] I9, 
	input logic  [0 : 0] I10, 
	input logic  [0 : 0] I11, 
	input logic  [0 : 0] I12, 
	input logic  [0 : 0] I13, 
	input logic  [0 : 0] I14, 
	input logic  [0 : 0] I15, 
	input logic  [0 : 0] I16, 
	input logic  [0 : 0] I17, 
	input logic  [0 : 0] I18, 
	input logic  [0 : 0] I19, 
	input logic  [0 : 0] I20, 
	input logic [20:0] valid_in,
	output logic [10:0] valid_out,
	output logic  [0 : 0] O0, 
	output logic  [0 : 0] O1, 
	output logic  [0 : 0] O2, 
	output logic  [0 : 0] O3, 
	output logic  [0 : 0] O4, 
	output logic  [0 : 0] O5, 
	output logic  [0 : 0] O6, 
	output logic  [0 : 0] O7, 
	output logic  [0 : 0] O8, 
	output logic  [0 : 0] O9, 
	output logic  [0 : 0] O10); 
	AO_CELL inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	AO_CELL inst_1_0 ( 
	.A1(out_sel[2]), 
	.A2(I2[0]), 
	.B1(out_sel[3]), 
	.B2(I3[0]), 
	.Z(O1[0])); 
	AO_CELL inst_2_0 ( 
	.A1(out_sel[4]), 
	.A2(I4[0]), 
	.B1(out_sel[5]), 
	.B2(I5[0]), 
	.Z(O2[0])); 
	AO_CELL inst_3_0 ( 
	.A1(out_sel[6]), 
	.A2(I6[0]), 
	.B1(out_sel[7]), 
	.B2(I7[0]), 
	.Z(O3[0])); 
	AO_CELL inst_4_0 ( 
	.A1(out_sel[8]), 
	.A2(I8[0]), 
	.B1(out_sel[9]), 
	.B2(I9[0]), 
	.Z(O4[0])); 
	AO_CELL inst_5_0 ( 
	.A1(out_sel[10]), 
	.A2(I10[0]), 
	.B1(out_sel[11]), 
	.B2(I11[0]), 
	.Z(O5[0])); 
	AO_CELL inst_6_0 ( 
	.A1(out_sel[12]), 
	.A2(I12[0]), 
	.B1(out_sel[13]), 
	.B2(I13[0]), 
	.Z(O6[0])); 
	AO_CELL inst_7_0 ( 
	.A1(out_sel[14]), 
	.A2(I14[0]), 
	.B1(out_sel[15]), 
	.B2(I15[0]), 
	.Z(O7[0])); 
	AO_CELL inst_8_0 ( 
	.A1(out_sel[16]), 
	.A2(I16[0]), 
	.B1(out_sel[17]), 
	.B2(I17[0]), 
	.Z(O8[0])); 
	AO_CELL inst_9_0 ( 
	.A1(out_sel[18]), 
	.A2(I18[0]), 
	.B1(out_sel[19]), 
	.B2(I19[0]), 
	.Z(O9[0])); 
	AO_CELL inst_10_0 ( 
	.A1(out_sel[20]), 
	.A2(I20[0]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(O10[0])); 
	AO_CELL inst_0_valid ( 
	.A1(out_sel[0]), 
	.A2(valid_in[0]), 
	.B1(out_sel[1]), 
	.B2(valid_in[1]), 
	.Z(valid_out[0])); 
	AO_CELL inst_1_valid ( 
	.A1(out_sel[2]), 
	.A2(valid_in[2]), 
	.B1(out_sel[3]), 
	.B2(valid_in[3]), 
	.Z(valid_out[1])); 
	AO_CELL inst_2_valid ( 
	.A1(out_sel[4]), 
	.A2(valid_in[4]), 
	.B1(out_sel[5]), 
	.B2(valid_in[5]), 
	.Z(valid_out[2])); 
	AO_CELL inst_3_valid ( 
	.A1(out_sel[6]), 
	.A2(valid_in[6]), 
	.B1(out_sel[7]), 
	.B2(valid_in[7]), 
	.Z(valid_out[3])); 
	AO_CELL inst_4_valid ( 
	.A1(out_sel[8]), 
	.A2(valid_in[8]), 
	.B1(out_sel[9]), 
	.B2(valid_in[9]), 
	.Z(valid_out[4])); 
	AO_CELL inst_5_valid ( 
	.A1(out_sel[10]), 
	.A2(valid_in[10]), 
	.B1(out_sel[11]), 
	.B2(valid_in[11]), 
	.Z(valid_out[5])); 
	AO_CELL inst_6_valid ( 
	.A1(out_sel[12]), 
	.A2(valid_in[12]), 
	.B1(out_sel[13]), 
	.B2(valid_in[13]), 
	.Z(valid_out[6])); 
	AO_CELL inst_7_valid ( 
	.A1(out_sel[14]), 
	.A2(valid_in[14]), 
	.B1(out_sel[15]), 
	.B2(valid_in[15]), 
	.Z(valid_out[7])); 
	AO_CELL inst_8_valid ( 
	.A1(out_sel[16]), 
	.A2(valid_in[16]), 
	.B1(out_sel[17]), 
	.B2(valid_in[17]), 
	.Z(valid_out[8])); 
	AO_CELL inst_9_valid ( 
	.A1(out_sel[18]), 
	.A2(valid_in[18]), 
	.B1(out_sel[19]), 
	.B2(valid_in[19]), 
	.Z(valid_out[9])); 
	AO_CELL inst_10_valid ( 
	.A1(out_sel[20]), 
	.A2(valid_in[20]), 
	.B1(out_sel[21]), 
	.B2(1'b0), 
	.Z(valid_out[10])); 
endmodule 

module mux_aoi_ready_valid_const_20_17 ( 
	input logic  [16 : 0] I[19:0], 
	input logic  [4 : 0] S ,
	input logic ready_in,
	output logic ready_out,
	input logic [19:0]  valid_in,
	output logic valid_out,
	output logic  [31 : 0] out_sel,
	output logic [16 : 0] O); 
	logic  [16 : 0] O_int0;
	logic  [16 : 0] O_int1;
	logic  [16 : 0] O_int2;
	logic  [16 : 0] O_int3;
	logic  [16 : 0] O_int4;
	logic  [16 : 0] O_int5;
	logic  [16 : 0] O_int6;
	logic  [16 : 0] O_int7;
	logic  [16 : 0] O_int8;
	logic  [16 : 0] O_int9;
	logic  [16 : 0] O_int10;
	logic [10:0] valid_out_temp;

precoder_17_20 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_17_20 u_mux_logic ( 
	.I0 (I[0]),
	.I1 (I[1]),
	.I2 (I[2]),
	.I3 (I[3]),
	.I4 (I[4]),
	.I5 (I[5]),
	.I6 (I[6]),
	.I7 (I[7]),
	.I8 (I[8]),
	.I9 (I[9]),
	.I10 (I[10]),
	.I11 (I[11]),
	.I12 (I[12]),
	.I13 (I[13]),
	.I14 (I[14]),
	.I15 (I[15]),
	.I16 (I[16]),
	.I17 (I[17]),
	.I18 (I[18]),
	.I19 (I[19]),
	.out_sel(out_sel), 
	.valid_in(valid_in),
	.valid_out(valid_out_temp),
	.O0(O_int0), 
	.O1(O_int1), 
	.O2(O_int2), 
	.O3(O_int3), 
	.O4(O_int4), 
	.O5(O_int5), 
	.O6(O_int6), 
	.O7(O_int7), 
	.O8(O_int8), 
	.O9(O_int9), 
	.O10(O_int10)); 
	assign O = (  	O_int0 | 	O_int1 | 	O_int2 | 	O_int3 | 	O_int4 | 	O_int5 | 	O_int6 | 	O_int7 | 	O_int8 | 	O_int9 | 	O_int10 	); 
	assign ready_out = ready_in;
	assign valid_out = |valid_out_temp;

endmodule 

module precoder_17_20 (
	input logic  [4 : 0] S ,
	output logic  [31 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		5'd0    :   out_sel = 32'b00000000000000000000000000000001;
		5'd1    :   out_sel = 32'b00000000000000000000000000000010;
		5'd2    :   out_sel = 32'b00000000000000000000000000000100;
		5'd3    :   out_sel = 32'b00000000000000000000000000001000;
		5'd4    :   out_sel = 32'b00000000000000000000000000010000;
		5'd5    :   out_sel = 32'b00000000000000000000000000100000;
		5'd6    :   out_sel = 32'b00000000000000000000000001000000;
		5'd7    :   out_sel = 32'b00000000000000000000000010000000;
		5'd8    :   out_sel = 32'b00000000000000000000000100000000;
		5'd9    :   out_sel = 32'b00000000000000000000001000000000;
		5'd10    :   out_sel = 32'b00000000000000000000010000000000;
		5'd11    :   out_sel = 32'b00000000000000000000100000000000;
		5'd12    :   out_sel = 32'b00000000000000000001000000000000;
		5'd13    :   out_sel = 32'b00000000000000000010000000000000;
		5'd14    :   out_sel = 32'b00000000000000000100000000000000;
		5'd15    :   out_sel = 32'b00000000000000001000000000000000;
		5'd16    :   out_sel = 32'b00000000000000010000000000000000;
		5'd17    :   out_sel = 32'b00000000000000100000000000000000;
		5'd18    :   out_sel = 32'b00000000000001000000000000000000;
		5'd19    :   out_sel = 32'b00000000000010000000000000000000;
		5'd20    :   out_sel = 32'b00000000000100000000000000000000;
		default :   out_sel = 32'b0;
	endcase 
end 

endmodule 

module mux_logic_17_20 ( 
	input logic  [31 : 0] out_sel,
	input logic  [16 : 0] I0, 
	input logic  [16 : 0] I1, 
	input logic  [16 : 0] I2, 
	input logic  [16 : 0] I3, 
	input logic  [16 : 0] I4, 
	input logic  [16 : 0] I5, 
	input logic  [16 : 0] I6, 
	input logic  [16 : 0] I7, 
	input logic  [16 : 0] I8, 
	input logic  [16 : 0] I9, 
	input logic  [16 : 0] I10, 
	input logic  [16 : 0] I11, 
	input logic  [16 : 0] I12, 
	input logic  [16 : 0] I13, 
	input logic  [16 : 0] I14, 
	input logic  [16 : 0] I15, 
	input logic  [16 : 0] I16, 
	input logic  [16 : 0] I17, 
	input logic  [16 : 0] I18, 
	input logic  [16 : 0] I19, 
	input logic [19:0] valid_in,
	output logic [10:0] valid_out,
	output logic  [16 : 0] O0, 
	output logic  [16 : 0] O1, 
	output logic  [16 : 0] O2, 
	output logic  [16 : 0] O3, 
	output logic  [16 : 0] O4, 
	output logic  [16 : 0] O5, 
	output logic  [16 : 0] O6, 
	output logic  [16 : 0] O7, 
	output logic  [16 : 0] O8, 
	output logic  [16 : 0] O9, 
	output logic  [16 : 0] O10); 
	AO_CELL inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	AO_CELL inst_1_0 ( 
	.A1(out_sel[2]), 
	.A2(I2[0]), 
	.B1(out_sel[3]), 
	.B2(I3[0]), 
	.Z(O1[0])); 
	AO_CELL inst_2_0 ( 
	.A1(out_sel[4]), 
	.A2(I4[0]), 
	.B1(out_sel[5]), 
	.B2(I5[0]), 
	.Z(O2[0])); 
	AO_CELL inst_3_0 ( 
	.A1(out_sel[6]), 
	.A2(I6[0]), 
	.B1(out_sel[7]), 
	.B2(I7[0]), 
	.Z(O3[0])); 
	AO_CELL inst_4_0 ( 
	.A1(out_sel[8]), 
	.A2(I8[0]), 
	.B1(out_sel[9]), 
	.B2(I9[0]), 
	.Z(O4[0])); 
	AO_CELL inst_5_0 ( 
	.A1(out_sel[10]), 
	.A2(I10[0]), 
	.B1(out_sel[11]), 
	.B2(I11[0]), 
	.Z(O5[0])); 
	AO_CELL inst_6_0 ( 
	.A1(out_sel[12]), 
	.A2(I12[0]), 
	.B1(out_sel[13]), 
	.B2(I13[0]), 
	.Z(O6[0])); 
	AO_CELL inst_7_0 ( 
	.A1(out_sel[14]), 
	.A2(I14[0]), 
	.B1(out_sel[15]), 
	.B2(I15[0]), 
	.Z(O7[0])); 
	AO_CELL inst_8_0 ( 
	.A1(out_sel[16]), 
	.A2(I16[0]), 
	.B1(out_sel[17]), 
	.B2(I17[0]), 
	.Z(O8[0])); 
	AO_CELL inst_9_0 ( 
	.A1(out_sel[18]), 
	.A2(I18[0]), 
	.B1(out_sel[19]), 
	.B2(I19[0]), 
	.Z(O9[0])); 
	AN_CELL inst_and_0 ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(O10[0])); 
	AO_CELL inst_0_1 ( 
	.A1(out_sel[0]), 
	.A2(I0[1]), 
	.B1(out_sel[1]), 
	.B2(I1[1]), 
	.Z(O0[1])); 
	AO_CELL inst_1_1 ( 
	.A1(out_sel[2]), 
	.A2(I2[1]), 
	.B1(out_sel[3]), 
	.B2(I3[1]), 
	.Z(O1[1])); 
	AO_CELL inst_2_1 ( 
	.A1(out_sel[4]), 
	.A2(I4[1]), 
	.B1(out_sel[5]), 
	.B2(I5[1]), 
	.Z(O2[1])); 
	AO_CELL inst_3_1 ( 
	.A1(out_sel[6]), 
	.A2(I6[1]), 
	.B1(out_sel[7]), 
	.B2(I7[1]), 
	.Z(O3[1])); 
	AO_CELL inst_4_1 ( 
	.A1(out_sel[8]), 
	.A2(I8[1]), 
	.B1(out_sel[9]), 
	.B2(I9[1]), 
	.Z(O4[1])); 
	AO_CELL inst_5_1 ( 
	.A1(out_sel[10]), 
	.A2(I10[1]), 
	.B1(out_sel[11]), 
	.B2(I11[1]), 
	.Z(O5[1])); 
	AO_CELL inst_6_1 ( 
	.A1(out_sel[12]), 
	.A2(I12[1]), 
	.B1(out_sel[13]), 
	.B2(I13[1]), 
	.Z(O6[1])); 
	AO_CELL inst_7_1 ( 
	.A1(out_sel[14]), 
	.A2(I14[1]), 
	.B1(out_sel[15]), 
	.B2(I15[1]), 
	.Z(O7[1])); 
	AO_CELL inst_8_1 ( 
	.A1(out_sel[16]), 
	.A2(I16[1]), 
	.B1(out_sel[17]), 
	.B2(I17[1]), 
	.Z(O8[1])); 
	AO_CELL inst_9_1 ( 
	.A1(out_sel[18]), 
	.A2(I18[1]), 
	.B1(out_sel[19]), 
	.B2(I19[1]), 
	.Z(O9[1])); 
	AN_CELL inst_and_1 ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(O10[1])); 
	AO_CELL inst_0_2 ( 
	.A1(out_sel[0]), 
	.A2(I0[2]), 
	.B1(out_sel[1]), 
	.B2(I1[2]), 
	.Z(O0[2])); 
	AO_CELL inst_1_2 ( 
	.A1(out_sel[2]), 
	.A2(I2[2]), 
	.B1(out_sel[3]), 
	.B2(I3[2]), 
	.Z(O1[2])); 
	AO_CELL inst_2_2 ( 
	.A1(out_sel[4]), 
	.A2(I4[2]), 
	.B1(out_sel[5]), 
	.B2(I5[2]), 
	.Z(O2[2])); 
	AO_CELL inst_3_2 ( 
	.A1(out_sel[6]), 
	.A2(I6[2]), 
	.B1(out_sel[7]), 
	.B2(I7[2]), 
	.Z(O3[2])); 
	AO_CELL inst_4_2 ( 
	.A1(out_sel[8]), 
	.A2(I8[2]), 
	.B1(out_sel[9]), 
	.B2(I9[2]), 
	.Z(O4[2])); 
	AO_CELL inst_5_2 ( 
	.A1(out_sel[10]), 
	.A2(I10[2]), 
	.B1(out_sel[11]), 
	.B2(I11[2]), 
	.Z(O5[2])); 
	AO_CELL inst_6_2 ( 
	.A1(out_sel[12]), 
	.A2(I12[2]), 
	.B1(out_sel[13]), 
	.B2(I13[2]), 
	.Z(O6[2])); 
	AO_CELL inst_7_2 ( 
	.A1(out_sel[14]), 
	.A2(I14[2]), 
	.B1(out_sel[15]), 
	.B2(I15[2]), 
	.Z(O7[2])); 
	AO_CELL inst_8_2 ( 
	.A1(out_sel[16]), 
	.A2(I16[2]), 
	.B1(out_sel[17]), 
	.B2(I17[2]), 
	.Z(O8[2])); 
	AO_CELL inst_9_2 ( 
	.A1(out_sel[18]), 
	.A2(I18[2]), 
	.B1(out_sel[19]), 
	.B2(I19[2]), 
	.Z(O9[2])); 
	AN_CELL inst_and_2 ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(O10[2])); 
	AO_CELL inst_0_3 ( 
	.A1(out_sel[0]), 
	.A2(I0[3]), 
	.B1(out_sel[1]), 
	.B2(I1[3]), 
	.Z(O0[3])); 
	AO_CELL inst_1_3 ( 
	.A1(out_sel[2]), 
	.A2(I2[3]), 
	.B1(out_sel[3]), 
	.B2(I3[3]), 
	.Z(O1[3])); 
	AO_CELL inst_2_3 ( 
	.A1(out_sel[4]), 
	.A2(I4[3]), 
	.B1(out_sel[5]), 
	.B2(I5[3]), 
	.Z(O2[3])); 
	AO_CELL inst_3_3 ( 
	.A1(out_sel[6]), 
	.A2(I6[3]), 
	.B1(out_sel[7]), 
	.B2(I7[3]), 
	.Z(O3[3])); 
	AO_CELL inst_4_3 ( 
	.A1(out_sel[8]), 
	.A2(I8[3]), 
	.B1(out_sel[9]), 
	.B2(I9[3]), 
	.Z(O4[3])); 
	AO_CELL inst_5_3 ( 
	.A1(out_sel[10]), 
	.A2(I10[3]), 
	.B1(out_sel[11]), 
	.B2(I11[3]), 
	.Z(O5[3])); 
	AO_CELL inst_6_3 ( 
	.A1(out_sel[12]), 
	.A2(I12[3]), 
	.B1(out_sel[13]), 
	.B2(I13[3]), 
	.Z(O6[3])); 
	AO_CELL inst_7_3 ( 
	.A1(out_sel[14]), 
	.A2(I14[3]), 
	.B1(out_sel[15]), 
	.B2(I15[3]), 
	.Z(O7[3])); 
	AO_CELL inst_8_3 ( 
	.A1(out_sel[16]), 
	.A2(I16[3]), 
	.B1(out_sel[17]), 
	.B2(I17[3]), 
	.Z(O8[3])); 
	AO_CELL inst_9_3 ( 
	.A1(out_sel[18]), 
	.A2(I18[3]), 
	.B1(out_sel[19]), 
	.B2(I19[3]), 
	.Z(O9[3])); 
	AN_CELL inst_and_3 ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(O10[3])); 
	AO_CELL inst_0_4 ( 
	.A1(out_sel[0]), 
	.A2(I0[4]), 
	.B1(out_sel[1]), 
	.B2(I1[4]), 
	.Z(O0[4])); 
	AO_CELL inst_1_4 ( 
	.A1(out_sel[2]), 
	.A2(I2[4]), 
	.B1(out_sel[3]), 
	.B2(I3[4]), 
	.Z(O1[4])); 
	AO_CELL inst_2_4 ( 
	.A1(out_sel[4]), 
	.A2(I4[4]), 
	.B1(out_sel[5]), 
	.B2(I5[4]), 
	.Z(O2[4])); 
	AO_CELL inst_3_4 ( 
	.A1(out_sel[6]), 
	.A2(I6[4]), 
	.B1(out_sel[7]), 
	.B2(I7[4]), 
	.Z(O3[4])); 
	AO_CELL inst_4_4 ( 
	.A1(out_sel[8]), 
	.A2(I8[4]), 
	.B1(out_sel[9]), 
	.B2(I9[4]), 
	.Z(O4[4])); 
	AO_CELL inst_5_4 ( 
	.A1(out_sel[10]), 
	.A2(I10[4]), 
	.B1(out_sel[11]), 
	.B2(I11[4]), 
	.Z(O5[4])); 
	AO_CELL inst_6_4 ( 
	.A1(out_sel[12]), 
	.A2(I12[4]), 
	.B1(out_sel[13]), 
	.B2(I13[4]), 
	.Z(O6[4])); 
	AO_CELL inst_7_4 ( 
	.A1(out_sel[14]), 
	.A2(I14[4]), 
	.B1(out_sel[15]), 
	.B2(I15[4]), 
	.Z(O7[4])); 
	AO_CELL inst_8_4 ( 
	.A1(out_sel[16]), 
	.A2(I16[4]), 
	.B1(out_sel[17]), 
	.B2(I17[4]), 
	.Z(O8[4])); 
	AO_CELL inst_9_4 ( 
	.A1(out_sel[18]), 
	.A2(I18[4]), 
	.B1(out_sel[19]), 
	.B2(I19[4]), 
	.Z(O9[4])); 
	AN_CELL inst_and_4 ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(O10[4])); 
	AO_CELL inst_0_5 ( 
	.A1(out_sel[0]), 
	.A2(I0[5]), 
	.B1(out_sel[1]), 
	.B2(I1[5]), 
	.Z(O0[5])); 
	AO_CELL inst_1_5 ( 
	.A1(out_sel[2]), 
	.A2(I2[5]), 
	.B1(out_sel[3]), 
	.B2(I3[5]), 
	.Z(O1[5])); 
	AO_CELL inst_2_5 ( 
	.A1(out_sel[4]), 
	.A2(I4[5]), 
	.B1(out_sel[5]), 
	.B2(I5[5]), 
	.Z(O2[5])); 
	AO_CELL inst_3_5 ( 
	.A1(out_sel[6]), 
	.A2(I6[5]), 
	.B1(out_sel[7]), 
	.B2(I7[5]), 
	.Z(O3[5])); 
	AO_CELL inst_4_5 ( 
	.A1(out_sel[8]), 
	.A2(I8[5]), 
	.B1(out_sel[9]), 
	.B2(I9[5]), 
	.Z(O4[5])); 
	AO_CELL inst_5_5 ( 
	.A1(out_sel[10]), 
	.A2(I10[5]), 
	.B1(out_sel[11]), 
	.B2(I11[5]), 
	.Z(O5[5])); 
	AO_CELL inst_6_5 ( 
	.A1(out_sel[12]), 
	.A2(I12[5]), 
	.B1(out_sel[13]), 
	.B2(I13[5]), 
	.Z(O6[5])); 
	AO_CELL inst_7_5 ( 
	.A1(out_sel[14]), 
	.A2(I14[5]), 
	.B1(out_sel[15]), 
	.B2(I15[5]), 
	.Z(O7[5])); 
	AO_CELL inst_8_5 ( 
	.A1(out_sel[16]), 
	.A2(I16[5]), 
	.B1(out_sel[17]), 
	.B2(I17[5]), 
	.Z(O8[5])); 
	AO_CELL inst_9_5 ( 
	.A1(out_sel[18]), 
	.A2(I18[5]), 
	.B1(out_sel[19]), 
	.B2(I19[5]), 
	.Z(O9[5])); 
	AN_CELL inst_and_5 ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(O10[5])); 
	AO_CELL inst_0_6 ( 
	.A1(out_sel[0]), 
	.A2(I0[6]), 
	.B1(out_sel[1]), 
	.B2(I1[6]), 
	.Z(O0[6])); 
	AO_CELL inst_1_6 ( 
	.A1(out_sel[2]), 
	.A2(I2[6]), 
	.B1(out_sel[3]), 
	.B2(I3[6]), 
	.Z(O1[6])); 
	AO_CELL inst_2_6 ( 
	.A1(out_sel[4]), 
	.A2(I4[6]), 
	.B1(out_sel[5]), 
	.B2(I5[6]), 
	.Z(O2[6])); 
	AO_CELL inst_3_6 ( 
	.A1(out_sel[6]), 
	.A2(I6[6]), 
	.B1(out_sel[7]), 
	.B2(I7[6]), 
	.Z(O3[6])); 
	AO_CELL inst_4_6 ( 
	.A1(out_sel[8]), 
	.A2(I8[6]), 
	.B1(out_sel[9]), 
	.B2(I9[6]), 
	.Z(O4[6])); 
	AO_CELL inst_5_6 ( 
	.A1(out_sel[10]), 
	.A2(I10[6]), 
	.B1(out_sel[11]), 
	.B2(I11[6]), 
	.Z(O5[6])); 
	AO_CELL inst_6_6 ( 
	.A1(out_sel[12]), 
	.A2(I12[6]), 
	.B1(out_sel[13]), 
	.B2(I13[6]), 
	.Z(O6[6])); 
	AO_CELL inst_7_6 ( 
	.A1(out_sel[14]), 
	.A2(I14[6]), 
	.B1(out_sel[15]), 
	.B2(I15[6]), 
	.Z(O7[6])); 
	AO_CELL inst_8_6 ( 
	.A1(out_sel[16]), 
	.A2(I16[6]), 
	.B1(out_sel[17]), 
	.B2(I17[6]), 
	.Z(O8[6])); 
	AO_CELL inst_9_6 ( 
	.A1(out_sel[18]), 
	.A2(I18[6]), 
	.B1(out_sel[19]), 
	.B2(I19[6]), 
	.Z(O9[6])); 
	AN_CELL inst_and_6 ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(O10[6])); 
	AO_CELL inst_0_7 ( 
	.A1(out_sel[0]), 
	.A2(I0[7]), 
	.B1(out_sel[1]), 
	.B2(I1[7]), 
	.Z(O0[7])); 
	AO_CELL inst_1_7 ( 
	.A1(out_sel[2]), 
	.A2(I2[7]), 
	.B1(out_sel[3]), 
	.B2(I3[7]), 
	.Z(O1[7])); 
	AO_CELL inst_2_7 ( 
	.A1(out_sel[4]), 
	.A2(I4[7]), 
	.B1(out_sel[5]), 
	.B2(I5[7]), 
	.Z(O2[7])); 
	AO_CELL inst_3_7 ( 
	.A1(out_sel[6]), 
	.A2(I6[7]), 
	.B1(out_sel[7]), 
	.B2(I7[7]), 
	.Z(O3[7])); 
	AO_CELL inst_4_7 ( 
	.A1(out_sel[8]), 
	.A2(I8[7]), 
	.B1(out_sel[9]), 
	.B2(I9[7]), 
	.Z(O4[7])); 
	AO_CELL inst_5_7 ( 
	.A1(out_sel[10]), 
	.A2(I10[7]), 
	.B1(out_sel[11]), 
	.B2(I11[7]), 
	.Z(O5[7])); 
	AO_CELL inst_6_7 ( 
	.A1(out_sel[12]), 
	.A2(I12[7]), 
	.B1(out_sel[13]), 
	.B2(I13[7]), 
	.Z(O6[7])); 
	AO_CELL inst_7_7 ( 
	.A1(out_sel[14]), 
	.A2(I14[7]), 
	.B1(out_sel[15]), 
	.B2(I15[7]), 
	.Z(O7[7])); 
	AO_CELL inst_8_7 ( 
	.A1(out_sel[16]), 
	.A2(I16[7]), 
	.B1(out_sel[17]), 
	.B2(I17[7]), 
	.Z(O8[7])); 
	AO_CELL inst_9_7 ( 
	.A1(out_sel[18]), 
	.A2(I18[7]), 
	.B1(out_sel[19]), 
	.B2(I19[7]), 
	.Z(O9[7])); 
	AN_CELL inst_and_7 ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(O10[7])); 
	AO_CELL inst_0_8 ( 
	.A1(out_sel[0]), 
	.A2(I0[8]), 
	.B1(out_sel[1]), 
	.B2(I1[8]), 
	.Z(O0[8])); 
	AO_CELL inst_1_8 ( 
	.A1(out_sel[2]), 
	.A2(I2[8]), 
	.B1(out_sel[3]), 
	.B2(I3[8]), 
	.Z(O1[8])); 
	AO_CELL inst_2_8 ( 
	.A1(out_sel[4]), 
	.A2(I4[8]), 
	.B1(out_sel[5]), 
	.B2(I5[8]), 
	.Z(O2[8])); 
	AO_CELL inst_3_8 ( 
	.A1(out_sel[6]), 
	.A2(I6[8]), 
	.B1(out_sel[7]), 
	.B2(I7[8]), 
	.Z(O3[8])); 
	AO_CELL inst_4_8 ( 
	.A1(out_sel[8]), 
	.A2(I8[8]), 
	.B1(out_sel[9]), 
	.B2(I9[8]), 
	.Z(O4[8])); 
	AO_CELL inst_5_8 ( 
	.A1(out_sel[10]), 
	.A2(I10[8]), 
	.B1(out_sel[11]), 
	.B2(I11[8]), 
	.Z(O5[8])); 
	AO_CELL inst_6_8 ( 
	.A1(out_sel[12]), 
	.A2(I12[8]), 
	.B1(out_sel[13]), 
	.B2(I13[8]), 
	.Z(O6[8])); 
	AO_CELL inst_7_8 ( 
	.A1(out_sel[14]), 
	.A2(I14[8]), 
	.B1(out_sel[15]), 
	.B2(I15[8]), 
	.Z(O7[8])); 
	AO_CELL inst_8_8 ( 
	.A1(out_sel[16]), 
	.A2(I16[8]), 
	.B1(out_sel[17]), 
	.B2(I17[8]), 
	.Z(O8[8])); 
	AO_CELL inst_9_8 ( 
	.A1(out_sel[18]), 
	.A2(I18[8]), 
	.B1(out_sel[19]), 
	.B2(I19[8]), 
	.Z(O9[8])); 
	AN_CELL inst_and_8 ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(O10[8])); 
	AO_CELL inst_0_9 ( 
	.A1(out_sel[0]), 
	.A2(I0[9]), 
	.B1(out_sel[1]), 
	.B2(I1[9]), 
	.Z(O0[9])); 
	AO_CELL inst_1_9 ( 
	.A1(out_sel[2]), 
	.A2(I2[9]), 
	.B1(out_sel[3]), 
	.B2(I3[9]), 
	.Z(O1[9])); 
	AO_CELL inst_2_9 ( 
	.A1(out_sel[4]), 
	.A2(I4[9]), 
	.B1(out_sel[5]), 
	.B2(I5[9]), 
	.Z(O2[9])); 
	AO_CELL inst_3_9 ( 
	.A1(out_sel[6]), 
	.A2(I6[9]), 
	.B1(out_sel[7]), 
	.B2(I7[9]), 
	.Z(O3[9])); 
	AO_CELL inst_4_9 ( 
	.A1(out_sel[8]), 
	.A2(I8[9]), 
	.B1(out_sel[9]), 
	.B2(I9[9]), 
	.Z(O4[9])); 
	AO_CELL inst_5_9 ( 
	.A1(out_sel[10]), 
	.A2(I10[9]), 
	.B1(out_sel[11]), 
	.B2(I11[9]), 
	.Z(O5[9])); 
	AO_CELL inst_6_9 ( 
	.A1(out_sel[12]), 
	.A2(I12[9]), 
	.B1(out_sel[13]), 
	.B2(I13[9]), 
	.Z(O6[9])); 
	AO_CELL inst_7_9 ( 
	.A1(out_sel[14]), 
	.A2(I14[9]), 
	.B1(out_sel[15]), 
	.B2(I15[9]), 
	.Z(O7[9])); 
	AO_CELL inst_8_9 ( 
	.A1(out_sel[16]), 
	.A2(I16[9]), 
	.B1(out_sel[17]), 
	.B2(I17[9]), 
	.Z(O8[9])); 
	AO_CELL inst_9_9 ( 
	.A1(out_sel[18]), 
	.A2(I18[9]), 
	.B1(out_sel[19]), 
	.B2(I19[9]), 
	.Z(O9[9])); 
	AN_CELL inst_and_9 ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(O10[9])); 
	AO_CELL inst_0_10 ( 
	.A1(out_sel[0]), 
	.A2(I0[10]), 
	.B1(out_sel[1]), 
	.B2(I1[10]), 
	.Z(O0[10])); 
	AO_CELL inst_1_10 ( 
	.A1(out_sel[2]), 
	.A2(I2[10]), 
	.B1(out_sel[3]), 
	.B2(I3[10]), 
	.Z(O1[10])); 
	AO_CELL inst_2_10 ( 
	.A1(out_sel[4]), 
	.A2(I4[10]), 
	.B1(out_sel[5]), 
	.B2(I5[10]), 
	.Z(O2[10])); 
	AO_CELL inst_3_10 ( 
	.A1(out_sel[6]), 
	.A2(I6[10]), 
	.B1(out_sel[7]), 
	.B2(I7[10]), 
	.Z(O3[10])); 
	AO_CELL inst_4_10 ( 
	.A1(out_sel[8]), 
	.A2(I8[10]), 
	.B1(out_sel[9]), 
	.B2(I9[10]), 
	.Z(O4[10])); 
	AO_CELL inst_5_10 ( 
	.A1(out_sel[10]), 
	.A2(I10[10]), 
	.B1(out_sel[11]), 
	.B2(I11[10]), 
	.Z(O5[10])); 
	AO_CELL inst_6_10 ( 
	.A1(out_sel[12]), 
	.A2(I12[10]), 
	.B1(out_sel[13]), 
	.B2(I13[10]), 
	.Z(O6[10])); 
	AO_CELL inst_7_10 ( 
	.A1(out_sel[14]), 
	.A2(I14[10]), 
	.B1(out_sel[15]), 
	.B2(I15[10]), 
	.Z(O7[10])); 
	AO_CELL inst_8_10 ( 
	.A1(out_sel[16]), 
	.A2(I16[10]), 
	.B1(out_sel[17]), 
	.B2(I17[10]), 
	.Z(O8[10])); 
	AO_CELL inst_9_10 ( 
	.A1(out_sel[18]), 
	.A2(I18[10]), 
	.B1(out_sel[19]), 
	.B2(I19[10]), 
	.Z(O9[10])); 
	AN_CELL inst_and_10 ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(O10[10])); 
	AO_CELL inst_0_11 ( 
	.A1(out_sel[0]), 
	.A2(I0[11]), 
	.B1(out_sel[1]), 
	.B2(I1[11]), 
	.Z(O0[11])); 
	AO_CELL inst_1_11 ( 
	.A1(out_sel[2]), 
	.A2(I2[11]), 
	.B1(out_sel[3]), 
	.B2(I3[11]), 
	.Z(O1[11])); 
	AO_CELL inst_2_11 ( 
	.A1(out_sel[4]), 
	.A2(I4[11]), 
	.B1(out_sel[5]), 
	.B2(I5[11]), 
	.Z(O2[11])); 
	AO_CELL inst_3_11 ( 
	.A1(out_sel[6]), 
	.A2(I6[11]), 
	.B1(out_sel[7]), 
	.B2(I7[11]), 
	.Z(O3[11])); 
	AO_CELL inst_4_11 ( 
	.A1(out_sel[8]), 
	.A2(I8[11]), 
	.B1(out_sel[9]), 
	.B2(I9[11]), 
	.Z(O4[11])); 
	AO_CELL inst_5_11 ( 
	.A1(out_sel[10]), 
	.A2(I10[11]), 
	.B1(out_sel[11]), 
	.B2(I11[11]), 
	.Z(O5[11])); 
	AO_CELL inst_6_11 ( 
	.A1(out_sel[12]), 
	.A2(I12[11]), 
	.B1(out_sel[13]), 
	.B2(I13[11]), 
	.Z(O6[11])); 
	AO_CELL inst_7_11 ( 
	.A1(out_sel[14]), 
	.A2(I14[11]), 
	.B1(out_sel[15]), 
	.B2(I15[11]), 
	.Z(O7[11])); 
	AO_CELL inst_8_11 ( 
	.A1(out_sel[16]), 
	.A2(I16[11]), 
	.B1(out_sel[17]), 
	.B2(I17[11]), 
	.Z(O8[11])); 
	AO_CELL inst_9_11 ( 
	.A1(out_sel[18]), 
	.A2(I18[11]), 
	.B1(out_sel[19]), 
	.B2(I19[11]), 
	.Z(O9[11])); 
	AN_CELL inst_and_11 ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(O10[11])); 
	AO_CELL inst_0_12 ( 
	.A1(out_sel[0]), 
	.A2(I0[12]), 
	.B1(out_sel[1]), 
	.B2(I1[12]), 
	.Z(O0[12])); 
	AO_CELL inst_1_12 ( 
	.A1(out_sel[2]), 
	.A2(I2[12]), 
	.B1(out_sel[3]), 
	.B2(I3[12]), 
	.Z(O1[12])); 
	AO_CELL inst_2_12 ( 
	.A1(out_sel[4]), 
	.A2(I4[12]), 
	.B1(out_sel[5]), 
	.B2(I5[12]), 
	.Z(O2[12])); 
	AO_CELL inst_3_12 ( 
	.A1(out_sel[6]), 
	.A2(I6[12]), 
	.B1(out_sel[7]), 
	.B2(I7[12]), 
	.Z(O3[12])); 
	AO_CELL inst_4_12 ( 
	.A1(out_sel[8]), 
	.A2(I8[12]), 
	.B1(out_sel[9]), 
	.B2(I9[12]), 
	.Z(O4[12])); 
	AO_CELL inst_5_12 ( 
	.A1(out_sel[10]), 
	.A2(I10[12]), 
	.B1(out_sel[11]), 
	.B2(I11[12]), 
	.Z(O5[12])); 
	AO_CELL inst_6_12 ( 
	.A1(out_sel[12]), 
	.A2(I12[12]), 
	.B1(out_sel[13]), 
	.B2(I13[12]), 
	.Z(O6[12])); 
	AO_CELL inst_7_12 ( 
	.A1(out_sel[14]), 
	.A2(I14[12]), 
	.B1(out_sel[15]), 
	.B2(I15[12]), 
	.Z(O7[12])); 
	AO_CELL inst_8_12 ( 
	.A1(out_sel[16]), 
	.A2(I16[12]), 
	.B1(out_sel[17]), 
	.B2(I17[12]), 
	.Z(O8[12])); 
	AO_CELL inst_9_12 ( 
	.A1(out_sel[18]), 
	.A2(I18[12]), 
	.B1(out_sel[19]), 
	.B2(I19[12]), 
	.Z(O9[12])); 
	AN_CELL inst_and_12 ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(O10[12])); 
	AO_CELL inst_0_13 ( 
	.A1(out_sel[0]), 
	.A2(I0[13]), 
	.B1(out_sel[1]), 
	.B2(I1[13]), 
	.Z(O0[13])); 
	AO_CELL inst_1_13 ( 
	.A1(out_sel[2]), 
	.A2(I2[13]), 
	.B1(out_sel[3]), 
	.B2(I3[13]), 
	.Z(O1[13])); 
	AO_CELL inst_2_13 ( 
	.A1(out_sel[4]), 
	.A2(I4[13]), 
	.B1(out_sel[5]), 
	.B2(I5[13]), 
	.Z(O2[13])); 
	AO_CELL inst_3_13 ( 
	.A1(out_sel[6]), 
	.A2(I6[13]), 
	.B1(out_sel[7]), 
	.B2(I7[13]), 
	.Z(O3[13])); 
	AO_CELL inst_4_13 ( 
	.A1(out_sel[8]), 
	.A2(I8[13]), 
	.B1(out_sel[9]), 
	.B2(I9[13]), 
	.Z(O4[13])); 
	AO_CELL inst_5_13 ( 
	.A1(out_sel[10]), 
	.A2(I10[13]), 
	.B1(out_sel[11]), 
	.B2(I11[13]), 
	.Z(O5[13])); 
	AO_CELL inst_6_13 ( 
	.A1(out_sel[12]), 
	.A2(I12[13]), 
	.B1(out_sel[13]), 
	.B2(I13[13]), 
	.Z(O6[13])); 
	AO_CELL inst_7_13 ( 
	.A1(out_sel[14]), 
	.A2(I14[13]), 
	.B1(out_sel[15]), 
	.B2(I15[13]), 
	.Z(O7[13])); 
	AO_CELL inst_8_13 ( 
	.A1(out_sel[16]), 
	.A2(I16[13]), 
	.B1(out_sel[17]), 
	.B2(I17[13]), 
	.Z(O8[13])); 
	AO_CELL inst_9_13 ( 
	.A1(out_sel[18]), 
	.A2(I18[13]), 
	.B1(out_sel[19]), 
	.B2(I19[13]), 
	.Z(O9[13])); 
	AN_CELL inst_and_13 ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(O10[13])); 
	AO_CELL inst_0_14 ( 
	.A1(out_sel[0]), 
	.A2(I0[14]), 
	.B1(out_sel[1]), 
	.B2(I1[14]), 
	.Z(O0[14])); 
	AO_CELL inst_1_14 ( 
	.A1(out_sel[2]), 
	.A2(I2[14]), 
	.B1(out_sel[3]), 
	.B2(I3[14]), 
	.Z(O1[14])); 
	AO_CELL inst_2_14 ( 
	.A1(out_sel[4]), 
	.A2(I4[14]), 
	.B1(out_sel[5]), 
	.B2(I5[14]), 
	.Z(O2[14])); 
	AO_CELL inst_3_14 ( 
	.A1(out_sel[6]), 
	.A2(I6[14]), 
	.B1(out_sel[7]), 
	.B2(I7[14]), 
	.Z(O3[14])); 
	AO_CELL inst_4_14 ( 
	.A1(out_sel[8]), 
	.A2(I8[14]), 
	.B1(out_sel[9]), 
	.B2(I9[14]), 
	.Z(O4[14])); 
	AO_CELL inst_5_14 ( 
	.A1(out_sel[10]), 
	.A2(I10[14]), 
	.B1(out_sel[11]), 
	.B2(I11[14]), 
	.Z(O5[14])); 
	AO_CELL inst_6_14 ( 
	.A1(out_sel[12]), 
	.A2(I12[14]), 
	.B1(out_sel[13]), 
	.B2(I13[14]), 
	.Z(O6[14])); 
	AO_CELL inst_7_14 ( 
	.A1(out_sel[14]), 
	.A2(I14[14]), 
	.B1(out_sel[15]), 
	.B2(I15[14]), 
	.Z(O7[14])); 
	AO_CELL inst_8_14 ( 
	.A1(out_sel[16]), 
	.A2(I16[14]), 
	.B1(out_sel[17]), 
	.B2(I17[14]), 
	.Z(O8[14])); 
	AO_CELL inst_9_14 ( 
	.A1(out_sel[18]), 
	.A2(I18[14]), 
	.B1(out_sel[19]), 
	.B2(I19[14]), 
	.Z(O9[14])); 
	AN_CELL inst_and_14 ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(O10[14])); 
	AO_CELL inst_0_15 ( 
	.A1(out_sel[0]), 
	.A2(I0[15]), 
	.B1(out_sel[1]), 
	.B2(I1[15]), 
	.Z(O0[15])); 
	AO_CELL inst_1_15 ( 
	.A1(out_sel[2]), 
	.A2(I2[15]), 
	.B1(out_sel[3]), 
	.B2(I3[15]), 
	.Z(O1[15])); 
	AO_CELL inst_2_15 ( 
	.A1(out_sel[4]), 
	.A2(I4[15]), 
	.B1(out_sel[5]), 
	.B2(I5[15]), 
	.Z(O2[15])); 
	AO_CELL inst_3_15 ( 
	.A1(out_sel[6]), 
	.A2(I6[15]), 
	.B1(out_sel[7]), 
	.B2(I7[15]), 
	.Z(O3[15])); 
	AO_CELL inst_4_15 ( 
	.A1(out_sel[8]), 
	.A2(I8[15]), 
	.B1(out_sel[9]), 
	.B2(I9[15]), 
	.Z(O4[15])); 
	AO_CELL inst_5_15 ( 
	.A1(out_sel[10]), 
	.A2(I10[15]), 
	.B1(out_sel[11]), 
	.B2(I11[15]), 
	.Z(O5[15])); 
	AO_CELL inst_6_15 ( 
	.A1(out_sel[12]), 
	.A2(I12[15]), 
	.B1(out_sel[13]), 
	.B2(I13[15]), 
	.Z(O6[15])); 
	AO_CELL inst_7_15 ( 
	.A1(out_sel[14]), 
	.A2(I14[15]), 
	.B1(out_sel[15]), 
	.B2(I15[15]), 
	.Z(O7[15])); 
	AO_CELL inst_8_15 ( 
	.A1(out_sel[16]), 
	.A2(I16[15]), 
	.B1(out_sel[17]), 
	.B2(I17[15]), 
	.Z(O8[15])); 
	AO_CELL inst_9_15 ( 
	.A1(out_sel[18]), 
	.A2(I18[15]), 
	.B1(out_sel[19]), 
	.B2(I19[15]), 
	.Z(O9[15])); 
	AN_CELL inst_and_15 ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(O10[15])); 
	AO_CELL inst_0_16 ( 
	.A1(out_sel[0]), 
	.A2(I0[16]), 
	.B1(out_sel[1]), 
	.B2(I1[16]), 
	.Z(O0[16])); 
	AO_CELL inst_1_16 ( 
	.A1(out_sel[2]), 
	.A2(I2[16]), 
	.B1(out_sel[3]), 
	.B2(I3[16]), 
	.Z(O1[16])); 
	AO_CELL inst_2_16 ( 
	.A1(out_sel[4]), 
	.A2(I4[16]), 
	.B1(out_sel[5]), 
	.B2(I5[16]), 
	.Z(O2[16])); 
	AO_CELL inst_3_16 ( 
	.A1(out_sel[6]), 
	.A2(I6[16]), 
	.B1(out_sel[7]), 
	.B2(I7[16]), 
	.Z(O3[16])); 
	AO_CELL inst_4_16 ( 
	.A1(out_sel[8]), 
	.A2(I8[16]), 
	.B1(out_sel[9]), 
	.B2(I9[16]), 
	.Z(O4[16])); 
	AO_CELL inst_5_16 ( 
	.A1(out_sel[10]), 
	.A2(I10[16]), 
	.B1(out_sel[11]), 
	.B2(I11[16]), 
	.Z(O5[16])); 
	AO_CELL inst_6_16 ( 
	.A1(out_sel[12]), 
	.A2(I12[16]), 
	.B1(out_sel[13]), 
	.B2(I13[16]), 
	.Z(O6[16])); 
	AO_CELL inst_7_16 ( 
	.A1(out_sel[14]), 
	.A2(I14[16]), 
	.B1(out_sel[15]), 
	.B2(I15[16]), 
	.Z(O7[16])); 
	AO_CELL inst_8_16 ( 
	.A1(out_sel[16]), 
	.A2(I16[16]), 
	.B1(out_sel[17]), 
	.B2(I17[16]), 
	.Z(O8[16])); 
	AO_CELL inst_9_16 ( 
	.A1(out_sel[18]), 
	.A2(I18[16]), 
	.B1(out_sel[19]), 
	.B2(I19[16]), 
	.Z(O9[16])); 
	AN_CELL inst_and_16 ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(O10[16])); 
	AO_CELL inst_0_valid ( 
	.A1(out_sel[0]), 
	.A2(valid_in[0]), 
	.B1(out_sel[1]), 
	.B2(valid_in[1]), 
	.Z(valid_out[0])); 
	AO_CELL inst_1_valid ( 
	.A1(out_sel[2]), 
	.A2(valid_in[2]), 
	.B1(out_sel[3]), 
	.B2(valid_in[3]), 
	.Z(valid_out[1])); 
	AO_CELL inst_2_valid ( 
	.A1(out_sel[4]), 
	.A2(valid_in[4]), 
	.B1(out_sel[5]), 
	.B2(valid_in[5]), 
	.Z(valid_out[2])); 
	AO_CELL inst_3_valid ( 
	.A1(out_sel[6]), 
	.A2(valid_in[6]), 
	.B1(out_sel[7]), 
	.B2(valid_in[7]), 
	.Z(valid_out[3])); 
	AO_CELL inst_4_valid ( 
	.A1(out_sel[8]), 
	.A2(valid_in[8]), 
	.B1(out_sel[9]), 
	.B2(valid_in[9]), 
	.Z(valid_out[4])); 
	AO_CELL inst_5_valid ( 
	.A1(out_sel[10]), 
	.A2(valid_in[10]), 
	.B1(out_sel[11]), 
	.B2(valid_in[11]), 
	.Z(valid_out[5])); 
	AO_CELL inst_6_valid ( 
	.A1(out_sel[12]), 
	.A2(valid_in[12]), 
	.B1(out_sel[13]), 
	.B2(valid_in[13]), 
	.Z(valid_out[6])); 
	AO_CELL inst_7_valid ( 
	.A1(out_sel[14]), 
	.A2(valid_in[14]), 
	.B1(out_sel[15]), 
	.B2(valid_in[15]), 
	.Z(valid_out[7])); 
	AO_CELL inst_8_valid ( 
	.A1(out_sel[16]), 
	.A2(valid_in[16]), 
	.B1(out_sel[17]), 
	.B2(valid_in[17]), 
	.Z(valid_out[8])); 
	AO_CELL inst_9_valid ( 
	.A1(out_sel[18]), 
	.A2(valid_in[18]), 
	.B1(out_sel[19]), 
	.B2(valid_in[19]), 
	.Z(valid_out[9])); 
	AN_CELL inst_and_10_valid ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(valid_out[10])); 
endmodule 

module mux_aoi_ready_valid_const_20_1 ( 
	input logic  [0 : 0] I[19:0], 
	input logic  [4 : 0] S ,
	input logic ready_in,
	output logic ready_out,
	input logic [19:0]  valid_in,
	output logic valid_out,
	output logic  [31 : 0] out_sel,
	output logic [0 : 0] O); 
	logic  [0 : 0] O_int0;
	logic  [0 : 0] O_int1;
	logic  [0 : 0] O_int2;
	logic  [0 : 0] O_int3;
	logic  [0 : 0] O_int4;
	logic  [0 : 0] O_int5;
	logic  [0 : 0] O_int6;
	logic  [0 : 0] O_int7;
	logic  [0 : 0] O_int8;
	logic  [0 : 0] O_int9;
	logic  [0 : 0] O_int10;
	logic [10:0] valid_out_temp;

precoder_1_20 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_1_20 u_mux_logic ( 
	.I0 (I[0]),
	.I1 (I[1]),
	.I2 (I[2]),
	.I3 (I[3]),
	.I4 (I[4]),
	.I5 (I[5]),
	.I6 (I[6]),
	.I7 (I[7]),
	.I8 (I[8]),
	.I9 (I[9]),
	.I10 (I[10]),
	.I11 (I[11]),
	.I12 (I[12]),
	.I13 (I[13]),
	.I14 (I[14]),
	.I15 (I[15]),
	.I16 (I[16]),
	.I17 (I[17]),
	.I18 (I[18]),
	.I19 (I[19]),
	.out_sel(out_sel), 
	.valid_in(valid_in),
	.valid_out(valid_out_temp),
	.O0(O_int0), 
	.O1(O_int1), 
	.O2(O_int2), 
	.O3(O_int3), 
	.O4(O_int4), 
	.O5(O_int5), 
	.O6(O_int6), 
	.O7(O_int7), 
	.O8(O_int8), 
	.O9(O_int9), 
	.O10(O_int10)); 
	assign O = (  	O_int0 | 	O_int1 | 	O_int2 | 	O_int3 | 	O_int4 | 	O_int5 | 	O_int6 | 	O_int7 | 	O_int8 | 	O_int9 | 	O_int10 	); 
	assign ready_out = ready_in;
	assign valid_out = |valid_out_temp;

endmodule 

module precoder_1_20 (
	input logic  [4 : 0] S ,
	output logic  [31 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		5'd0    :   out_sel = 32'b00000000000000000000000000000001;
		5'd1    :   out_sel = 32'b00000000000000000000000000000010;
		5'd2    :   out_sel = 32'b00000000000000000000000000000100;
		5'd3    :   out_sel = 32'b00000000000000000000000000001000;
		5'd4    :   out_sel = 32'b00000000000000000000000000010000;
		5'd5    :   out_sel = 32'b00000000000000000000000000100000;
		5'd6    :   out_sel = 32'b00000000000000000000000001000000;
		5'd7    :   out_sel = 32'b00000000000000000000000010000000;
		5'd8    :   out_sel = 32'b00000000000000000000000100000000;
		5'd9    :   out_sel = 32'b00000000000000000000001000000000;
		5'd10    :   out_sel = 32'b00000000000000000000010000000000;
		5'd11    :   out_sel = 32'b00000000000000000000100000000000;
		5'd12    :   out_sel = 32'b00000000000000000001000000000000;
		5'd13    :   out_sel = 32'b00000000000000000010000000000000;
		5'd14    :   out_sel = 32'b00000000000000000100000000000000;
		5'd15    :   out_sel = 32'b00000000000000001000000000000000;
		5'd16    :   out_sel = 32'b00000000000000010000000000000000;
		5'd17    :   out_sel = 32'b00000000000000100000000000000000;
		5'd18    :   out_sel = 32'b00000000000001000000000000000000;
		5'd19    :   out_sel = 32'b00000000000010000000000000000000;
		5'd20    :   out_sel = 32'b00000000000100000000000000000000;
		default :   out_sel = 32'b0;
	endcase 
end 

endmodule 

module mux_logic_1_20 ( 
	input logic  [31 : 0] out_sel,
	input logic  [0 : 0] I0, 
	input logic  [0 : 0] I1, 
	input logic  [0 : 0] I2, 
	input logic  [0 : 0] I3, 
	input logic  [0 : 0] I4, 
	input logic  [0 : 0] I5, 
	input logic  [0 : 0] I6, 
	input logic  [0 : 0] I7, 
	input logic  [0 : 0] I8, 
	input logic  [0 : 0] I9, 
	input logic  [0 : 0] I10, 
	input logic  [0 : 0] I11, 
	input logic  [0 : 0] I12, 
	input logic  [0 : 0] I13, 
	input logic  [0 : 0] I14, 
	input logic  [0 : 0] I15, 
	input logic  [0 : 0] I16, 
	input logic  [0 : 0] I17, 
	input logic  [0 : 0] I18, 
	input logic  [0 : 0] I19, 
	input logic [19:0] valid_in,
	output logic [10:0] valid_out,
	output logic  [0 : 0] O0, 
	output logic  [0 : 0] O1, 
	output logic  [0 : 0] O2, 
	output logic  [0 : 0] O3, 
	output logic  [0 : 0] O4, 
	output logic  [0 : 0] O5, 
	output logic  [0 : 0] O6, 
	output logic  [0 : 0] O7, 
	output logic  [0 : 0] O8, 
	output logic  [0 : 0] O9, 
	output logic  [0 : 0] O10); 
	AO_CELL inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	AO_CELL inst_1_0 ( 
	.A1(out_sel[2]), 
	.A2(I2[0]), 
	.B1(out_sel[3]), 
	.B2(I3[0]), 
	.Z(O1[0])); 
	AO_CELL inst_2_0 ( 
	.A1(out_sel[4]), 
	.A2(I4[0]), 
	.B1(out_sel[5]), 
	.B2(I5[0]), 
	.Z(O2[0])); 
	AO_CELL inst_3_0 ( 
	.A1(out_sel[6]), 
	.A2(I6[0]), 
	.B1(out_sel[7]), 
	.B2(I7[0]), 
	.Z(O3[0])); 
	AO_CELL inst_4_0 ( 
	.A1(out_sel[8]), 
	.A2(I8[0]), 
	.B1(out_sel[9]), 
	.B2(I9[0]), 
	.Z(O4[0])); 
	AO_CELL inst_5_0 ( 
	.A1(out_sel[10]), 
	.A2(I10[0]), 
	.B1(out_sel[11]), 
	.B2(I11[0]), 
	.Z(O5[0])); 
	AO_CELL inst_6_0 ( 
	.A1(out_sel[12]), 
	.A2(I12[0]), 
	.B1(out_sel[13]), 
	.B2(I13[0]), 
	.Z(O6[0])); 
	AO_CELL inst_7_0 ( 
	.A1(out_sel[14]), 
	.A2(I14[0]), 
	.B1(out_sel[15]), 
	.B2(I15[0]), 
	.Z(O7[0])); 
	AO_CELL inst_8_0 ( 
	.A1(out_sel[16]), 
	.A2(I16[0]), 
	.B1(out_sel[17]), 
	.B2(I17[0]), 
	.Z(O8[0])); 
	AO_CELL inst_9_0 ( 
	.A1(out_sel[18]), 
	.A2(I18[0]), 
	.B1(out_sel[19]), 
	.B2(I19[0]), 
	.Z(O9[0])); 
	AN_CELL inst_and_0 ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(O10[0])); 
	AO_CELL inst_0_valid ( 
	.A1(out_sel[0]), 
	.A2(valid_in[0]), 
	.B1(out_sel[1]), 
	.B2(valid_in[1]), 
	.Z(valid_out[0])); 
	AO_CELL inst_1_valid ( 
	.A1(out_sel[2]), 
	.A2(valid_in[2]), 
	.B1(out_sel[3]), 
	.B2(valid_in[3]), 
	.Z(valid_out[1])); 
	AO_CELL inst_2_valid ( 
	.A1(out_sel[4]), 
	.A2(valid_in[4]), 
	.B1(out_sel[5]), 
	.B2(valid_in[5]), 
	.Z(valid_out[2])); 
	AO_CELL inst_3_valid ( 
	.A1(out_sel[6]), 
	.A2(valid_in[6]), 
	.B1(out_sel[7]), 
	.B2(valid_in[7]), 
	.Z(valid_out[3])); 
	AO_CELL inst_4_valid ( 
	.A1(out_sel[8]), 
	.A2(valid_in[8]), 
	.B1(out_sel[9]), 
	.B2(valid_in[9]), 
	.Z(valid_out[4])); 
	AO_CELL inst_5_valid ( 
	.A1(out_sel[10]), 
	.A2(valid_in[10]), 
	.B1(out_sel[11]), 
	.B2(valid_in[11]), 
	.Z(valid_out[5])); 
	AO_CELL inst_6_valid ( 
	.A1(out_sel[12]), 
	.A2(valid_in[12]), 
	.B1(out_sel[13]), 
	.B2(valid_in[13]), 
	.Z(valid_out[6])); 
	AO_CELL inst_7_valid ( 
	.A1(out_sel[14]), 
	.A2(valid_in[14]), 
	.B1(out_sel[15]), 
	.B2(valid_in[15]), 
	.Z(valid_out[7])); 
	AO_CELL inst_8_valid ( 
	.A1(out_sel[16]), 
	.A2(valid_in[16]), 
	.B1(out_sel[17]), 
	.B2(valid_in[17]), 
	.Z(valid_out[8])); 
	AO_CELL inst_9_valid ( 
	.A1(out_sel[18]), 
	.A2(valid_in[18]), 
	.B1(out_sel[19]), 
	.B2(valid_in[19]), 
	.Z(valid_out[9])); 
	AN_CELL inst_and_10_valid ( 
	.A1(out_sel[20]), 
	.A2(1'b0), 
	.Z(valid_out[10])); 
endmodule 

module mux_aoi_ready_valid_7_17 ( 
	input logic  [16 : 0] I[6:0], 
	input logic  [2 : 0] S ,
	input logic ready_in,
	output logic ready_out,
	input logic [6:0]  valid_in,
	output logic valid_out,
	output logic  [7 : 0] out_sel,
	output logic [16 : 0] O); 
	logic  [16 : 0] O_int0;
	logic  [16 : 0] O_int1;
	logic  [16 : 0] O_int2;
	logic  [16 : 0] O_int3;
	logic [3:0] valid_out_temp;

precoder_17_7 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_17_7 u_mux_logic ( 
	.I0 (I[0]),
	.I1 (I[1]),
	.I2 (I[2]),
	.I3 (I[3]),
	.I4 (I[4]),
	.I5 (I[5]),
	.I6 (I[6]),
	.out_sel(out_sel), 
	.valid_in(valid_in),
	.valid_out(valid_out_temp),
	.O0(O_int0), 
	.O1(O_int1), 
	.O2(O_int2), 
	.O3(O_int3)); 
	assign O = (  	O_int0 | 	O_int1 | 	O_int2 | 	O_int3 	); 
	assign ready_out = ready_in;
	assign valid_out = |valid_out_temp;

endmodule 

module precoder_17_7 (
	input logic  [2 : 0] S ,
	output logic  [7 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		3'd0    :   out_sel = 8'b00000001;
		3'd1    :   out_sel = 8'b00000010;
		3'd2    :   out_sel = 8'b00000100;
		3'd3    :   out_sel = 8'b00001000;
		3'd4    :   out_sel = 8'b00010000;
		3'd5    :   out_sel = 8'b00100000;
		3'd6    :   out_sel = 8'b01000000;
		default :   out_sel = 8'b0;
	endcase 
end 

endmodule 

module mux_logic_17_7 ( 
	input logic  [7 : 0] out_sel,
	input logic  [16 : 0] I0, 
	input logic  [16 : 0] I1, 
	input logic  [16 : 0] I2, 
	input logic  [16 : 0] I3, 
	input logic  [16 : 0] I4, 
	input logic  [16 : 0] I5, 
	input logic  [16 : 0] I6, 
	input logic [6:0] valid_in,
	output logic [3:0] valid_out,
	output logic  [16 : 0] O0, 
	output logic  [16 : 0] O1, 
	output logic  [16 : 0] O2, 
	output logic  [16 : 0] O3); 
	AO_CELL inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	AO_CELL inst_1_0 ( 
	.A1(out_sel[2]), 
	.A2(I2[0]), 
	.B1(out_sel[3]), 
	.B2(I3[0]), 
	.Z(O1[0])); 
	AO_CELL inst_2_0 ( 
	.A1(out_sel[4]), 
	.A2(I4[0]), 
	.B1(out_sel[5]), 
	.B2(I5[0]), 
	.Z(O2[0])); 
	AN_CELL inst_and_0 ( 
	.A1(out_sel[6]), 
	.A2(I6[0]), 
	.Z(O3[0])); 
	AO_CELL inst_0_1 ( 
	.A1(out_sel[0]), 
	.A2(I0[1]), 
	.B1(out_sel[1]), 
	.B2(I1[1]), 
	.Z(O0[1])); 
	AO_CELL inst_1_1 ( 
	.A1(out_sel[2]), 
	.A2(I2[1]), 
	.B1(out_sel[3]), 
	.B2(I3[1]), 
	.Z(O1[1])); 
	AO_CELL inst_2_1 ( 
	.A1(out_sel[4]), 
	.A2(I4[1]), 
	.B1(out_sel[5]), 
	.B2(I5[1]), 
	.Z(O2[1])); 
	AN_CELL inst_and_1 ( 
	.A1(out_sel[6]), 
	.A2(I6[1]), 
	.Z(O3[1])); 
	AO_CELL inst_0_2 ( 
	.A1(out_sel[0]), 
	.A2(I0[2]), 
	.B1(out_sel[1]), 
	.B2(I1[2]), 
	.Z(O0[2])); 
	AO_CELL inst_1_2 ( 
	.A1(out_sel[2]), 
	.A2(I2[2]), 
	.B1(out_sel[3]), 
	.B2(I3[2]), 
	.Z(O1[2])); 
	AO_CELL inst_2_2 ( 
	.A1(out_sel[4]), 
	.A2(I4[2]), 
	.B1(out_sel[5]), 
	.B2(I5[2]), 
	.Z(O2[2])); 
	AN_CELL inst_and_2 ( 
	.A1(out_sel[6]), 
	.A2(I6[2]), 
	.Z(O3[2])); 
	AO_CELL inst_0_3 ( 
	.A1(out_sel[0]), 
	.A2(I0[3]), 
	.B1(out_sel[1]), 
	.B2(I1[3]), 
	.Z(O0[3])); 
	AO_CELL inst_1_3 ( 
	.A1(out_sel[2]), 
	.A2(I2[3]), 
	.B1(out_sel[3]), 
	.B2(I3[3]), 
	.Z(O1[3])); 
	AO_CELL inst_2_3 ( 
	.A1(out_sel[4]), 
	.A2(I4[3]), 
	.B1(out_sel[5]), 
	.B2(I5[3]), 
	.Z(O2[3])); 
	AN_CELL inst_and_3 ( 
	.A1(out_sel[6]), 
	.A2(I6[3]), 
	.Z(O3[3])); 
	AO_CELL inst_0_4 ( 
	.A1(out_sel[0]), 
	.A2(I0[4]), 
	.B1(out_sel[1]), 
	.B2(I1[4]), 
	.Z(O0[4])); 
	AO_CELL inst_1_4 ( 
	.A1(out_sel[2]), 
	.A2(I2[4]), 
	.B1(out_sel[3]), 
	.B2(I3[4]), 
	.Z(O1[4])); 
	AO_CELL inst_2_4 ( 
	.A1(out_sel[4]), 
	.A2(I4[4]), 
	.B1(out_sel[5]), 
	.B2(I5[4]), 
	.Z(O2[4])); 
	AN_CELL inst_and_4 ( 
	.A1(out_sel[6]), 
	.A2(I6[4]), 
	.Z(O3[4])); 
	AO_CELL inst_0_5 ( 
	.A1(out_sel[0]), 
	.A2(I0[5]), 
	.B1(out_sel[1]), 
	.B2(I1[5]), 
	.Z(O0[5])); 
	AO_CELL inst_1_5 ( 
	.A1(out_sel[2]), 
	.A2(I2[5]), 
	.B1(out_sel[3]), 
	.B2(I3[5]), 
	.Z(O1[5])); 
	AO_CELL inst_2_5 ( 
	.A1(out_sel[4]), 
	.A2(I4[5]), 
	.B1(out_sel[5]), 
	.B2(I5[5]), 
	.Z(O2[5])); 
	AN_CELL inst_and_5 ( 
	.A1(out_sel[6]), 
	.A2(I6[5]), 
	.Z(O3[5])); 
	AO_CELL inst_0_6 ( 
	.A1(out_sel[0]), 
	.A2(I0[6]), 
	.B1(out_sel[1]), 
	.B2(I1[6]), 
	.Z(O0[6])); 
	AO_CELL inst_1_6 ( 
	.A1(out_sel[2]), 
	.A2(I2[6]), 
	.B1(out_sel[3]), 
	.B2(I3[6]), 
	.Z(O1[6])); 
	AO_CELL inst_2_6 ( 
	.A1(out_sel[4]), 
	.A2(I4[6]), 
	.B1(out_sel[5]), 
	.B2(I5[6]), 
	.Z(O2[6])); 
	AN_CELL inst_and_6 ( 
	.A1(out_sel[6]), 
	.A2(I6[6]), 
	.Z(O3[6])); 
	AO_CELL inst_0_7 ( 
	.A1(out_sel[0]), 
	.A2(I0[7]), 
	.B1(out_sel[1]), 
	.B2(I1[7]), 
	.Z(O0[7])); 
	AO_CELL inst_1_7 ( 
	.A1(out_sel[2]), 
	.A2(I2[7]), 
	.B1(out_sel[3]), 
	.B2(I3[7]), 
	.Z(O1[7])); 
	AO_CELL inst_2_7 ( 
	.A1(out_sel[4]), 
	.A2(I4[7]), 
	.B1(out_sel[5]), 
	.B2(I5[7]), 
	.Z(O2[7])); 
	AN_CELL inst_and_7 ( 
	.A1(out_sel[6]), 
	.A2(I6[7]), 
	.Z(O3[7])); 
	AO_CELL inst_0_8 ( 
	.A1(out_sel[0]), 
	.A2(I0[8]), 
	.B1(out_sel[1]), 
	.B2(I1[8]), 
	.Z(O0[8])); 
	AO_CELL inst_1_8 ( 
	.A1(out_sel[2]), 
	.A2(I2[8]), 
	.B1(out_sel[3]), 
	.B2(I3[8]), 
	.Z(O1[8])); 
	AO_CELL inst_2_8 ( 
	.A1(out_sel[4]), 
	.A2(I4[8]), 
	.B1(out_sel[5]), 
	.B2(I5[8]), 
	.Z(O2[8])); 
	AN_CELL inst_and_8 ( 
	.A1(out_sel[6]), 
	.A2(I6[8]), 
	.Z(O3[8])); 
	AO_CELL inst_0_9 ( 
	.A1(out_sel[0]), 
	.A2(I0[9]), 
	.B1(out_sel[1]), 
	.B2(I1[9]), 
	.Z(O0[9])); 
	AO_CELL inst_1_9 ( 
	.A1(out_sel[2]), 
	.A2(I2[9]), 
	.B1(out_sel[3]), 
	.B2(I3[9]), 
	.Z(O1[9])); 
	AO_CELL inst_2_9 ( 
	.A1(out_sel[4]), 
	.A2(I4[9]), 
	.B1(out_sel[5]), 
	.B2(I5[9]), 
	.Z(O2[9])); 
	AN_CELL inst_and_9 ( 
	.A1(out_sel[6]), 
	.A2(I6[9]), 
	.Z(O3[9])); 
	AO_CELL inst_0_10 ( 
	.A1(out_sel[0]), 
	.A2(I0[10]), 
	.B1(out_sel[1]), 
	.B2(I1[10]), 
	.Z(O0[10])); 
	AO_CELL inst_1_10 ( 
	.A1(out_sel[2]), 
	.A2(I2[10]), 
	.B1(out_sel[3]), 
	.B2(I3[10]), 
	.Z(O1[10])); 
	AO_CELL inst_2_10 ( 
	.A1(out_sel[4]), 
	.A2(I4[10]), 
	.B1(out_sel[5]), 
	.B2(I5[10]), 
	.Z(O2[10])); 
	AN_CELL inst_and_10 ( 
	.A1(out_sel[6]), 
	.A2(I6[10]), 
	.Z(O3[10])); 
	AO_CELL inst_0_11 ( 
	.A1(out_sel[0]), 
	.A2(I0[11]), 
	.B1(out_sel[1]), 
	.B2(I1[11]), 
	.Z(O0[11])); 
	AO_CELL inst_1_11 ( 
	.A1(out_sel[2]), 
	.A2(I2[11]), 
	.B1(out_sel[3]), 
	.B2(I3[11]), 
	.Z(O1[11])); 
	AO_CELL inst_2_11 ( 
	.A1(out_sel[4]), 
	.A2(I4[11]), 
	.B1(out_sel[5]), 
	.B2(I5[11]), 
	.Z(O2[11])); 
	AN_CELL inst_and_11 ( 
	.A1(out_sel[6]), 
	.A2(I6[11]), 
	.Z(O3[11])); 
	AO_CELL inst_0_12 ( 
	.A1(out_sel[0]), 
	.A2(I0[12]), 
	.B1(out_sel[1]), 
	.B2(I1[12]), 
	.Z(O0[12])); 
	AO_CELL inst_1_12 ( 
	.A1(out_sel[2]), 
	.A2(I2[12]), 
	.B1(out_sel[3]), 
	.B2(I3[12]), 
	.Z(O1[12])); 
	AO_CELL inst_2_12 ( 
	.A1(out_sel[4]), 
	.A2(I4[12]), 
	.B1(out_sel[5]), 
	.B2(I5[12]), 
	.Z(O2[12])); 
	AN_CELL inst_and_12 ( 
	.A1(out_sel[6]), 
	.A2(I6[12]), 
	.Z(O3[12])); 
	AO_CELL inst_0_13 ( 
	.A1(out_sel[0]), 
	.A2(I0[13]), 
	.B1(out_sel[1]), 
	.B2(I1[13]), 
	.Z(O0[13])); 
	AO_CELL inst_1_13 ( 
	.A1(out_sel[2]), 
	.A2(I2[13]), 
	.B1(out_sel[3]), 
	.B2(I3[13]), 
	.Z(O1[13])); 
	AO_CELL inst_2_13 ( 
	.A1(out_sel[4]), 
	.A2(I4[13]), 
	.B1(out_sel[5]), 
	.B2(I5[13]), 
	.Z(O2[13])); 
	AN_CELL inst_and_13 ( 
	.A1(out_sel[6]), 
	.A2(I6[13]), 
	.Z(O3[13])); 
	AO_CELL inst_0_14 ( 
	.A1(out_sel[0]), 
	.A2(I0[14]), 
	.B1(out_sel[1]), 
	.B2(I1[14]), 
	.Z(O0[14])); 
	AO_CELL inst_1_14 ( 
	.A1(out_sel[2]), 
	.A2(I2[14]), 
	.B1(out_sel[3]), 
	.B2(I3[14]), 
	.Z(O1[14])); 
	AO_CELL inst_2_14 ( 
	.A1(out_sel[4]), 
	.A2(I4[14]), 
	.B1(out_sel[5]), 
	.B2(I5[14]), 
	.Z(O2[14])); 
	AN_CELL inst_and_14 ( 
	.A1(out_sel[6]), 
	.A2(I6[14]), 
	.Z(O3[14])); 
	AO_CELL inst_0_15 ( 
	.A1(out_sel[0]), 
	.A2(I0[15]), 
	.B1(out_sel[1]), 
	.B2(I1[15]), 
	.Z(O0[15])); 
	AO_CELL inst_1_15 ( 
	.A1(out_sel[2]), 
	.A2(I2[15]), 
	.B1(out_sel[3]), 
	.B2(I3[15]), 
	.Z(O1[15])); 
	AO_CELL inst_2_15 ( 
	.A1(out_sel[4]), 
	.A2(I4[15]), 
	.B1(out_sel[5]), 
	.B2(I5[15]), 
	.Z(O2[15])); 
	AN_CELL inst_and_15 ( 
	.A1(out_sel[6]), 
	.A2(I6[15]), 
	.Z(O3[15])); 
	AO_CELL inst_0_16 ( 
	.A1(out_sel[0]), 
	.A2(I0[16]), 
	.B1(out_sel[1]), 
	.B2(I1[16]), 
	.Z(O0[16])); 
	AO_CELL inst_1_16 ( 
	.A1(out_sel[2]), 
	.A2(I2[16]), 
	.B1(out_sel[3]), 
	.B2(I3[16]), 
	.Z(O1[16])); 
	AO_CELL inst_2_16 ( 
	.A1(out_sel[4]), 
	.A2(I4[16]), 
	.B1(out_sel[5]), 
	.B2(I5[16]), 
	.Z(O2[16])); 
	AN_CELL inst_and_16 ( 
	.A1(out_sel[6]), 
	.A2(I6[16]), 
	.Z(O3[16])); 
	AO_CELL inst_0_valid ( 
	.A1(out_sel[0]), 
	.A2(valid_in[0]), 
	.B1(out_sel[1]), 
	.B2(valid_in[1]), 
	.Z(valid_out[0])); 
	AO_CELL inst_1_valid ( 
	.A1(out_sel[2]), 
	.A2(valid_in[2]), 
	.B1(out_sel[3]), 
	.B2(valid_in[3]), 
	.Z(valid_out[1])); 
	AO_CELL inst_2_valid ( 
	.A1(out_sel[4]), 
	.A2(valid_in[4]), 
	.B1(out_sel[5]), 
	.B2(valid_in[5]), 
	.Z(valid_out[2])); 
	AN_CELL inst_and_3_valid ( 
	.A1(out_sel[6]), 
	.A2(valid_in[6]), 
	.Z(valid_out[3])); 
endmodule 

module mux_aoi_ready_valid_6_17 ( 
	input logic  [16 : 0] I[5:0], 
	input logic  [2 : 0] S ,
	input logic ready_in,
	output logic ready_out,
	input logic [5:0]  valid_in,
	output logic valid_out,
	output logic  [7 : 0] out_sel,
	output logic [16 : 0] O); 
	logic  [16 : 0] O_int0;
	logic  [16 : 0] O_int1;
	logic  [16 : 0] O_int2;
	logic [2:0] valid_out_temp;

precoder_17_6 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_17_6 u_mux_logic ( 
	.I0 (I[0]),
	.I1 (I[1]),
	.I2 (I[2]),
	.I3 (I[3]),
	.I4 (I[4]),
	.I5 (I[5]),
	.out_sel(out_sel), 
	.valid_in(valid_in),
	.valid_out(valid_out_temp),
	.O0(O_int0), 
	.O1(O_int1), 
	.O2(O_int2)); 
	assign O = (  	O_int0 | 	O_int1 | 	O_int2 	); 
	assign ready_out = ready_in;
	assign valid_out = |valid_out_temp;

endmodule 

module precoder_17_6 (
	input logic  [2 : 0] S ,
	output logic  [7 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		3'd0    :   out_sel = 8'b00000001;
		3'd1    :   out_sel = 8'b00000010;
		3'd2    :   out_sel = 8'b00000100;
		3'd3    :   out_sel = 8'b00001000;
		3'd4    :   out_sel = 8'b00010000;
		3'd5    :   out_sel = 8'b00100000;
		default :   out_sel = 8'b0;
	endcase 
end 

endmodule 

module mux_logic_17_6 ( 
	input logic  [7 : 0] out_sel,
	input logic  [16 : 0] I0, 
	input logic  [16 : 0] I1, 
	input logic  [16 : 0] I2, 
	input logic  [16 : 0] I3, 
	input logic  [16 : 0] I4, 
	input logic  [16 : 0] I5, 
	input logic [5:0] valid_in,
	output logic [2:0] valid_out,
	output logic  [16 : 0] O0, 
	output logic  [16 : 0] O1, 
	output logic  [16 : 0] O2); 
	AO_CELL inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	AO_CELL inst_1_0 ( 
	.A1(out_sel[2]), 
	.A2(I2[0]), 
	.B1(out_sel[3]), 
	.B2(I3[0]), 
	.Z(O1[0])); 
	AO_CELL inst_2_0 ( 
	.A1(out_sel[4]), 
	.A2(I4[0]), 
	.B1(out_sel[5]), 
	.B2(I5[0]), 
	.Z(O2[0])); 
	AO_CELL inst_0_1 ( 
	.A1(out_sel[0]), 
	.A2(I0[1]), 
	.B1(out_sel[1]), 
	.B2(I1[1]), 
	.Z(O0[1])); 
	AO_CELL inst_1_1 ( 
	.A1(out_sel[2]), 
	.A2(I2[1]), 
	.B1(out_sel[3]), 
	.B2(I3[1]), 
	.Z(O1[1])); 
	AO_CELL inst_2_1 ( 
	.A1(out_sel[4]), 
	.A2(I4[1]), 
	.B1(out_sel[5]), 
	.B2(I5[1]), 
	.Z(O2[1])); 
	AO_CELL inst_0_2 ( 
	.A1(out_sel[0]), 
	.A2(I0[2]), 
	.B1(out_sel[1]), 
	.B2(I1[2]), 
	.Z(O0[2])); 
	AO_CELL inst_1_2 ( 
	.A1(out_sel[2]), 
	.A2(I2[2]), 
	.B1(out_sel[3]), 
	.B2(I3[2]), 
	.Z(O1[2])); 
	AO_CELL inst_2_2 ( 
	.A1(out_sel[4]), 
	.A2(I4[2]), 
	.B1(out_sel[5]), 
	.B2(I5[2]), 
	.Z(O2[2])); 
	AO_CELL inst_0_3 ( 
	.A1(out_sel[0]), 
	.A2(I0[3]), 
	.B1(out_sel[1]), 
	.B2(I1[3]), 
	.Z(O0[3])); 
	AO_CELL inst_1_3 ( 
	.A1(out_sel[2]), 
	.A2(I2[3]), 
	.B1(out_sel[3]), 
	.B2(I3[3]), 
	.Z(O1[3])); 
	AO_CELL inst_2_3 ( 
	.A1(out_sel[4]), 
	.A2(I4[3]), 
	.B1(out_sel[5]), 
	.B2(I5[3]), 
	.Z(O2[3])); 
	AO_CELL inst_0_4 ( 
	.A1(out_sel[0]), 
	.A2(I0[4]), 
	.B1(out_sel[1]), 
	.B2(I1[4]), 
	.Z(O0[4])); 
	AO_CELL inst_1_4 ( 
	.A1(out_sel[2]), 
	.A2(I2[4]), 
	.B1(out_sel[3]), 
	.B2(I3[4]), 
	.Z(O1[4])); 
	AO_CELL inst_2_4 ( 
	.A1(out_sel[4]), 
	.A2(I4[4]), 
	.B1(out_sel[5]), 
	.B2(I5[4]), 
	.Z(O2[4])); 
	AO_CELL inst_0_5 ( 
	.A1(out_sel[0]), 
	.A2(I0[5]), 
	.B1(out_sel[1]), 
	.B2(I1[5]), 
	.Z(O0[5])); 
	AO_CELL inst_1_5 ( 
	.A1(out_sel[2]), 
	.A2(I2[5]), 
	.B1(out_sel[3]), 
	.B2(I3[5]), 
	.Z(O1[5])); 
	AO_CELL inst_2_5 ( 
	.A1(out_sel[4]), 
	.A2(I4[5]), 
	.B1(out_sel[5]), 
	.B2(I5[5]), 
	.Z(O2[5])); 
	AO_CELL inst_0_6 ( 
	.A1(out_sel[0]), 
	.A2(I0[6]), 
	.B1(out_sel[1]), 
	.B2(I1[6]), 
	.Z(O0[6])); 
	AO_CELL inst_1_6 ( 
	.A1(out_sel[2]), 
	.A2(I2[6]), 
	.B1(out_sel[3]), 
	.B2(I3[6]), 
	.Z(O1[6])); 
	AO_CELL inst_2_6 ( 
	.A1(out_sel[4]), 
	.A2(I4[6]), 
	.B1(out_sel[5]), 
	.B2(I5[6]), 
	.Z(O2[6])); 
	AO_CELL inst_0_7 ( 
	.A1(out_sel[0]), 
	.A2(I0[7]), 
	.B1(out_sel[1]), 
	.B2(I1[7]), 
	.Z(O0[7])); 
	AO_CELL inst_1_7 ( 
	.A1(out_sel[2]), 
	.A2(I2[7]), 
	.B1(out_sel[3]), 
	.B2(I3[7]), 
	.Z(O1[7])); 
	AO_CELL inst_2_7 ( 
	.A1(out_sel[4]), 
	.A2(I4[7]), 
	.B1(out_sel[5]), 
	.B2(I5[7]), 
	.Z(O2[7])); 
	AO_CELL inst_0_8 ( 
	.A1(out_sel[0]), 
	.A2(I0[8]), 
	.B1(out_sel[1]), 
	.B2(I1[8]), 
	.Z(O0[8])); 
	AO_CELL inst_1_8 ( 
	.A1(out_sel[2]), 
	.A2(I2[8]), 
	.B1(out_sel[3]), 
	.B2(I3[8]), 
	.Z(O1[8])); 
	AO_CELL inst_2_8 ( 
	.A1(out_sel[4]), 
	.A2(I4[8]), 
	.B1(out_sel[5]), 
	.B2(I5[8]), 
	.Z(O2[8])); 
	AO_CELL inst_0_9 ( 
	.A1(out_sel[0]), 
	.A2(I0[9]), 
	.B1(out_sel[1]), 
	.B2(I1[9]), 
	.Z(O0[9])); 
	AO_CELL inst_1_9 ( 
	.A1(out_sel[2]), 
	.A2(I2[9]), 
	.B1(out_sel[3]), 
	.B2(I3[9]), 
	.Z(O1[9])); 
	AO_CELL inst_2_9 ( 
	.A1(out_sel[4]), 
	.A2(I4[9]), 
	.B1(out_sel[5]), 
	.B2(I5[9]), 
	.Z(O2[9])); 
	AO_CELL inst_0_10 ( 
	.A1(out_sel[0]), 
	.A2(I0[10]), 
	.B1(out_sel[1]), 
	.B2(I1[10]), 
	.Z(O0[10])); 
	AO_CELL inst_1_10 ( 
	.A1(out_sel[2]), 
	.A2(I2[10]), 
	.B1(out_sel[3]), 
	.B2(I3[10]), 
	.Z(O1[10])); 
	AO_CELL inst_2_10 ( 
	.A1(out_sel[4]), 
	.A2(I4[10]), 
	.B1(out_sel[5]), 
	.B2(I5[10]), 
	.Z(O2[10])); 
	AO_CELL inst_0_11 ( 
	.A1(out_sel[0]), 
	.A2(I0[11]), 
	.B1(out_sel[1]), 
	.B2(I1[11]), 
	.Z(O0[11])); 
	AO_CELL inst_1_11 ( 
	.A1(out_sel[2]), 
	.A2(I2[11]), 
	.B1(out_sel[3]), 
	.B2(I3[11]), 
	.Z(O1[11])); 
	AO_CELL inst_2_11 ( 
	.A1(out_sel[4]), 
	.A2(I4[11]), 
	.B1(out_sel[5]), 
	.B2(I5[11]), 
	.Z(O2[11])); 
	AO_CELL inst_0_12 ( 
	.A1(out_sel[0]), 
	.A2(I0[12]), 
	.B1(out_sel[1]), 
	.B2(I1[12]), 
	.Z(O0[12])); 
	AO_CELL inst_1_12 ( 
	.A1(out_sel[2]), 
	.A2(I2[12]), 
	.B1(out_sel[3]), 
	.B2(I3[12]), 
	.Z(O1[12])); 
	AO_CELL inst_2_12 ( 
	.A1(out_sel[4]), 
	.A2(I4[12]), 
	.B1(out_sel[5]), 
	.B2(I5[12]), 
	.Z(O2[12])); 
	AO_CELL inst_0_13 ( 
	.A1(out_sel[0]), 
	.A2(I0[13]), 
	.B1(out_sel[1]), 
	.B2(I1[13]), 
	.Z(O0[13])); 
	AO_CELL inst_1_13 ( 
	.A1(out_sel[2]), 
	.A2(I2[13]), 
	.B1(out_sel[3]), 
	.B2(I3[13]), 
	.Z(O1[13])); 
	AO_CELL inst_2_13 ( 
	.A1(out_sel[4]), 
	.A2(I4[13]), 
	.B1(out_sel[5]), 
	.B2(I5[13]), 
	.Z(O2[13])); 
	AO_CELL inst_0_14 ( 
	.A1(out_sel[0]), 
	.A2(I0[14]), 
	.B1(out_sel[1]), 
	.B2(I1[14]), 
	.Z(O0[14])); 
	AO_CELL inst_1_14 ( 
	.A1(out_sel[2]), 
	.A2(I2[14]), 
	.B1(out_sel[3]), 
	.B2(I3[14]), 
	.Z(O1[14])); 
	AO_CELL inst_2_14 ( 
	.A1(out_sel[4]), 
	.A2(I4[14]), 
	.B1(out_sel[5]), 
	.B2(I5[14]), 
	.Z(O2[14])); 
	AO_CELL inst_0_15 ( 
	.A1(out_sel[0]), 
	.A2(I0[15]), 
	.B1(out_sel[1]), 
	.B2(I1[15]), 
	.Z(O0[15])); 
	AO_CELL inst_1_15 ( 
	.A1(out_sel[2]), 
	.A2(I2[15]), 
	.B1(out_sel[3]), 
	.B2(I3[15]), 
	.Z(O1[15])); 
	AO_CELL inst_2_15 ( 
	.A1(out_sel[4]), 
	.A2(I4[15]), 
	.B1(out_sel[5]), 
	.B2(I5[15]), 
	.Z(O2[15])); 
	AO_CELL inst_0_16 ( 
	.A1(out_sel[0]), 
	.A2(I0[16]), 
	.B1(out_sel[1]), 
	.B2(I1[16]), 
	.Z(O0[16])); 
	AO_CELL inst_1_16 ( 
	.A1(out_sel[2]), 
	.A2(I2[16]), 
	.B1(out_sel[3]), 
	.B2(I3[16]), 
	.Z(O1[16])); 
	AO_CELL inst_2_16 ( 
	.A1(out_sel[4]), 
	.A2(I4[16]), 
	.B1(out_sel[5]), 
	.B2(I5[16]), 
	.Z(O2[16])); 
	AO_CELL inst_0_valid ( 
	.A1(out_sel[0]), 
	.A2(valid_in[0]), 
	.B1(out_sel[1]), 
	.B2(valid_in[1]), 
	.Z(valid_out[0])); 
	AO_CELL inst_1_valid ( 
	.A1(out_sel[2]), 
	.A2(valid_in[2]), 
	.B1(out_sel[3]), 
	.B2(valid_in[3]), 
	.Z(valid_out[1])); 
	AO_CELL inst_2_valid ( 
	.A1(out_sel[4]), 
	.A2(valid_in[4]), 
	.B1(out_sel[5]), 
	.B2(valid_in[5]), 
	.Z(valid_out[2])); 
endmodule 

module mux_aoi_ready_valid_6_1 ( 
	input logic  [0 : 0] I[5:0], 
	input logic  [2 : 0] S ,
	input logic ready_in,
	output logic ready_out,
	input logic [5:0]  valid_in,
	output logic valid_out,
	output logic  [7 : 0] out_sel,
	output logic [0 : 0] O); 
	logic  [0 : 0] O_int0;
	logic  [0 : 0] O_int1;
	logic  [0 : 0] O_int2;
	logic [2:0] valid_out_temp;

precoder_1_6 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_1_6 u_mux_logic ( 
	.I0 (I[0]),
	.I1 (I[1]),
	.I2 (I[2]),
	.I3 (I[3]),
	.I4 (I[4]),
	.I5 (I[5]),
	.out_sel(out_sel), 
	.valid_in(valid_in),
	.valid_out(valid_out_temp),
	.O0(O_int0), 
	.O1(O_int1), 
	.O2(O_int2)); 
	assign O = (  	O_int0 | 	O_int1 | 	O_int2 	); 
	assign ready_out = ready_in;
	assign valid_out = |valid_out_temp;

endmodule 

module precoder_1_6 (
	input logic  [2 : 0] S ,
	output logic  [7 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		3'd0    :   out_sel = 8'b00000001;
		3'd1    :   out_sel = 8'b00000010;
		3'd2    :   out_sel = 8'b00000100;
		3'd3    :   out_sel = 8'b00001000;
		3'd4    :   out_sel = 8'b00010000;
		3'd5    :   out_sel = 8'b00100000;
		default :   out_sel = 8'b0;
	endcase 
end 

endmodule 

module mux_logic_1_6 ( 
	input logic  [7 : 0] out_sel,
	input logic  [0 : 0] I0, 
	input logic  [0 : 0] I1, 
	input logic  [0 : 0] I2, 
	input logic  [0 : 0] I3, 
	input logic  [0 : 0] I4, 
	input logic  [0 : 0] I5, 
	input logic [5:0] valid_in,
	output logic [2:0] valid_out,
	output logic  [0 : 0] O0, 
	output logic  [0 : 0] O1, 
	output logic  [0 : 0] O2); 
	AO_CELL inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	AO_CELL inst_1_0 ( 
	.A1(out_sel[2]), 
	.A2(I2[0]), 
	.B1(out_sel[3]), 
	.B2(I3[0]), 
	.Z(O1[0])); 
	AO_CELL inst_2_0 ( 
	.A1(out_sel[4]), 
	.A2(I4[0]), 
	.B1(out_sel[5]), 
	.B2(I5[0]), 
	.Z(O2[0])); 
	AO_CELL inst_0_valid ( 
	.A1(out_sel[0]), 
	.A2(valid_in[0]), 
	.B1(out_sel[1]), 
	.B2(valid_in[1]), 
	.Z(valid_out[0])); 
	AO_CELL inst_1_valid ( 
	.A1(out_sel[2]), 
	.A2(valid_in[2]), 
	.B1(out_sel[3]), 
	.B2(valid_in[3]), 
	.Z(valid_out[1])); 
	AO_CELL inst_2_valid ( 
	.A1(out_sel[4]), 
	.A2(valid_in[4]), 
	.B1(out_sel[5]), 
	.B2(valid_in[5]), 
	.Z(valid_out[2])); 
endmodule 

module mux_aoi_ready_valid_2_17 ( 
	input logic  [16 : 0] I[1:0], 
input logic S, 
	input logic ready_in,
	output logic ready_out,
	input logic [1:0]  valid_in,
	output logic valid_out,
	output logic  [1 : 0] out_sel,
	output logic [16 : 0] O); 
	logic  [16 : 0] O_int0;
	logic [0:0] valid_out_temp;

precoder_17_2 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_17_2 u_mux_logic ( 
	.I0 (I[0]),
	.I1 (I[1]),
	.out_sel(out_sel), 
	.valid_in(valid_in),
	.valid_out(valid_out_temp),
	.O0(O_int0)); 
	assign O = (  	O_int0 	); 
	assign ready_out = ready_in;
	assign valid_out = |valid_out_temp;

endmodule 

module precoder_17_2 (
	input logic  [0 : 0] S ,
	output logic  [1 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		1'd0    :   out_sel = 2'b01;
		1'd1    :   out_sel = 2'b10;
		default :   out_sel = 2'b0;
	endcase 
end 

endmodule 

module mux_logic_17_2 ( 
	input logic  [1 : 0] out_sel,
	input logic  [16 : 0] I0, 
	input logic  [16 : 0] I1, 
	input logic [1:0] valid_in,
	output logic [0:0] valid_out,
	output logic  [16 : 0] O0); 
	AO_CELL inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	AO_CELL inst_0_1 ( 
	.A1(out_sel[0]), 
	.A2(I0[1]), 
	.B1(out_sel[1]), 
	.B2(I1[1]), 
	.Z(O0[1])); 
	AO_CELL inst_0_2 ( 
	.A1(out_sel[0]), 
	.A2(I0[2]), 
	.B1(out_sel[1]), 
	.B2(I1[2]), 
	.Z(O0[2])); 
	AO_CELL inst_0_3 ( 
	.A1(out_sel[0]), 
	.A2(I0[3]), 
	.B1(out_sel[1]), 
	.B2(I1[3]), 
	.Z(O0[3])); 
	AO_CELL inst_0_4 ( 
	.A1(out_sel[0]), 
	.A2(I0[4]), 
	.B1(out_sel[1]), 
	.B2(I1[4]), 
	.Z(O0[4])); 
	AO_CELL inst_0_5 ( 
	.A1(out_sel[0]), 
	.A2(I0[5]), 
	.B1(out_sel[1]), 
	.B2(I1[5]), 
	.Z(O0[5])); 
	AO_CELL inst_0_6 ( 
	.A1(out_sel[0]), 
	.A2(I0[6]), 
	.B1(out_sel[1]), 
	.B2(I1[6]), 
	.Z(O0[6])); 
	AO_CELL inst_0_7 ( 
	.A1(out_sel[0]), 
	.A2(I0[7]), 
	.B1(out_sel[1]), 
	.B2(I1[7]), 
	.Z(O0[7])); 
	AO_CELL inst_0_8 ( 
	.A1(out_sel[0]), 
	.A2(I0[8]), 
	.B1(out_sel[1]), 
	.B2(I1[8]), 
	.Z(O0[8])); 
	AO_CELL inst_0_9 ( 
	.A1(out_sel[0]), 
	.A2(I0[9]), 
	.B1(out_sel[1]), 
	.B2(I1[9]), 
	.Z(O0[9])); 
	AO_CELL inst_0_10 ( 
	.A1(out_sel[0]), 
	.A2(I0[10]), 
	.B1(out_sel[1]), 
	.B2(I1[10]), 
	.Z(O0[10])); 
	AO_CELL inst_0_11 ( 
	.A1(out_sel[0]), 
	.A2(I0[11]), 
	.B1(out_sel[1]), 
	.B2(I1[11]), 
	.Z(O0[11])); 
	AO_CELL inst_0_12 ( 
	.A1(out_sel[0]), 
	.A2(I0[12]), 
	.B1(out_sel[1]), 
	.B2(I1[12]), 
	.Z(O0[12])); 
	AO_CELL inst_0_13 ( 
	.A1(out_sel[0]), 
	.A2(I0[13]), 
	.B1(out_sel[1]), 
	.B2(I1[13]), 
	.Z(O0[13])); 
	AO_CELL inst_0_14 ( 
	.A1(out_sel[0]), 
	.A2(I0[14]), 
	.B1(out_sel[1]), 
	.B2(I1[14]), 
	.Z(O0[14])); 
	AO_CELL inst_0_15 ( 
	.A1(out_sel[0]), 
	.A2(I0[15]), 
	.B1(out_sel[1]), 
	.B2(I1[15]), 
	.Z(O0[15])); 
	AO_CELL inst_0_16 ( 
	.A1(out_sel[0]), 
	.A2(I0[16]), 
	.B1(out_sel[1]), 
	.B2(I1[16]), 
	.Z(O0[16])); 
	AO_CELL inst_0_valid ( 
	.A1(out_sel[0]), 
	.A2(valid_in[0]), 
	.B1(out_sel[1]), 
	.B2(valid_in[1]), 
	.Z(valid_out[0])); 
endmodule 

module mux_aoi_ready_valid_2_1 ( 
	input logic  [0 : 0] I[1:0], 
input logic S, 
	input logic ready_in,
	output logic ready_out,
	input logic [1:0]  valid_in,
	output logic valid_out,
	output logic  [1 : 0] out_sel,
	output logic [0 : 0] O); 
	logic  [0 : 0] O_int0;
	logic [0:0] valid_out_temp;

precoder_1_2 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_1_2 u_mux_logic ( 
	.I0 (I[0]),
	.I1 (I[1]),
	.out_sel(out_sel), 
	.valid_in(valid_in),
	.valid_out(valid_out_temp),
	.O0(O_int0)); 
	assign O = (  	O_int0 	); 
	assign ready_out = ready_in;
	assign valid_out = |valid_out_temp;

endmodule 

module precoder_1_2 (
	input logic  [0 : 0] S ,
	output logic  [1 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		1'd0    :   out_sel = 2'b01;
		1'd1    :   out_sel = 2'b10;
		default :   out_sel = 2'b0;
	endcase 
end 

endmodule 

module mux_logic_1_2 ( 
	input logic  [1 : 0] out_sel,
	input logic  [0 : 0] I0, 
	input logic  [0 : 0] I1, 
	input logic [1:0] valid_in,
	output logic [0:0] valid_out,
	output logic  [0 : 0] O0); 
	AO_CELL inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	AO_CELL inst_0_valid ( 
	.A1(out_sel[0]), 
	.A2(valid_in[0]), 
	.B1(out_sel[1]), 
	.B2(valid_in[1]), 
	.Z(valid_out[0])); 
endmodule 

module mux_aoi_7_32 ( 
	input logic  [31 : 0] I[6:0], 
	input logic  [2 : 0] S ,
	output logic  [7 : 0] out_sel,
	output logic [31 : 0] O); 
	logic  [31 : 0] O_int0;
	logic  [31 : 0] O_int1;
	logic  [31 : 0] O_int2;
	logic  [31 : 0] O_int3;

precoder_32_7 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_32_7 u_mux_logic ( 
	.I0 (I[0]),
	.I1 (I[1]),
	.I2 (I[2]),
	.I3 (I[3]),
	.I4 (I[4]),
	.I5 (I[5]),
	.I6 (I[6]),
	.out_sel(out_sel), 
	.O0(O_int0), 
	.O1(O_int1), 
	.O2(O_int2), 
	.O3(O_int3)); 
	assign O = (  	O_int0 | 	O_int1 | 	O_int2 | 	O_int3 	); 

endmodule 

module precoder_32_7 (
	input logic  [2 : 0] S ,
	output logic  [7 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		3'd0    :   out_sel = 8'b00000001;
		3'd1    :   out_sel = 8'b00000010;
		3'd2    :   out_sel = 8'b00000100;
		3'd3    :   out_sel = 8'b00001000;
		3'd4    :   out_sel = 8'b00010000;
		3'd5    :   out_sel = 8'b00100000;
		3'd6    :   out_sel = 8'b01000000;
		default :   out_sel = 8'b0;
	endcase 
end 

endmodule 

module mux_logic_32_7 ( 
	input logic  [7 : 0] out_sel,
	input logic  [31 : 0] I0, 
	input logic  [31 : 0] I1, 
	input logic  [31 : 0] I2, 
	input logic  [31 : 0] I3, 
	input logic  [31 : 0] I4, 
	input logic  [31 : 0] I5, 
	input logic  [31 : 0] I6, 
	output logic  [31 : 0] O0, 
	output logic  [31 : 0] O1, 
	output logic  [31 : 0] O2, 
	output logic  [31 : 0] O3); 
	AO_CELL inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	AO_CELL inst_1_0 ( 
	.A1(out_sel[2]), 
	.A2(I2[0]), 
	.B1(out_sel[3]), 
	.B2(I3[0]), 
	.Z(O1[0])); 
	AO_CELL inst_2_0 ( 
	.A1(out_sel[4]), 
	.A2(I4[0]), 
	.B1(out_sel[5]), 
	.B2(I5[0]), 
	.Z(O2[0])); 
	AN_CELL inst_and_0 ( 
	.A1(out_sel[6]), 
	.A2(I6[0]), 
	.Z(O3[0])); 
	AO_CELL inst_0_1 ( 
	.A1(out_sel[0]), 
	.A2(I0[1]), 
	.B1(out_sel[1]), 
	.B2(I1[1]), 
	.Z(O0[1])); 
	AO_CELL inst_1_1 ( 
	.A1(out_sel[2]), 
	.A2(I2[1]), 
	.B1(out_sel[3]), 
	.B2(I3[1]), 
	.Z(O1[1])); 
	AO_CELL inst_2_1 ( 
	.A1(out_sel[4]), 
	.A2(I4[1]), 
	.B1(out_sel[5]), 
	.B2(I5[1]), 
	.Z(O2[1])); 
	AN_CELL inst_and_1 ( 
	.A1(out_sel[6]), 
	.A2(I6[1]), 
	.Z(O3[1])); 
	AO_CELL inst_0_2 ( 
	.A1(out_sel[0]), 
	.A2(I0[2]), 
	.B1(out_sel[1]), 
	.B2(I1[2]), 
	.Z(O0[2])); 
	AO_CELL inst_1_2 ( 
	.A1(out_sel[2]), 
	.A2(I2[2]), 
	.B1(out_sel[3]), 
	.B2(I3[2]), 
	.Z(O1[2])); 
	AO_CELL inst_2_2 ( 
	.A1(out_sel[4]), 
	.A2(I4[2]), 
	.B1(out_sel[5]), 
	.B2(I5[2]), 
	.Z(O2[2])); 
	AN_CELL inst_and_2 ( 
	.A1(out_sel[6]), 
	.A2(I6[2]), 
	.Z(O3[2])); 
	AO_CELL inst_0_3 ( 
	.A1(out_sel[0]), 
	.A2(I0[3]), 
	.B1(out_sel[1]), 
	.B2(I1[3]), 
	.Z(O0[3])); 
	AO_CELL inst_1_3 ( 
	.A1(out_sel[2]), 
	.A2(I2[3]), 
	.B1(out_sel[3]), 
	.B2(I3[3]), 
	.Z(O1[3])); 
	AO_CELL inst_2_3 ( 
	.A1(out_sel[4]), 
	.A2(I4[3]), 
	.B1(out_sel[5]), 
	.B2(I5[3]), 
	.Z(O2[3])); 
	AN_CELL inst_and_3 ( 
	.A1(out_sel[6]), 
	.A2(I6[3]), 
	.Z(O3[3])); 
	AO_CELL inst_0_4 ( 
	.A1(out_sel[0]), 
	.A2(I0[4]), 
	.B1(out_sel[1]), 
	.B2(I1[4]), 
	.Z(O0[4])); 
	AO_CELL inst_1_4 ( 
	.A1(out_sel[2]), 
	.A2(I2[4]), 
	.B1(out_sel[3]), 
	.B2(I3[4]), 
	.Z(O1[4])); 
	AO_CELL inst_2_4 ( 
	.A1(out_sel[4]), 
	.A2(I4[4]), 
	.B1(out_sel[5]), 
	.B2(I5[4]), 
	.Z(O2[4])); 
	AN_CELL inst_and_4 ( 
	.A1(out_sel[6]), 
	.A2(I6[4]), 
	.Z(O3[4])); 
	AO_CELL inst_0_5 ( 
	.A1(out_sel[0]), 
	.A2(I0[5]), 
	.B1(out_sel[1]), 
	.B2(I1[5]), 
	.Z(O0[5])); 
	AO_CELL inst_1_5 ( 
	.A1(out_sel[2]), 
	.A2(I2[5]), 
	.B1(out_sel[3]), 
	.B2(I3[5]), 
	.Z(O1[5])); 
	AO_CELL inst_2_5 ( 
	.A1(out_sel[4]), 
	.A2(I4[5]), 
	.B1(out_sel[5]), 
	.B2(I5[5]), 
	.Z(O2[5])); 
	AN_CELL inst_and_5 ( 
	.A1(out_sel[6]), 
	.A2(I6[5]), 
	.Z(O3[5])); 
	AO_CELL inst_0_6 ( 
	.A1(out_sel[0]), 
	.A2(I0[6]), 
	.B1(out_sel[1]), 
	.B2(I1[6]), 
	.Z(O0[6])); 
	AO_CELL inst_1_6 ( 
	.A1(out_sel[2]), 
	.A2(I2[6]), 
	.B1(out_sel[3]), 
	.B2(I3[6]), 
	.Z(O1[6])); 
	AO_CELL inst_2_6 ( 
	.A1(out_sel[4]), 
	.A2(I4[6]), 
	.B1(out_sel[5]), 
	.B2(I5[6]), 
	.Z(O2[6])); 
	AN_CELL inst_and_6 ( 
	.A1(out_sel[6]), 
	.A2(I6[6]), 
	.Z(O3[6])); 
	AO_CELL inst_0_7 ( 
	.A1(out_sel[0]), 
	.A2(I0[7]), 
	.B1(out_sel[1]), 
	.B2(I1[7]), 
	.Z(O0[7])); 
	AO_CELL inst_1_7 ( 
	.A1(out_sel[2]), 
	.A2(I2[7]), 
	.B1(out_sel[3]), 
	.B2(I3[7]), 
	.Z(O1[7])); 
	AO_CELL inst_2_7 ( 
	.A1(out_sel[4]), 
	.A2(I4[7]), 
	.B1(out_sel[5]), 
	.B2(I5[7]), 
	.Z(O2[7])); 
	AN_CELL inst_and_7 ( 
	.A1(out_sel[6]), 
	.A2(I6[7]), 
	.Z(O3[7])); 
	AO_CELL inst_0_8 ( 
	.A1(out_sel[0]), 
	.A2(I0[8]), 
	.B1(out_sel[1]), 
	.B2(I1[8]), 
	.Z(O0[8])); 
	AO_CELL inst_1_8 ( 
	.A1(out_sel[2]), 
	.A2(I2[8]), 
	.B1(out_sel[3]), 
	.B2(I3[8]), 
	.Z(O1[8])); 
	AO_CELL inst_2_8 ( 
	.A1(out_sel[4]), 
	.A2(I4[8]), 
	.B1(out_sel[5]), 
	.B2(I5[8]), 
	.Z(O2[8])); 
	AN_CELL inst_and_8 ( 
	.A1(out_sel[6]), 
	.A2(I6[8]), 
	.Z(O3[8])); 
	AO_CELL inst_0_9 ( 
	.A1(out_sel[0]), 
	.A2(I0[9]), 
	.B1(out_sel[1]), 
	.B2(I1[9]), 
	.Z(O0[9])); 
	AO_CELL inst_1_9 ( 
	.A1(out_sel[2]), 
	.A2(I2[9]), 
	.B1(out_sel[3]), 
	.B2(I3[9]), 
	.Z(O1[9])); 
	AO_CELL inst_2_9 ( 
	.A1(out_sel[4]), 
	.A2(I4[9]), 
	.B1(out_sel[5]), 
	.B2(I5[9]), 
	.Z(O2[9])); 
	AN_CELL inst_and_9 ( 
	.A1(out_sel[6]), 
	.A2(I6[9]), 
	.Z(O3[9])); 
	AO_CELL inst_0_10 ( 
	.A1(out_sel[0]), 
	.A2(I0[10]), 
	.B1(out_sel[1]), 
	.B2(I1[10]), 
	.Z(O0[10])); 
	AO_CELL inst_1_10 ( 
	.A1(out_sel[2]), 
	.A2(I2[10]), 
	.B1(out_sel[3]), 
	.B2(I3[10]), 
	.Z(O1[10])); 
	AO_CELL inst_2_10 ( 
	.A1(out_sel[4]), 
	.A2(I4[10]), 
	.B1(out_sel[5]), 
	.B2(I5[10]), 
	.Z(O2[10])); 
	AN_CELL inst_and_10 ( 
	.A1(out_sel[6]), 
	.A2(I6[10]), 
	.Z(O3[10])); 
	AO_CELL inst_0_11 ( 
	.A1(out_sel[0]), 
	.A2(I0[11]), 
	.B1(out_sel[1]), 
	.B2(I1[11]), 
	.Z(O0[11])); 
	AO_CELL inst_1_11 ( 
	.A1(out_sel[2]), 
	.A2(I2[11]), 
	.B1(out_sel[3]), 
	.B2(I3[11]), 
	.Z(O1[11])); 
	AO_CELL inst_2_11 ( 
	.A1(out_sel[4]), 
	.A2(I4[11]), 
	.B1(out_sel[5]), 
	.B2(I5[11]), 
	.Z(O2[11])); 
	AN_CELL inst_and_11 ( 
	.A1(out_sel[6]), 
	.A2(I6[11]), 
	.Z(O3[11])); 
	AO_CELL inst_0_12 ( 
	.A1(out_sel[0]), 
	.A2(I0[12]), 
	.B1(out_sel[1]), 
	.B2(I1[12]), 
	.Z(O0[12])); 
	AO_CELL inst_1_12 ( 
	.A1(out_sel[2]), 
	.A2(I2[12]), 
	.B1(out_sel[3]), 
	.B2(I3[12]), 
	.Z(O1[12])); 
	AO_CELL inst_2_12 ( 
	.A1(out_sel[4]), 
	.A2(I4[12]), 
	.B1(out_sel[5]), 
	.B2(I5[12]), 
	.Z(O2[12])); 
	AN_CELL inst_and_12 ( 
	.A1(out_sel[6]), 
	.A2(I6[12]), 
	.Z(O3[12])); 
	AO_CELL inst_0_13 ( 
	.A1(out_sel[0]), 
	.A2(I0[13]), 
	.B1(out_sel[1]), 
	.B2(I1[13]), 
	.Z(O0[13])); 
	AO_CELL inst_1_13 ( 
	.A1(out_sel[2]), 
	.A2(I2[13]), 
	.B1(out_sel[3]), 
	.B2(I3[13]), 
	.Z(O1[13])); 
	AO_CELL inst_2_13 ( 
	.A1(out_sel[4]), 
	.A2(I4[13]), 
	.B1(out_sel[5]), 
	.B2(I5[13]), 
	.Z(O2[13])); 
	AN_CELL inst_and_13 ( 
	.A1(out_sel[6]), 
	.A2(I6[13]), 
	.Z(O3[13])); 
	AO_CELL inst_0_14 ( 
	.A1(out_sel[0]), 
	.A2(I0[14]), 
	.B1(out_sel[1]), 
	.B2(I1[14]), 
	.Z(O0[14])); 
	AO_CELL inst_1_14 ( 
	.A1(out_sel[2]), 
	.A2(I2[14]), 
	.B1(out_sel[3]), 
	.B2(I3[14]), 
	.Z(O1[14])); 
	AO_CELL inst_2_14 ( 
	.A1(out_sel[4]), 
	.A2(I4[14]), 
	.B1(out_sel[5]), 
	.B2(I5[14]), 
	.Z(O2[14])); 
	AN_CELL inst_and_14 ( 
	.A1(out_sel[6]), 
	.A2(I6[14]), 
	.Z(O3[14])); 
	AO_CELL inst_0_15 ( 
	.A1(out_sel[0]), 
	.A2(I0[15]), 
	.B1(out_sel[1]), 
	.B2(I1[15]), 
	.Z(O0[15])); 
	AO_CELL inst_1_15 ( 
	.A1(out_sel[2]), 
	.A2(I2[15]), 
	.B1(out_sel[3]), 
	.B2(I3[15]), 
	.Z(O1[15])); 
	AO_CELL inst_2_15 ( 
	.A1(out_sel[4]), 
	.A2(I4[15]), 
	.B1(out_sel[5]), 
	.B2(I5[15]), 
	.Z(O2[15])); 
	AN_CELL inst_and_15 ( 
	.A1(out_sel[6]), 
	.A2(I6[15]), 
	.Z(O3[15])); 
	AO_CELL inst_0_16 ( 
	.A1(out_sel[0]), 
	.A2(I0[16]), 
	.B1(out_sel[1]), 
	.B2(I1[16]), 
	.Z(O0[16])); 
	AO_CELL inst_1_16 ( 
	.A1(out_sel[2]), 
	.A2(I2[16]), 
	.B1(out_sel[3]), 
	.B2(I3[16]), 
	.Z(O1[16])); 
	AO_CELL inst_2_16 ( 
	.A1(out_sel[4]), 
	.A2(I4[16]), 
	.B1(out_sel[5]), 
	.B2(I5[16]), 
	.Z(O2[16])); 
	AN_CELL inst_and_16 ( 
	.A1(out_sel[6]), 
	.A2(I6[16]), 
	.Z(O3[16])); 
	AO_CELL inst_0_17 ( 
	.A1(out_sel[0]), 
	.A2(I0[17]), 
	.B1(out_sel[1]), 
	.B2(I1[17]), 
	.Z(O0[17])); 
	AO_CELL inst_1_17 ( 
	.A1(out_sel[2]), 
	.A2(I2[17]), 
	.B1(out_sel[3]), 
	.B2(I3[17]), 
	.Z(O1[17])); 
	AO_CELL inst_2_17 ( 
	.A1(out_sel[4]), 
	.A2(I4[17]), 
	.B1(out_sel[5]), 
	.B2(I5[17]), 
	.Z(O2[17])); 
	AN_CELL inst_and_17 ( 
	.A1(out_sel[6]), 
	.A2(I6[17]), 
	.Z(O3[17])); 
	AO_CELL inst_0_18 ( 
	.A1(out_sel[0]), 
	.A2(I0[18]), 
	.B1(out_sel[1]), 
	.B2(I1[18]), 
	.Z(O0[18])); 
	AO_CELL inst_1_18 ( 
	.A1(out_sel[2]), 
	.A2(I2[18]), 
	.B1(out_sel[3]), 
	.B2(I3[18]), 
	.Z(O1[18])); 
	AO_CELL inst_2_18 ( 
	.A1(out_sel[4]), 
	.A2(I4[18]), 
	.B1(out_sel[5]), 
	.B2(I5[18]), 
	.Z(O2[18])); 
	AN_CELL inst_and_18 ( 
	.A1(out_sel[6]), 
	.A2(I6[18]), 
	.Z(O3[18])); 
	AO_CELL inst_0_19 ( 
	.A1(out_sel[0]), 
	.A2(I0[19]), 
	.B1(out_sel[1]), 
	.B2(I1[19]), 
	.Z(O0[19])); 
	AO_CELL inst_1_19 ( 
	.A1(out_sel[2]), 
	.A2(I2[19]), 
	.B1(out_sel[3]), 
	.B2(I3[19]), 
	.Z(O1[19])); 
	AO_CELL inst_2_19 ( 
	.A1(out_sel[4]), 
	.A2(I4[19]), 
	.B1(out_sel[5]), 
	.B2(I5[19]), 
	.Z(O2[19])); 
	AN_CELL inst_and_19 ( 
	.A1(out_sel[6]), 
	.A2(I6[19]), 
	.Z(O3[19])); 
	AO_CELL inst_0_20 ( 
	.A1(out_sel[0]), 
	.A2(I0[20]), 
	.B1(out_sel[1]), 
	.B2(I1[20]), 
	.Z(O0[20])); 
	AO_CELL inst_1_20 ( 
	.A1(out_sel[2]), 
	.A2(I2[20]), 
	.B1(out_sel[3]), 
	.B2(I3[20]), 
	.Z(O1[20])); 
	AO_CELL inst_2_20 ( 
	.A1(out_sel[4]), 
	.A2(I4[20]), 
	.B1(out_sel[5]), 
	.B2(I5[20]), 
	.Z(O2[20])); 
	AN_CELL inst_and_20 ( 
	.A1(out_sel[6]), 
	.A2(I6[20]), 
	.Z(O3[20])); 
	AO_CELL inst_0_21 ( 
	.A1(out_sel[0]), 
	.A2(I0[21]), 
	.B1(out_sel[1]), 
	.B2(I1[21]), 
	.Z(O0[21])); 
	AO_CELL inst_1_21 ( 
	.A1(out_sel[2]), 
	.A2(I2[21]), 
	.B1(out_sel[3]), 
	.B2(I3[21]), 
	.Z(O1[21])); 
	AO_CELL inst_2_21 ( 
	.A1(out_sel[4]), 
	.A2(I4[21]), 
	.B1(out_sel[5]), 
	.B2(I5[21]), 
	.Z(O2[21])); 
	AN_CELL inst_and_21 ( 
	.A1(out_sel[6]), 
	.A2(I6[21]), 
	.Z(O3[21])); 
	AO_CELL inst_0_22 ( 
	.A1(out_sel[0]), 
	.A2(I0[22]), 
	.B1(out_sel[1]), 
	.B2(I1[22]), 
	.Z(O0[22])); 
	AO_CELL inst_1_22 ( 
	.A1(out_sel[2]), 
	.A2(I2[22]), 
	.B1(out_sel[3]), 
	.B2(I3[22]), 
	.Z(O1[22])); 
	AO_CELL inst_2_22 ( 
	.A1(out_sel[4]), 
	.A2(I4[22]), 
	.B1(out_sel[5]), 
	.B2(I5[22]), 
	.Z(O2[22])); 
	AN_CELL inst_and_22 ( 
	.A1(out_sel[6]), 
	.A2(I6[22]), 
	.Z(O3[22])); 
	AO_CELL inst_0_23 ( 
	.A1(out_sel[0]), 
	.A2(I0[23]), 
	.B1(out_sel[1]), 
	.B2(I1[23]), 
	.Z(O0[23])); 
	AO_CELL inst_1_23 ( 
	.A1(out_sel[2]), 
	.A2(I2[23]), 
	.B1(out_sel[3]), 
	.B2(I3[23]), 
	.Z(O1[23])); 
	AO_CELL inst_2_23 ( 
	.A1(out_sel[4]), 
	.A2(I4[23]), 
	.B1(out_sel[5]), 
	.B2(I5[23]), 
	.Z(O2[23])); 
	AN_CELL inst_and_23 ( 
	.A1(out_sel[6]), 
	.A2(I6[23]), 
	.Z(O3[23])); 
	AO_CELL inst_0_24 ( 
	.A1(out_sel[0]), 
	.A2(I0[24]), 
	.B1(out_sel[1]), 
	.B2(I1[24]), 
	.Z(O0[24])); 
	AO_CELL inst_1_24 ( 
	.A1(out_sel[2]), 
	.A2(I2[24]), 
	.B1(out_sel[3]), 
	.B2(I3[24]), 
	.Z(O1[24])); 
	AO_CELL inst_2_24 ( 
	.A1(out_sel[4]), 
	.A2(I4[24]), 
	.B1(out_sel[5]), 
	.B2(I5[24]), 
	.Z(O2[24])); 
	AN_CELL inst_and_24 ( 
	.A1(out_sel[6]), 
	.A2(I6[24]), 
	.Z(O3[24])); 
	AO_CELL inst_0_25 ( 
	.A1(out_sel[0]), 
	.A2(I0[25]), 
	.B1(out_sel[1]), 
	.B2(I1[25]), 
	.Z(O0[25])); 
	AO_CELL inst_1_25 ( 
	.A1(out_sel[2]), 
	.A2(I2[25]), 
	.B1(out_sel[3]), 
	.B2(I3[25]), 
	.Z(O1[25])); 
	AO_CELL inst_2_25 ( 
	.A1(out_sel[4]), 
	.A2(I4[25]), 
	.B1(out_sel[5]), 
	.B2(I5[25]), 
	.Z(O2[25])); 
	AN_CELL inst_and_25 ( 
	.A1(out_sel[6]), 
	.A2(I6[25]), 
	.Z(O3[25])); 
	AO_CELL inst_0_26 ( 
	.A1(out_sel[0]), 
	.A2(I0[26]), 
	.B1(out_sel[1]), 
	.B2(I1[26]), 
	.Z(O0[26])); 
	AO_CELL inst_1_26 ( 
	.A1(out_sel[2]), 
	.A2(I2[26]), 
	.B1(out_sel[3]), 
	.B2(I3[26]), 
	.Z(O1[26])); 
	AO_CELL inst_2_26 ( 
	.A1(out_sel[4]), 
	.A2(I4[26]), 
	.B1(out_sel[5]), 
	.B2(I5[26]), 
	.Z(O2[26])); 
	AN_CELL inst_and_26 ( 
	.A1(out_sel[6]), 
	.A2(I6[26]), 
	.Z(O3[26])); 
	AO_CELL inst_0_27 ( 
	.A1(out_sel[0]), 
	.A2(I0[27]), 
	.B1(out_sel[1]), 
	.B2(I1[27]), 
	.Z(O0[27])); 
	AO_CELL inst_1_27 ( 
	.A1(out_sel[2]), 
	.A2(I2[27]), 
	.B1(out_sel[3]), 
	.B2(I3[27]), 
	.Z(O1[27])); 
	AO_CELL inst_2_27 ( 
	.A1(out_sel[4]), 
	.A2(I4[27]), 
	.B1(out_sel[5]), 
	.B2(I5[27]), 
	.Z(O2[27])); 
	AN_CELL inst_and_27 ( 
	.A1(out_sel[6]), 
	.A2(I6[27]), 
	.Z(O3[27])); 
	AO_CELL inst_0_28 ( 
	.A1(out_sel[0]), 
	.A2(I0[28]), 
	.B1(out_sel[1]), 
	.B2(I1[28]), 
	.Z(O0[28])); 
	AO_CELL inst_1_28 ( 
	.A1(out_sel[2]), 
	.A2(I2[28]), 
	.B1(out_sel[3]), 
	.B2(I3[28]), 
	.Z(O1[28])); 
	AO_CELL inst_2_28 ( 
	.A1(out_sel[4]), 
	.A2(I4[28]), 
	.B1(out_sel[5]), 
	.B2(I5[28]), 
	.Z(O2[28])); 
	AN_CELL inst_and_28 ( 
	.A1(out_sel[6]), 
	.A2(I6[28]), 
	.Z(O3[28])); 
	AO_CELL inst_0_29 ( 
	.A1(out_sel[0]), 
	.A2(I0[29]), 
	.B1(out_sel[1]), 
	.B2(I1[29]), 
	.Z(O0[29])); 
	AO_CELL inst_1_29 ( 
	.A1(out_sel[2]), 
	.A2(I2[29]), 
	.B1(out_sel[3]), 
	.B2(I3[29]), 
	.Z(O1[29])); 
	AO_CELL inst_2_29 ( 
	.A1(out_sel[4]), 
	.A2(I4[29]), 
	.B1(out_sel[5]), 
	.B2(I5[29]), 
	.Z(O2[29])); 
	AN_CELL inst_and_29 ( 
	.A1(out_sel[6]), 
	.A2(I6[29]), 
	.Z(O3[29])); 
	AO_CELL inst_0_30 ( 
	.A1(out_sel[0]), 
	.A2(I0[30]), 
	.B1(out_sel[1]), 
	.B2(I1[30]), 
	.Z(O0[30])); 
	AO_CELL inst_1_30 ( 
	.A1(out_sel[2]), 
	.A2(I2[30]), 
	.B1(out_sel[3]), 
	.B2(I3[30]), 
	.Z(O1[30])); 
	AO_CELL inst_2_30 ( 
	.A1(out_sel[4]), 
	.A2(I4[30]), 
	.B1(out_sel[5]), 
	.B2(I5[30]), 
	.Z(O2[30])); 
	AN_CELL inst_and_30 ( 
	.A1(out_sel[6]), 
	.A2(I6[30]), 
	.Z(O3[30])); 
	AO_CELL inst_0_31 ( 
	.A1(out_sel[0]), 
	.A2(I0[31]), 
	.B1(out_sel[1]), 
	.B2(I1[31]), 
	.Z(O0[31])); 
	AO_CELL inst_1_31 ( 
	.A1(out_sel[2]), 
	.A2(I2[31]), 
	.B1(out_sel[3]), 
	.B2(I3[31]), 
	.Z(O1[31])); 
	AO_CELL inst_2_31 ( 
	.A1(out_sel[4]), 
	.A2(I4[31]), 
	.B1(out_sel[5]), 
	.B2(I5[31]), 
	.Z(O2[31])); 
	AN_CELL inst_and_31 ( 
	.A1(out_sel[6]), 
	.A2(I6[31]), 
	.Z(O3[31])); 
endmodule 

module mux_aoi_6_32 ( 
	input logic  [31 : 0] I[5:0], 
	input logic  [2 : 0] S ,
	output logic  [7 : 0] out_sel,
	output logic [31 : 0] O); 
	logic  [31 : 0] O_int0;
	logic  [31 : 0] O_int1;
	logic  [31 : 0] O_int2;

precoder_32_6 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_32_6 u_mux_logic ( 
	.I0 (I[0]),
	.I1 (I[1]),
	.I2 (I[2]),
	.I3 (I[3]),
	.I4 (I[4]),
	.I5 (I[5]),
	.out_sel(out_sel), 
	.O0(O_int0), 
	.O1(O_int1), 
	.O2(O_int2)); 
	assign O = (  	O_int0 | 	O_int1 | 	O_int2 	); 

endmodule 

module precoder_32_6 (
	input logic  [2 : 0] S ,
	output logic  [7 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		3'd0    :   out_sel = 8'b00000001;
		3'd1    :   out_sel = 8'b00000010;
		3'd2    :   out_sel = 8'b00000100;
		3'd3    :   out_sel = 8'b00001000;
		3'd4    :   out_sel = 8'b00010000;
		3'd5    :   out_sel = 8'b00100000;
		default :   out_sel = 8'b0;
	endcase 
end 

endmodule 

module mux_logic_32_6 ( 
	input logic  [7 : 0] out_sel,
	input logic  [31 : 0] I0, 
	input logic  [31 : 0] I1, 
	input logic  [31 : 0] I2, 
	input logic  [31 : 0] I3, 
	input logic  [31 : 0] I4, 
	input logic  [31 : 0] I5, 
	output logic  [31 : 0] O0, 
	output logic  [31 : 0] O1, 
	output logic  [31 : 0] O2); 
	AO_CELL inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	AO_CELL inst_1_0 ( 
	.A1(out_sel[2]), 
	.A2(I2[0]), 
	.B1(out_sel[3]), 
	.B2(I3[0]), 
	.Z(O1[0])); 
	AO_CELL inst_2_0 ( 
	.A1(out_sel[4]), 
	.A2(I4[0]), 
	.B1(out_sel[5]), 
	.B2(I5[0]), 
	.Z(O2[0])); 
	AO_CELL inst_0_1 ( 
	.A1(out_sel[0]), 
	.A2(I0[1]), 
	.B1(out_sel[1]), 
	.B2(I1[1]), 
	.Z(O0[1])); 
	AO_CELL inst_1_1 ( 
	.A1(out_sel[2]), 
	.A2(I2[1]), 
	.B1(out_sel[3]), 
	.B2(I3[1]), 
	.Z(O1[1])); 
	AO_CELL inst_2_1 ( 
	.A1(out_sel[4]), 
	.A2(I4[1]), 
	.B1(out_sel[5]), 
	.B2(I5[1]), 
	.Z(O2[1])); 
	AO_CELL inst_0_2 ( 
	.A1(out_sel[0]), 
	.A2(I0[2]), 
	.B1(out_sel[1]), 
	.B2(I1[2]), 
	.Z(O0[2])); 
	AO_CELL inst_1_2 ( 
	.A1(out_sel[2]), 
	.A2(I2[2]), 
	.B1(out_sel[3]), 
	.B2(I3[2]), 
	.Z(O1[2])); 
	AO_CELL inst_2_2 ( 
	.A1(out_sel[4]), 
	.A2(I4[2]), 
	.B1(out_sel[5]), 
	.B2(I5[2]), 
	.Z(O2[2])); 
	AO_CELL inst_0_3 ( 
	.A1(out_sel[0]), 
	.A2(I0[3]), 
	.B1(out_sel[1]), 
	.B2(I1[3]), 
	.Z(O0[3])); 
	AO_CELL inst_1_3 ( 
	.A1(out_sel[2]), 
	.A2(I2[3]), 
	.B1(out_sel[3]), 
	.B2(I3[3]), 
	.Z(O1[3])); 
	AO_CELL inst_2_3 ( 
	.A1(out_sel[4]), 
	.A2(I4[3]), 
	.B1(out_sel[5]), 
	.B2(I5[3]), 
	.Z(O2[3])); 
	AO_CELL inst_0_4 ( 
	.A1(out_sel[0]), 
	.A2(I0[4]), 
	.B1(out_sel[1]), 
	.B2(I1[4]), 
	.Z(O0[4])); 
	AO_CELL inst_1_4 ( 
	.A1(out_sel[2]), 
	.A2(I2[4]), 
	.B1(out_sel[3]), 
	.B2(I3[4]), 
	.Z(O1[4])); 
	AO_CELL inst_2_4 ( 
	.A1(out_sel[4]), 
	.A2(I4[4]), 
	.B1(out_sel[5]), 
	.B2(I5[4]), 
	.Z(O2[4])); 
	AO_CELL inst_0_5 ( 
	.A1(out_sel[0]), 
	.A2(I0[5]), 
	.B1(out_sel[1]), 
	.B2(I1[5]), 
	.Z(O0[5])); 
	AO_CELL inst_1_5 ( 
	.A1(out_sel[2]), 
	.A2(I2[5]), 
	.B1(out_sel[3]), 
	.B2(I3[5]), 
	.Z(O1[5])); 
	AO_CELL inst_2_5 ( 
	.A1(out_sel[4]), 
	.A2(I4[5]), 
	.B1(out_sel[5]), 
	.B2(I5[5]), 
	.Z(O2[5])); 
	AO_CELL inst_0_6 ( 
	.A1(out_sel[0]), 
	.A2(I0[6]), 
	.B1(out_sel[1]), 
	.B2(I1[6]), 
	.Z(O0[6])); 
	AO_CELL inst_1_6 ( 
	.A1(out_sel[2]), 
	.A2(I2[6]), 
	.B1(out_sel[3]), 
	.B2(I3[6]), 
	.Z(O1[6])); 
	AO_CELL inst_2_6 ( 
	.A1(out_sel[4]), 
	.A2(I4[6]), 
	.B1(out_sel[5]), 
	.B2(I5[6]), 
	.Z(O2[6])); 
	AO_CELL inst_0_7 ( 
	.A1(out_sel[0]), 
	.A2(I0[7]), 
	.B1(out_sel[1]), 
	.B2(I1[7]), 
	.Z(O0[7])); 
	AO_CELL inst_1_7 ( 
	.A1(out_sel[2]), 
	.A2(I2[7]), 
	.B1(out_sel[3]), 
	.B2(I3[7]), 
	.Z(O1[7])); 
	AO_CELL inst_2_7 ( 
	.A1(out_sel[4]), 
	.A2(I4[7]), 
	.B1(out_sel[5]), 
	.B2(I5[7]), 
	.Z(O2[7])); 
	AO_CELL inst_0_8 ( 
	.A1(out_sel[0]), 
	.A2(I0[8]), 
	.B1(out_sel[1]), 
	.B2(I1[8]), 
	.Z(O0[8])); 
	AO_CELL inst_1_8 ( 
	.A1(out_sel[2]), 
	.A2(I2[8]), 
	.B1(out_sel[3]), 
	.B2(I3[8]), 
	.Z(O1[8])); 
	AO_CELL inst_2_8 ( 
	.A1(out_sel[4]), 
	.A2(I4[8]), 
	.B1(out_sel[5]), 
	.B2(I5[8]), 
	.Z(O2[8])); 
	AO_CELL inst_0_9 ( 
	.A1(out_sel[0]), 
	.A2(I0[9]), 
	.B1(out_sel[1]), 
	.B2(I1[9]), 
	.Z(O0[9])); 
	AO_CELL inst_1_9 ( 
	.A1(out_sel[2]), 
	.A2(I2[9]), 
	.B1(out_sel[3]), 
	.B2(I3[9]), 
	.Z(O1[9])); 
	AO_CELL inst_2_9 ( 
	.A1(out_sel[4]), 
	.A2(I4[9]), 
	.B1(out_sel[5]), 
	.B2(I5[9]), 
	.Z(O2[9])); 
	AO_CELL inst_0_10 ( 
	.A1(out_sel[0]), 
	.A2(I0[10]), 
	.B1(out_sel[1]), 
	.B2(I1[10]), 
	.Z(O0[10])); 
	AO_CELL inst_1_10 ( 
	.A1(out_sel[2]), 
	.A2(I2[10]), 
	.B1(out_sel[3]), 
	.B2(I3[10]), 
	.Z(O1[10])); 
	AO_CELL inst_2_10 ( 
	.A1(out_sel[4]), 
	.A2(I4[10]), 
	.B1(out_sel[5]), 
	.B2(I5[10]), 
	.Z(O2[10])); 
	AO_CELL inst_0_11 ( 
	.A1(out_sel[0]), 
	.A2(I0[11]), 
	.B1(out_sel[1]), 
	.B2(I1[11]), 
	.Z(O0[11])); 
	AO_CELL inst_1_11 ( 
	.A1(out_sel[2]), 
	.A2(I2[11]), 
	.B1(out_sel[3]), 
	.B2(I3[11]), 
	.Z(O1[11])); 
	AO_CELL inst_2_11 ( 
	.A1(out_sel[4]), 
	.A2(I4[11]), 
	.B1(out_sel[5]), 
	.B2(I5[11]), 
	.Z(O2[11])); 
	AO_CELL inst_0_12 ( 
	.A1(out_sel[0]), 
	.A2(I0[12]), 
	.B1(out_sel[1]), 
	.B2(I1[12]), 
	.Z(O0[12])); 
	AO_CELL inst_1_12 ( 
	.A1(out_sel[2]), 
	.A2(I2[12]), 
	.B1(out_sel[3]), 
	.B2(I3[12]), 
	.Z(O1[12])); 
	AO_CELL inst_2_12 ( 
	.A1(out_sel[4]), 
	.A2(I4[12]), 
	.B1(out_sel[5]), 
	.B2(I5[12]), 
	.Z(O2[12])); 
	AO_CELL inst_0_13 ( 
	.A1(out_sel[0]), 
	.A2(I0[13]), 
	.B1(out_sel[1]), 
	.B2(I1[13]), 
	.Z(O0[13])); 
	AO_CELL inst_1_13 ( 
	.A1(out_sel[2]), 
	.A2(I2[13]), 
	.B1(out_sel[3]), 
	.B2(I3[13]), 
	.Z(O1[13])); 
	AO_CELL inst_2_13 ( 
	.A1(out_sel[4]), 
	.A2(I4[13]), 
	.B1(out_sel[5]), 
	.B2(I5[13]), 
	.Z(O2[13])); 
	AO_CELL inst_0_14 ( 
	.A1(out_sel[0]), 
	.A2(I0[14]), 
	.B1(out_sel[1]), 
	.B2(I1[14]), 
	.Z(O0[14])); 
	AO_CELL inst_1_14 ( 
	.A1(out_sel[2]), 
	.A2(I2[14]), 
	.B1(out_sel[3]), 
	.B2(I3[14]), 
	.Z(O1[14])); 
	AO_CELL inst_2_14 ( 
	.A1(out_sel[4]), 
	.A2(I4[14]), 
	.B1(out_sel[5]), 
	.B2(I5[14]), 
	.Z(O2[14])); 
	AO_CELL inst_0_15 ( 
	.A1(out_sel[0]), 
	.A2(I0[15]), 
	.B1(out_sel[1]), 
	.B2(I1[15]), 
	.Z(O0[15])); 
	AO_CELL inst_1_15 ( 
	.A1(out_sel[2]), 
	.A2(I2[15]), 
	.B1(out_sel[3]), 
	.B2(I3[15]), 
	.Z(O1[15])); 
	AO_CELL inst_2_15 ( 
	.A1(out_sel[4]), 
	.A2(I4[15]), 
	.B1(out_sel[5]), 
	.B2(I5[15]), 
	.Z(O2[15])); 
	AO_CELL inst_0_16 ( 
	.A1(out_sel[0]), 
	.A2(I0[16]), 
	.B1(out_sel[1]), 
	.B2(I1[16]), 
	.Z(O0[16])); 
	AO_CELL inst_1_16 ( 
	.A1(out_sel[2]), 
	.A2(I2[16]), 
	.B1(out_sel[3]), 
	.B2(I3[16]), 
	.Z(O1[16])); 
	AO_CELL inst_2_16 ( 
	.A1(out_sel[4]), 
	.A2(I4[16]), 
	.B1(out_sel[5]), 
	.B2(I5[16]), 
	.Z(O2[16])); 
	AO_CELL inst_0_17 ( 
	.A1(out_sel[0]), 
	.A2(I0[17]), 
	.B1(out_sel[1]), 
	.B2(I1[17]), 
	.Z(O0[17])); 
	AO_CELL inst_1_17 ( 
	.A1(out_sel[2]), 
	.A2(I2[17]), 
	.B1(out_sel[3]), 
	.B2(I3[17]), 
	.Z(O1[17])); 
	AO_CELL inst_2_17 ( 
	.A1(out_sel[4]), 
	.A2(I4[17]), 
	.B1(out_sel[5]), 
	.B2(I5[17]), 
	.Z(O2[17])); 
	AO_CELL inst_0_18 ( 
	.A1(out_sel[0]), 
	.A2(I0[18]), 
	.B1(out_sel[1]), 
	.B2(I1[18]), 
	.Z(O0[18])); 
	AO_CELL inst_1_18 ( 
	.A1(out_sel[2]), 
	.A2(I2[18]), 
	.B1(out_sel[3]), 
	.B2(I3[18]), 
	.Z(O1[18])); 
	AO_CELL inst_2_18 ( 
	.A1(out_sel[4]), 
	.A2(I4[18]), 
	.B1(out_sel[5]), 
	.B2(I5[18]), 
	.Z(O2[18])); 
	AO_CELL inst_0_19 ( 
	.A1(out_sel[0]), 
	.A2(I0[19]), 
	.B1(out_sel[1]), 
	.B2(I1[19]), 
	.Z(O0[19])); 
	AO_CELL inst_1_19 ( 
	.A1(out_sel[2]), 
	.A2(I2[19]), 
	.B1(out_sel[3]), 
	.B2(I3[19]), 
	.Z(O1[19])); 
	AO_CELL inst_2_19 ( 
	.A1(out_sel[4]), 
	.A2(I4[19]), 
	.B1(out_sel[5]), 
	.B2(I5[19]), 
	.Z(O2[19])); 
	AO_CELL inst_0_20 ( 
	.A1(out_sel[0]), 
	.A2(I0[20]), 
	.B1(out_sel[1]), 
	.B2(I1[20]), 
	.Z(O0[20])); 
	AO_CELL inst_1_20 ( 
	.A1(out_sel[2]), 
	.A2(I2[20]), 
	.B1(out_sel[3]), 
	.B2(I3[20]), 
	.Z(O1[20])); 
	AO_CELL inst_2_20 ( 
	.A1(out_sel[4]), 
	.A2(I4[20]), 
	.B1(out_sel[5]), 
	.B2(I5[20]), 
	.Z(O2[20])); 
	AO_CELL inst_0_21 ( 
	.A1(out_sel[0]), 
	.A2(I0[21]), 
	.B1(out_sel[1]), 
	.B2(I1[21]), 
	.Z(O0[21])); 
	AO_CELL inst_1_21 ( 
	.A1(out_sel[2]), 
	.A2(I2[21]), 
	.B1(out_sel[3]), 
	.B2(I3[21]), 
	.Z(O1[21])); 
	AO_CELL inst_2_21 ( 
	.A1(out_sel[4]), 
	.A2(I4[21]), 
	.B1(out_sel[5]), 
	.B2(I5[21]), 
	.Z(O2[21])); 
	AO_CELL inst_0_22 ( 
	.A1(out_sel[0]), 
	.A2(I0[22]), 
	.B1(out_sel[1]), 
	.B2(I1[22]), 
	.Z(O0[22])); 
	AO_CELL inst_1_22 ( 
	.A1(out_sel[2]), 
	.A2(I2[22]), 
	.B1(out_sel[3]), 
	.B2(I3[22]), 
	.Z(O1[22])); 
	AO_CELL inst_2_22 ( 
	.A1(out_sel[4]), 
	.A2(I4[22]), 
	.B1(out_sel[5]), 
	.B2(I5[22]), 
	.Z(O2[22])); 
	AO_CELL inst_0_23 ( 
	.A1(out_sel[0]), 
	.A2(I0[23]), 
	.B1(out_sel[1]), 
	.B2(I1[23]), 
	.Z(O0[23])); 
	AO_CELL inst_1_23 ( 
	.A1(out_sel[2]), 
	.A2(I2[23]), 
	.B1(out_sel[3]), 
	.B2(I3[23]), 
	.Z(O1[23])); 
	AO_CELL inst_2_23 ( 
	.A1(out_sel[4]), 
	.A2(I4[23]), 
	.B1(out_sel[5]), 
	.B2(I5[23]), 
	.Z(O2[23])); 
	AO_CELL inst_0_24 ( 
	.A1(out_sel[0]), 
	.A2(I0[24]), 
	.B1(out_sel[1]), 
	.B2(I1[24]), 
	.Z(O0[24])); 
	AO_CELL inst_1_24 ( 
	.A1(out_sel[2]), 
	.A2(I2[24]), 
	.B1(out_sel[3]), 
	.B2(I3[24]), 
	.Z(O1[24])); 
	AO_CELL inst_2_24 ( 
	.A1(out_sel[4]), 
	.A2(I4[24]), 
	.B1(out_sel[5]), 
	.B2(I5[24]), 
	.Z(O2[24])); 
	AO_CELL inst_0_25 ( 
	.A1(out_sel[0]), 
	.A2(I0[25]), 
	.B1(out_sel[1]), 
	.B2(I1[25]), 
	.Z(O0[25])); 
	AO_CELL inst_1_25 ( 
	.A1(out_sel[2]), 
	.A2(I2[25]), 
	.B1(out_sel[3]), 
	.B2(I3[25]), 
	.Z(O1[25])); 
	AO_CELL inst_2_25 ( 
	.A1(out_sel[4]), 
	.A2(I4[25]), 
	.B1(out_sel[5]), 
	.B2(I5[25]), 
	.Z(O2[25])); 
	AO_CELL inst_0_26 ( 
	.A1(out_sel[0]), 
	.A2(I0[26]), 
	.B1(out_sel[1]), 
	.B2(I1[26]), 
	.Z(O0[26])); 
	AO_CELL inst_1_26 ( 
	.A1(out_sel[2]), 
	.A2(I2[26]), 
	.B1(out_sel[3]), 
	.B2(I3[26]), 
	.Z(O1[26])); 
	AO_CELL inst_2_26 ( 
	.A1(out_sel[4]), 
	.A2(I4[26]), 
	.B1(out_sel[5]), 
	.B2(I5[26]), 
	.Z(O2[26])); 
	AO_CELL inst_0_27 ( 
	.A1(out_sel[0]), 
	.A2(I0[27]), 
	.B1(out_sel[1]), 
	.B2(I1[27]), 
	.Z(O0[27])); 
	AO_CELL inst_1_27 ( 
	.A1(out_sel[2]), 
	.A2(I2[27]), 
	.B1(out_sel[3]), 
	.B2(I3[27]), 
	.Z(O1[27])); 
	AO_CELL inst_2_27 ( 
	.A1(out_sel[4]), 
	.A2(I4[27]), 
	.B1(out_sel[5]), 
	.B2(I5[27]), 
	.Z(O2[27])); 
	AO_CELL inst_0_28 ( 
	.A1(out_sel[0]), 
	.A2(I0[28]), 
	.B1(out_sel[1]), 
	.B2(I1[28]), 
	.Z(O0[28])); 
	AO_CELL inst_1_28 ( 
	.A1(out_sel[2]), 
	.A2(I2[28]), 
	.B1(out_sel[3]), 
	.B2(I3[28]), 
	.Z(O1[28])); 
	AO_CELL inst_2_28 ( 
	.A1(out_sel[4]), 
	.A2(I4[28]), 
	.B1(out_sel[5]), 
	.B2(I5[28]), 
	.Z(O2[28])); 
	AO_CELL inst_0_29 ( 
	.A1(out_sel[0]), 
	.A2(I0[29]), 
	.B1(out_sel[1]), 
	.B2(I1[29]), 
	.Z(O0[29])); 
	AO_CELL inst_1_29 ( 
	.A1(out_sel[2]), 
	.A2(I2[29]), 
	.B1(out_sel[3]), 
	.B2(I3[29]), 
	.Z(O1[29])); 
	AO_CELL inst_2_29 ( 
	.A1(out_sel[4]), 
	.A2(I4[29]), 
	.B1(out_sel[5]), 
	.B2(I5[29]), 
	.Z(O2[29])); 
	AO_CELL inst_0_30 ( 
	.A1(out_sel[0]), 
	.A2(I0[30]), 
	.B1(out_sel[1]), 
	.B2(I1[30]), 
	.Z(O0[30])); 
	AO_CELL inst_1_30 ( 
	.A1(out_sel[2]), 
	.A2(I2[30]), 
	.B1(out_sel[3]), 
	.B2(I3[30]), 
	.Z(O1[30])); 
	AO_CELL inst_2_30 ( 
	.A1(out_sel[4]), 
	.A2(I4[30]), 
	.B1(out_sel[5]), 
	.B2(I5[30]), 
	.Z(O2[30])); 
	AO_CELL inst_0_31 ( 
	.A1(out_sel[0]), 
	.A2(I0[31]), 
	.B1(out_sel[1]), 
	.B2(I1[31]), 
	.Z(O0[31])); 
	AO_CELL inst_1_31 ( 
	.A1(out_sel[2]), 
	.A2(I2[31]), 
	.B1(out_sel[3]), 
	.B2(I3[31]), 
	.Z(O1[31])); 
	AO_CELL inst_2_31 ( 
	.A1(out_sel[4]), 
	.A2(I4[31]), 
	.B1(out_sel[5]), 
	.B2(I5[31]), 
	.Z(O2[31])); 
endmodule 

module mux_aoi_47_32 ( 
	input logic  [31 : 0] I[46:0], 
	input logic  [5 : 0] S ,
	output logic  [63 : 0] out_sel,
	output logic [31 : 0] O); 
	logic  [31 : 0] O_int0;
	logic  [31 : 0] O_int1;
	logic  [31 : 0] O_int2;
	logic  [31 : 0] O_int3;
	logic  [31 : 0] O_int4;
	logic  [31 : 0] O_int5;
	logic  [31 : 0] O_int6;
	logic  [31 : 0] O_int7;
	logic  [31 : 0] O_int8;
	logic  [31 : 0] O_int9;
	logic  [31 : 0] O_int10;
	logic  [31 : 0] O_int11;
	logic  [31 : 0] O_int12;
	logic  [31 : 0] O_int13;
	logic  [31 : 0] O_int14;
	logic  [31 : 0] O_int15;
	logic  [31 : 0] O_int16;
	logic  [31 : 0] O_int17;
	logic  [31 : 0] O_int18;
	logic  [31 : 0] O_int19;
	logic  [31 : 0] O_int20;
	logic  [31 : 0] O_int21;
	logic  [31 : 0] O_int22;
	logic  [31 : 0] O_int23;

precoder_32_47 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_32_47 u_mux_logic ( 
	.I0 (I[0]),
	.I1 (I[1]),
	.I2 (I[2]),
	.I3 (I[3]),
	.I4 (I[4]),
	.I5 (I[5]),
	.I6 (I[6]),
	.I7 (I[7]),
	.I8 (I[8]),
	.I9 (I[9]),
	.I10 (I[10]),
	.I11 (I[11]),
	.I12 (I[12]),
	.I13 (I[13]),
	.I14 (I[14]),
	.I15 (I[15]),
	.I16 (I[16]),
	.I17 (I[17]),
	.I18 (I[18]),
	.I19 (I[19]),
	.I20 (I[20]),
	.I21 (I[21]),
	.I22 (I[22]),
	.I23 (I[23]),
	.I24 (I[24]),
	.I25 (I[25]),
	.I26 (I[26]),
	.I27 (I[27]),
	.I28 (I[28]),
	.I29 (I[29]),
	.I30 (I[30]),
	.I31 (I[31]),
	.I32 (I[32]),
	.I33 (I[33]),
	.I34 (I[34]),
	.I35 (I[35]),
	.I36 (I[36]),
	.I37 (I[37]),
	.I38 (I[38]),
	.I39 (I[39]),
	.I40 (I[40]),
	.I41 (I[41]),
	.I42 (I[42]),
	.I43 (I[43]),
	.I44 (I[44]),
	.I45 (I[45]),
	.I46 (I[46]),
	.out_sel(out_sel), 
	.O0(O_int0), 
	.O1(O_int1), 
	.O2(O_int2), 
	.O3(O_int3), 
	.O4(O_int4), 
	.O5(O_int5), 
	.O6(O_int6), 
	.O7(O_int7), 
	.O8(O_int8), 
	.O9(O_int9), 
	.O10(O_int10), 
	.O11(O_int11), 
	.O12(O_int12), 
	.O13(O_int13), 
	.O14(O_int14), 
	.O15(O_int15), 
	.O16(O_int16), 
	.O17(O_int17), 
	.O18(O_int18), 
	.O19(O_int19), 
	.O20(O_int20), 
	.O21(O_int21), 
	.O22(O_int22), 
	.O23(O_int23)); 
	assign O = (  	O_int0 | 	O_int1 | 	O_int2 | 	O_int3 | 	O_int4 | 	O_int5 | 	O_int6 | 	O_int7 | 	O_int8 | 	O_int9 | 	O_int10 | 	O_int11 | 	O_int12 | 	O_int13 | 	O_int14 | 	O_int15 | 	O_int16 | 	O_int17 | 	O_int18 | 	O_int19 | 	O_int20 | 	O_int21 | 	O_int22 | 	O_int23 	); 

endmodule 

module precoder_32_47 (
	input logic  [5 : 0] S ,
	output logic  [63 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		6'd0    :   out_sel = 64'b0000000000000000000000000000000000000000000000000000000000000001;
		6'd1    :   out_sel = 64'b0000000000000000000000000000000000000000000000000000000000000010;
		6'd2    :   out_sel = 64'b0000000000000000000000000000000000000000000000000000000000000100;
		6'd3    :   out_sel = 64'b0000000000000000000000000000000000000000000000000000000000001000;
		6'd4    :   out_sel = 64'b0000000000000000000000000000000000000000000000000000000000010000;
		6'd5    :   out_sel = 64'b0000000000000000000000000000000000000000000000000000000000100000;
		6'd6    :   out_sel = 64'b0000000000000000000000000000000000000000000000000000000001000000;
		6'd7    :   out_sel = 64'b0000000000000000000000000000000000000000000000000000000010000000;
		6'd8    :   out_sel = 64'b0000000000000000000000000000000000000000000000000000000100000000;
		6'd9    :   out_sel = 64'b0000000000000000000000000000000000000000000000000000001000000000;
		6'd10    :   out_sel = 64'b0000000000000000000000000000000000000000000000000000010000000000;
		6'd11    :   out_sel = 64'b0000000000000000000000000000000000000000000000000000100000000000;
		6'd12    :   out_sel = 64'b0000000000000000000000000000000000000000000000000001000000000000;
		6'd13    :   out_sel = 64'b0000000000000000000000000000000000000000000000000010000000000000;
		6'd14    :   out_sel = 64'b0000000000000000000000000000000000000000000000000100000000000000;
		6'd15    :   out_sel = 64'b0000000000000000000000000000000000000000000000001000000000000000;
		6'd16    :   out_sel = 64'b0000000000000000000000000000000000000000000000010000000000000000;
		6'd17    :   out_sel = 64'b0000000000000000000000000000000000000000000000100000000000000000;
		6'd18    :   out_sel = 64'b0000000000000000000000000000000000000000000001000000000000000000;
		6'd19    :   out_sel = 64'b0000000000000000000000000000000000000000000010000000000000000000;
		6'd20    :   out_sel = 64'b0000000000000000000000000000000000000000000100000000000000000000;
		6'd21    :   out_sel = 64'b0000000000000000000000000000000000000000001000000000000000000000;
		6'd22    :   out_sel = 64'b0000000000000000000000000000000000000000010000000000000000000000;
		6'd23    :   out_sel = 64'b0000000000000000000000000000000000000000100000000000000000000000;
		6'd24    :   out_sel = 64'b0000000000000000000000000000000000000001000000000000000000000000;
		6'd25    :   out_sel = 64'b0000000000000000000000000000000000000010000000000000000000000000;
		6'd26    :   out_sel = 64'b0000000000000000000000000000000000000100000000000000000000000000;
		6'd27    :   out_sel = 64'b0000000000000000000000000000000000001000000000000000000000000000;
		6'd28    :   out_sel = 64'b0000000000000000000000000000000000010000000000000000000000000000;
		6'd29    :   out_sel = 64'b0000000000000000000000000000000000100000000000000000000000000000;
		6'd30    :   out_sel = 64'b0000000000000000000000000000000001000000000000000000000000000000;
		6'd31    :   out_sel = 64'b0000000000000000000000000000000010000000000000000000000000000000;
		6'd32    :   out_sel = 64'b0000000000000000000000000000000100000000000000000000000000000000;
		6'd33    :   out_sel = 64'b0000000000000000000000000000001000000000000000000000000000000000;
		6'd34    :   out_sel = 64'b0000000000000000000000000000010000000000000000000000000000000000;
		6'd35    :   out_sel = 64'b0000000000000000000000000000100000000000000000000000000000000000;
		6'd36    :   out_sel = 64'b0000000000000000000000000001000000000000000000000000000000000000;
		6'd37    :   out_sel = 64'b0000000000000000000000000010000000000000000000000000000000000000;
		6'd38    :   out_sel = 64'b0000000000000000000000000100000000000000000000000000000000000000;
		6'd39    :   out_sel = 64'b0000000000000000000000001000000000000000000000000000000000000000;
		6'd40    :   out_sel = 64'b0000000000000000000000010000000000000000000000000000000000000000;
		6'd41    :   out_sel = 64'b0000000000000000000000100000000000000000000000000000000000000000;
		6'd42    :   out_sel = 64'b0000000000000000000001000000000000000000000000000000000000000000;
		6'd43    :   out_sel = 64'b0000000000000000000010000000000000000000000000000000000000000000;
		6'd44    :   out_sel = 64'b0000000000000000000100000000000000000000000000000000000000000000;
		6'd45    :   out_sel = 64'b0000000000000000001000000000000000000000000000000000000000000000;
		6'd46    :   out_sel = 64'b0000000000000000010000000000000000000000000000000000000000000000;
		default :   out_sel = 64'b0;
	endcase 
end 

endmodule 

module mux_logic_32_47 ( 
	input logic  [63 : 0] out_sel,
	input logic  [31 : 0] I0, 
	input logic  [31 : 0] I1, 
	input logic  [31 : 0] I2, 
	input logic  [31 : 0] I3, 
	input logic  [31 : 0] I4, 
	input logic  [31 : 0] I5, 
	input logic  [31 : 0] I6, 
	input logic  [31 : 0] I7, 
	input logic  [31 : 0] I8, 
	input logic  [31 : 0] I9, 
	input logic  [31 : 0] I10, 
	input logic  [31 : 0] I11, 
	input logic  [31 : 0] I12, 
	input logic  [31 : 0] I13, 
	input logic  [31 : 0] I14, 
	input logic  [31 : 0] I15, 
	input logic  [31 : 0] I16, 
	input logic  [31 : 0] I17, 
	input logic  [31 : 0] I18, 
	input logic  [31 : 0] I19, 
	input logic  [31 : 0] I20, 
	input logic  [31 : 0] I21, 
	input logic  [31 : 0] I22, 
	input logic  [31 : 0] I23, 
	input logic  [31 : 0] I24, 
	input logic  [31 : 0] I25, 
	input logic  [31 : 0] I26, 
	input logic  [31 : 0] I27, 
	input logic  [31 : 0] I28, 
	input logic  [31 : 0] I29, 
	input logic  [31 : 0] I30, 
	input logic  [31 : 0] I31, 
	input logic  [31 : 0] I32, 
	input logic  [31 : 0] I33, 
	input logic  [31 : 0] I34, 
	input logic  [31 : 0] I35, 
	input logic  [31 : 0] I36, 
	input logic  [31 : 0] I37, 
	input logic  [31 : 0] I38, 
	input logic  [31 : 0] I39, 
	input logic  [31 : 0] I40, 
	input logic  [31 : 0] I41, 
	input logic  [31 : 0] I42, 
	input logic  [31 : 0] I43, 
	input logic  [31 : 0] I44, 
	input logic  [31 : 0] I45, 
	input logic  [31 : 0] I46, 
	output logic  [31 : 0] O0, 
	output logic  [31 : 0] O1, 
	output logic  [31 : 0] O2, 
	output logic  [31 : 0] O3, 
	output logic  [31 : 0] O4, 
	output logic  [31 : 0] O5, 
	output logic  [31 : 0] O6, 
	output logic  [31 : 0] O7, 
	output logic  [31 : 0] O8, 
	output logic  [31 : 0] O9, 
	output logic  [31 : 0] O10, 
	output logic  [31 : 0] O11, 
	output logic  [31 : 0] O12, 
	output logic  [31 : 0] O13, 
	output logic  [31 : 0] O14, 
	output logic  [31 : 0] O15, 
	output logic  [31 : 0] O16, 
	output logic  [31 : 0] O17, 
	output logic  [31 : 0] O18, 
	output logic  [31 : 0] O19, 
	output logic  [31 : 0] O20, 
	output logic  [31 : 0] O21, 
	output logic  [31 : 0] O22, 
	output logic  [31 : 0] O23); 
	AO_CELL inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	AO_CELL inst_1_0 ( 
	.A1(out_sel[2]), 
	.A2(I2[0]), 
	.B1(out_sel[3]), 
	.B2(I3[0]), 
	.Z(O1[0])); 
	AO_CELL inst_2_0 ( 
	.A1(out_sel[4]), 
	.A2(I4[0]), 
	.B1(out_sel[5]), 
	.B2(I5[0]), 
	.Z(O2[0])); 
	AO_CELL inst_3_0 ( 
	.A1(out_sel[6]), 
	.A2(I6[0]), 
	.B1(out_sel[7]), 
	.B2(I7[0]), 
	.Z(O3[0])); 
	AO_CELL inst_4_0 ( 
	.A1(out_sel[8]), 
	.A2(I8[0]), 
	.B1(out_sel[9]), 
	.B2(I9[0]), 
	.Z(O4[0])); 
	AO_CELL inst_5_0 ( 
	.A1(out_sel[10]), 
	.A2(I10[0]), 
	.B1(out_sel[11]), 
	.B2(I11[0]), 
	.Z(O5[0])); 
	AO_CELL inst_6_0 ( 
	.A1(out_sel[12]), 
	.A2(I12[0]), 
	.B1(out_sel[13]), 
	.B2(I13[0]), 
	.Z(O6[0])); 
	AO_CELL inst_7_0 ( 
	.A1(out_sel[14]), 
	.A2(I14[0]), 
	.B1(out_sel[15]), 
	.B2(I15[0]), 
	.Z(O7[0])); 
	AO_CELL inst_8_0 ( 
	.A1(out_sel[16]), 
	.A2(I16[0]), 
	.B1(out_sel[17]), 
	.B2(I17[0]), 
	.Z(O8[0])); 
	AO_CELL inst_9_0 ( 
	.A1(out_sel[18]), 
	.A2(I18[0]), 
	.B1(out_sel[19]), 
	.B2(I19[0]), 
	.Z(O9[0])); 
	AO_CELL inst_10_0 ( 
	.A1(out_sel[20]), 
	.A2(I20[0]), 
	.B1(out_sel[21]), 
	.B2(I21[0]), 
	.Z(O10[0])); 
	AO_CELL inst_11_0 ( 
	.A1(out_sel[22]), 
	.A2(I22[0]), 
	.B1(out_sel[23]), 
	.B2(I23[0]), 
	.Z(O11[0])); 
	AO_CELL inst_12_0 ( 
	.A1(out_sel[24]), 
	.A2(I24[0]), 
	.B1(out_sel[25]), 
	.B2(I25[0]), 
	.Z(O12[0])); 
	AO_CELL inst_13_0 ( 
	.A1(out_sel[26]), 
	.A2(I26[0]), 
	.B1(out_sel[27]), 
	.B2(I27[0]), 
	.Z(O13[0])); 
	AO_CELL inst_14_0 ( 
	.A1(out_sel[28]), 
	.A2(I28[0]), 
	.B1(out_sel[29]), 
	.B2(I29[0]), 
	.Z(O14[0])); 
	AO_CELL inst_15_0 ( 
	.A1(out_sel[30]), 
	.A2(I30[0]), 
	.B1(out_sel[31]), 
	.B2(I31[0]), 
	.Z(O15[0])); 
	AO_CELL inst_16_0 ( 
	.A1(out_sel[32]), 
	.A2(I32[0]), 
	.B1(out_sel[33]), 
	.B2(I33[0]), 
	.Z(O16[0])); 
	AO_CELL inst_17_0 ( 
	.A1(out_sel[34]), 
	.A2(I34[0]), 
	.B1(out_sel[35]), 
	.B2(I35[0]), 
	.Z(O17[0])); 
	AO_CELL inst_18_0 ( 
	.A1(out_sel[36]), 
	.A2(I36[0]), 
	.B1(out_sel[37]), 
	.B2(I37[0]), 
	.Z(O18[0])); 
	AO_CELL inst_19_0 ( 
	.A1(out_sel[38]), 
	.A2(I38[0]), 
	.B1(out_sel[39]), 
	.B2(I39[0]), 
	.Z(O19[0])); 
	AO_CELL inst_20_0 ( 
	.A1(out_sel[40]), 
	.A2(I40[0]), 
	.B1(out_sel[41]), 
	.B2(I41[0]), 
	.Z(O20[0])); 
	AO_CELL inst_21_0 ( 
	.A1(out_sel[42]), 
	.A2(I42[0]), 
	.B1(out_sel[43]), 
	.B2(I43[0]), 
	.Z(O21[0])); 
	AO_CELL inst_22_0 ( 
	.A1(out_sel[44]), 
	.A2(I44[0]), 
	.B1(out_sel[45]), 
	.B2(I45[0]), 
	.Z(O22[0])); 
	AN_CELL inst_and_0 ( 
	.A1(out_sel[46]), 
	.A2(I46[0]), 
	.Z(O23[0])); 
	AO_CELL inst_0_1 ( 
	.A1(out_sel[0]), 
	.A2(I0[1]), 
	.B1(out_sel[1]), 
	.B2(I1[1]), 
	.Z(O0[1])); 
	AO_CELL inst_1_1 ( 
	.A1(out_sel[2]), 
	.A2(I2[1]), 
	.B1(out_sel[3]), 
	.B2(I3[1]), 
	.Z(O1[1])); 
	AO_CELL inst_2_1 ( 
	.A1(out_sel[4]), 
	.A2(I4[1]), 
	.B1(out_sel[5]), 
	.B2(I5[1]), 
	.Z(O2[1])); 
	AO_CELL inst_3_1 ( 
	.A1(out_sel[6]), 
	.A2(I6[1]), 
	.B1(out_sel[7]), 
	.B2(I7[1]), 
	.Z(O3[1])); 
	AO_CELL inst_4_1 ( 
	.A1(out_sel[8]), 
	.A2(I8[1]), 
	.B1(out_sel[9]), 
	.B2(I9[1]), 
	.Z(O4[1])); 
	AO_CELL inst_5_1 ( 
	.A1(out_sel[10]), 
	.A2(I10[1]), 
	.B1(out_sel[11]), 
	.B2(I11[1]), 
	.Z(O5[1])); 
	AO_CELL inst_6_1 ( 
	.A1(out_sel[12]), 
	.A2(I12[1]), 
	.B1(out_sel[13]), 
	.B2(I13[1]), 
	.Z(O6[1])); 
	AO_CELL inst_7_1 ( 
	.A1(out_sel[14]), 
	.A2(I14[1]), 
	.B1(out_sel[15]), 
	.B2(I15[1]), 
	.Z(O7[1])); 
	AO_CELL inst_8_1 ( 
	.A1(out_sel[16]), 
	.A2(I16[1]), 
	.B1(out_sel[17]), 
	.B2(I17[1]), 
	.Z(O8[1])); 
	AO_CELL inst_9_1 ( 
	.A1(out_sel[18]), 
	.A2(I18[1]), 
	.B1(out_sel[19]), 
	.B2(I19[1]), 
	.Z(O9[1])); 
	AO_CELL inst_10_1 ( 
	.A1(out_sel[20]), 
	.A2(I20[1]), 
	.B1(out_sel[21]), 
	.B2(I21[1]), 
	.Z(O10[1])); 
	AO_CELL inst_11_1 ( 
	.A1(out_sel[22]), 
	.A2(I22[1]), 
	.B1(out_sel[23]), 
	.B2(I23[1]), 
	.Z(O11[1])); 
	AO_CELL inst_12_1 ( 
	.A1(out_sel[24]), 
	.A2(I24[1]), 
	.B1(out_sel[25]), 
	.B2(I25[1]), 
	.Z(O12[1])); 
	AO_CELL inst_13_1 ( 
	.A1(out_sel[26]), 
	.A2(I26[1]), 
	.B1(out_sel[27]), 
	.B2(I27[1]), 
	.Z(O13[1])); 
	AO_CELL inst_14_1 ( 
	.A1(out_sel[28]), 
	.A2(I28[1]), 
	.B1(out_sel[29]), 
	.B2(I29[1]), 
	.Z(O14[1])); 
	AO_CELL inst_15_1 ( 
	.A1(out_sel[30]), 
	.A2(I30[1]), 
	.B1(out_sel[31]), 
	.B2(I31[1]), 
	.Z(O15[1])); 
	AO_CELL inst_16_1 ( 
	.A1(out_sel[32]), 
	.A2(I32[1]), 
	.B1(out_sel[33]), 
	.B2(I33[1]), 
	.Z(O16[1])); 
	AO_CELL inst_17_1 ( 
	.A1(out_sel[34]), 
	.A2(I34[1]), 
	.B1(out_sel[35]), 
	.B2(I35[1]), 
	.Z(O17[1])); 
	AO_CELL inst_18_1 ( 
	.A1(out_sel[36]), 
	.A2(I36[1]), 
	.B1(out_sel[37]), 
	.B2(I37[1]), 
	.Z(O18[1])); 
	AO_CELL inst_19_1 ( 
	.A1(out_sel[38]), 
	.A2(I38[1]), 
	.B1(out_sel[39]), 
	.B2(I39[1]), 
	.Z(O19[1])); 
	AO_CELL inst_20_1 ( 
	.A1(out_sel[40]), 
	.A2(I40[1]), 
	.B1(out_sel[41]), 
	.B2(I41[1]), 
	.Z(O20[1])); 
	AO_CELL inst_21_1 ( 
	.A1(out_sel[42]), 
	.A2(I42[1]), 
	.B1(out_sel[43]), 
	.B2(I43[1]), 
	.Z(O21[1])); 
	AO_CELL inst_22_1 ( 
	.A1(out_sel[44]), 
	.A2(I44[1]), 
	.B1(out_sel[45]), 
	.B2(I45[1]), 
	.Z(O22[1])); 
	AN_CELL inst_and_1 ( 
	.A1(out_sel[46]), 
	.A2(I46[1]), 
	.Z(O23[1])); 
	AO_CELL inst_0_2 ( 
	.A1(out_sel[0]), 
	.A2(I0[2]), 
	.B1(out_sel[1]), 
	.B2(I1[2]), 
	.Z(O0[2])); 
	AO_CELL inst_1_2 ( 
	.A1(out_sel[2]), 
	.A2(I2[2]), 
	.B1(out_sel[3]), 
	.B2(I3[2]), 
	.Z(O1[2])); 
	AO_CELL inst_2_2 ( 
	.A1(out_sel[4]), 
	.A2(I4[2]), 
	.B1(out_sel[5]), 
	.B2(I5[2]), 
	.Z(O2[2])); 
	AO_CELL inst_3_2 ( 
	.A1(out_sel[6]), 
	.A2(I6[2]), 
	.B1(out_sel[7]), 
	.B2(I7[2]), 
	.Z(O3[2])); 
	AO_CELL inst_4_2 ( 
	.A1(out_sel[8]), 
	.A2(I8[2]), 
	.B1(out_sel[9]), 
	.B2(I9[2]), 
	.Z(O4[2])); 
	AO_CELL inst_5_2 ( 
	.A1(out_sel[10]), 
	.A2(I10[2]), 
	.B1(out_sel[11]), 
	.B2(I11[2]), 
	.Z(O5[2])); 
	AO_CELL inst_6_2 ( 
	.A1(out_sel[12]), 
	.A2(I12[2]), 
	.B1(out_sel[13]), 
	.B2(I13[2]), 
	.Z(O6[2])); 
	AO_CELL inst_7_2 ( 
	.A1(out_sel[14]), 
	.A2(I14[2]), 
	.B1(out_sel[15]), 
	.B2(I15[2]), 
	.Z(O7[2])); 
	AO_CELL inst_8_2 ( 
	.A1(out_sel[16]), 
	.A2(I16[2]), 
	.B1(out_sel[17]), 
	.B2(I17[2]), 
	.Z(O8[2])); 
	AO_CELL inst_9_2 ( 
	.A1(out_sel[18]), 
	.A2(I18[2]), 
	.B1(out_sel[19]), 
	.B2(I19[2]), 
	.Z(O9[2])); 
	AO_CELL inst_10_2 ( 
	.A1(out_sel[20]), 
	.A2(I20[2]), 
	.B1(out_sel[21]), 
	.B2(I21[2]), 
	.Z(O10[2])); 
	AO_CELL inst_11_2 ( 
	.A1(out_sel[22]), 
	.A2(I22[2]), 
	.B1(out_sel[23]), 
	.B2(I23[2]), 
	.Z(O11[2])); 
	AO_CELL inst_12_2 ( 
	.A1(out_sel[24]), 
	.A2(I24[2]), 
	.B1(out_sel[25]), 
	.B2(I25[2]), 
	.Z(O12[2])); 
	AO_CELL inst_13_2 ( 
	.A1(out_sel[26]), 
	.A2(I26[2]), 
	.B1(out_sel[27]), 
	.B2(I27[2]), 
	.Z(O13[2])); 
	AO_CELL inst_14_2 ( 
	.A1(out_sel[28]), 
	.A2(I28[2]), 
	.B1(out_sel[29]), 
	.B2(I29[2]), 
	.Z(O14[2])); 
	AO_CELL inst_15_2 ( 
	.A1(out_sel[30]), 
	.A2(I30[2]), 
	.B1(out_sel[31]), 
	.B2(I31[2]), 
	.Z(O15[2])); 
	AO_CELL inst_16_2 ( 
	.A1(out_sel[32]), 
	.A2(I32[2]), 
	.B1(out_sel[33]), 
	.B2(I33[2]), 
	.Z(O16[2])); 
	AO_CELL inst_17_2 ( 
	.A1(out_sel[34]), 
	.A2(I34[2]), 
	.B1(out_sel[35]), 
	.B2(I35[2]), 
	.Z(O17[2])); 
	AO_CELL inst_18_2 ( 
	.A1(out_sel[36]), 
	.A2(I36[2]), 
	.B1(out_sel[37]), 
	.B2(I37[2]), 
	.Z(O18[2])); 
	AO_CELL inst_19_2 ( 
	.A1(out_sel[38]), 
	.A2(I38[2]), 
	.B1(out_sel[39]), 
	.B2(I39[2]), 
	.Z(O19[2])); 
	AO_CELL inst_20_2 ( 
	.A1(out_sel[40]), 
	.A2(I40[2]), 
	.B1(out_sel[41]), 
	.B2(I41[2]), 
	.Z(O20[2])); 
	AO_CELL inst_21_2 ( 
	.A1(out_sel[42]), 
	.A2(I42[2]), 
	.B1(out_sel[43]), 
	.B2(I43[2]), 
	.Z(O21[2])); 
	AO_CELL inst_22_2 ( 
	.A1(out_sel[44]), 
	.A2(I44[2]), 
	.B1(out_sel[45]), 
	.B2(I45[2]), 
	.Z(O22[2])); 
	AN_CELL inst_and_2 ( 
	.A1(out_sel[46]), 
	.A2(I46[2]), 
	.Z(O23[2])); 
	AO_CELL inst_0_3 ( 
	.A1(out_sel[0]), 
	.A2(I0[3]), 
	.B1(out_sel[1]), 
	.B2(I1[3]), 
	.Z(O0[3])); 
	AO_CELL inst_1_3 ( 
	.A1(out_sel[2]), 
	.A2(I2[3]), 
	.B1(out_sel[3]), 
	.B2(I3[3]), 
	.Z(O1[3])); 
	AO_CELL inst_2_3 ( 
	.A1(out_sel[4]), 
	.A2(I4[3]), 
	.B1(out_sel[5]), 
	.B2(I5[3]), 
	.Z(O2[3])); 
	AO_CELL inst_3_3 ( 
	.A1(out_sel[6]), 
	.A2(I6[3]), 
	.B1(out_sel[7]), 
	.B2(I7[3]), 
	.Z(O3[3])); 
	AO_CELL inst_4_3 ( 
	.A1(out_sel[8]), 
	.A2(I8[3]), 
	.B1(out_sel[9]), 
	.B2(I9[3]), 
	.Z(O4[3])); 
	AO_CELL inst_5_3 ( 
	.A1(out_sel[10]), 
	.A2(I10[3]), 
	.B1(out_sel[11]), 
	.B2(I11[3]), 
	.Z(O5[3])); 
	AO_CELL inst_6_3 ( 
	.A1(out_sel[12]), 
	.A2(I12[3]), 
	.B1(out_sel[13]), 
	.B2(I13[3]), 
	.Z(O6[3])); 
	AO_CELL inst_7_3 ( 
	.A1(out_sel[14]), 
	.A2(I14[3]), 
	.B1(out_sel[15]), 
	.B2(I15[3]), 
	.Z(O7[3])); 
	AO_CELL inst_8_3 ( 
	.A1(out_sel[16]), 
	.A2(I16[3]), 
	.B1(out_sel[17]), 
	.B2(I17[3]), 
	.Z(O8[3])); 
	AO_CELL inst_9_3 ( 
	.A1(out_sel[18]), 
	.A2(I18[3]), 
	.B1(out_sel[19]), 
	.B2(I19[3]), 
	.Z(O9[3])); 
	AO_CELL inst_10_3 ( 
	.A1(out_sel[20]), 
	.A2(I20[3]), 
	.B1(out_sel[21]), 
	.B2(I21[3]), 
	.Z(O10[3])); 
	AO_CELL inst_11_3 ( 
	.A1(out_sel[22]), 
	.A2(I22[3]), 
	.B1(out_sel[23]), 
	.B2(I23[3]), 
	.Z(O11[3])); 
	AO_CELL inst_12_3 ( 
	.A1(out_sel[24]), 
	.A2(I24[3]), 
	.B1(out_sel[25]), 
	.B2(I25[3]), 
	.Z(O12[3])); 
	AO_CELL inst_13_3 ( 
	.A1(out_sel[26]), 
	.A2(I26[3]), 
	.B1(out_sel[27]), 
	.B2(I27[3]), 
	.Z(O13[3])); 
	AO_CELL inst_14_3 ( 
	.A1(out_sel[28]), 
	.A2(I28[3]), 
	.B1(out_sel[29]), 
	.B2(I29[3]), 
	.Z(O14[3])); 
	AO_CELL inst_15_3 ( 
	.A1(out_sel[30]), 
	.A2(I30[3]), 
	.B1(out_sel[31]), 
	.B2(I31[3]), 
	.Z(O15[3])); 
	AO_CELL inst_16_3 ( 
	.A1(out_sel[32]), 
	.A2(I32[3]), 
	.B1(out_sel[33]), 
	.B2(I33[3]), 
	.Z(O16[3])); 
	AO_CELL inst_17_3 ( 
	.A1(out_sel[34]), 
	.A2(I34[3]), 
	.B1(out_sel[35]), 
	.B2(I35[3]), 
	.Z(O17[3])); 
	AO_CELL inst_18_3 ( 
	.A1(out_sel[36]), 
	.A2(I36[3]), 
	.B1(out_sel[37]), 
	.B2(I37[3]), 
	.Z(O18[3])); 
	AO_CELL inst_19_3 ( 
	.A1(out_sel[38]), 
	.A2(I38[3]), 
	.B1(out_sel[39]), 
	.B2(I39[3]), 
	.Z(O19[3])); 
	AO_CELL inst_20_3 ( 
	.A1(out_sel[40]), 
	.A2(I40[3]), 
	.B1(out_sel[41]), 
	.B2(I41[3]), 
	.Z(O20[3])); 
	AO_CELL inst_21_3 ( 
	.A1(out_sel[42]), 
	.A2(I42[3]), 
	.B1(out_sel[43]), 
	.B2(I43[3]), 
	.Z(O21[3])); 
	AO_CELL inst_22_3 ( 
	.A1(out_sel[44]), 
	.A2(I44[3]), 
	.B1(out_sel[45]), 
	.B2(I45[3]), 
	.Z(O22[3])); 
	AN_CELL inst_and_3 ( 
	.A1(out_sel[46]), 
	.A2(I46[3]), 
	.Z(O23[3])); 
	AO_CELL inst_0_4 ( 
	.A1(out_sel[0]), 
	.A2(I0[4]), 
	.B1(out_sel[1]), 
	.B2(I1[4]), 
	.Z(O0[4])); 
	AO_CELL inst_1_4 ( 
	.A1(out_sel[2]), 
	.A2(I2[4]), 
	.B1(out_sel[3]), 
	.B2(I3[4]), 
	.Z(O1[4])); 
	AO_CELL inst_2_4 ( 
	.A1(out_sel[4]), 
	.A2(I4[4]), 
	.B1(out_sel[5]), 
	.B2(I5[4]), 
	.Z(O2[4])); 
	AO_CELL inst_3_4 ( 
	.A1(out_sel[6]), 
	.A2(I6[4]), 
	.B1(out_sel[7]), 
	.B2(I7[4]), 
	.Z(O3[4])); 
	AO_CELL inst_4_4 ( 
	.A1(out_sel[8]), 
	.A2(I8[4]), 
	.B1(out_sel[9]), 
	.B2(I9[4]), 
	.Z(O4[4])); 
	AO_CELL inst_5_4 ( 
	.A1(out_sel[10]), 
	.A2(I10[4]), 
	.B1(out_sel[11]), 
	.B2(I11[4]), 
	.Z(O5[4])); 
	AO_CELL inst_6_4 ( 
	.A1(out_sel[12]), 
	.A2(I12[4]), 
	.B1(out_sel[13]), 
	.B2(I13[4]), 
	.Z(O6[4])); 
	AO_CELL inst_7_4 ( 
	.A1(out_sel[14]), 
	.A2(I14[4]), 
	.B1(out_sel[15]), 
	.B2(I15[4]), 
	.Z(O7[4])); 
	AO_CELL inst_8_4 ( 
	.A1(out_sel[16]), 
	.A2(I16[4]), 
	.B1(out_sel[17]), 
	.B2(I17[4]), 
	.Z(O8[4])); 
	AO_CELL inst_9_4 ( 
	.A1(out_sel[18]), 
	.A2(I18[4]), 
	.B1(out_sel[19]), 
	.B2(I19[4]), 
	.Z(O9[4])); 
	AO_CELL inst_10_4 ( 
	.A1(out_sel[20]), 
	.A2(I20[4]), 
	.B1(out_sel[21]), 
	.B2(I21[4]), 
	.Z(O10[4])); 
	AO_CELL inst_11_4 ( 
	.A1(out_sel[22]), 
	.A2(I22[4]), 
	.B1(out_sel[23]), 
	.B2(I23[4]), 
	.Z(O11[4])); 
	AO_CELL inst_12_4 ( 
	.A1(out_sel[24]), 
	.A2(I24[4]), 
	.B1(out_sel[25]), 
	.B2(I25[4]), 
	.Z(O12[4])); 
	AO_CELL inst_13_4 ( 
	.A1(out_sel[26]), 
	.A2(I26[4]), 
	.B1(out_sel[27]), 
	.B2(I27[4]), 
	.Z(O13[4])); 
	AO_CELL inst_14_4 ( 
	.A1(out_sel[28]), 
	.A2(I28[4]), 
	.B1(out_sel[29]), 
	.B2(I29[4]), 
	.Z(O14[4])); 
	AO_CELL inst_15_4 ( 
	.A1(out_sel[30]), 
	.A2(I30[4]), 
	.B1(out_sel[31]), 
	.B2(I31[4]), 
	.Z(O15[4])); 
	AO_CELL inst_16_4 ( 
	.A1(out_sel[32]), 
	.A2(I32[4]), 
	.B1(out_sel[33]), 
	.B2(I33[4]), 
	.Z(O16[4])); 
	AO_CELL inst_17_4 ( 
	.A1(out_sel[34]), 
	.A2(I34[4]), 
	.B1(out_sel[35]), 
	.B2(I35[4]), 
	.Z(O17[4])); 
	AO_CELL inst_18_4 ( 
	.A1(out_sel[36]), 
	.A2(I36[4]), 
	.B1(out_sel[37]), 
	.B2(I37[4]), 
	.Z(O18[4])); 
	AO_CELL inst_19_4 ( 
	.A1(out_sel[38]), 
	.A2(I38[4]), 
	.B1(out_sel[39]), 
	.B2(I39[4]), 
	.Z(O19[4])); 
	AO_CELL inst_20_4 ( 
	.A1(out_sel[40]), 
	.A2(I40[4]), 
	.B1(out_sel[41]), 
	.B2(I41[4]), 
	.Z(O20[4])); 
	AO_CELL inst_21_4 ( 
	.A1(out_sel[42]), 
	.A2(I42[4]), 
	.B1(out_sel[43]), 
	.B2(I43[4]), 
	.Z(O21[4])); 
	AO_CELL inst_22_4 ( 
	.A1(out_sel[44]), 
	.A2(I44[4]), 
	.B1(out_sel[45]), 
	.B2(I45[4]), 
	.Z(O22[4])); 
	AN_CELL inst_and_4 ( 
	.A1(out_sel[46]), 
	.A2(I46[4]), 
	.Z(O23[4])); 
	AO_CELL inst_0_5 ( 
	.A1(out_sel[0]), 
	.A2(I0[5]), 
	.B1(out_sel[1]), 
	.B2(I1[5]), 
	.Z(O0[5])); 
	AO_CELL inst_1_5 ( 
	.A1(out_sel[2]), 
	.A2(I2[5]), 
	.B1(out_sel[3]), 
	.B2(I3[5]), 
	.Z(O1[5])); 
	AO_CELL inst_2_5 ( 
	.A1(out_sel[4]), 
	.A2(I4[5]), 
	.B1(out_sel[5]), 
	.B2(I5[5]), 
	.Z(O2[5])); 
	AO_CELL inst_3_5 ( 
	.A1(out_sel[6]), 
	.A2(I6[5]), 
	.B1(out_sel[7]), 
	.B2(I7[5]), 
	.Z(O3[5])); 
	AO_CELL inst_4_5 ( 
	.A1(out_sel[8]), 
	.A2(I8[5]), 
	.B1(out_sel[9]), 
	.B2(I9[5]), 
	.Z(O4[5])); 
	AO_CELL inst_5_5 ( 
	.A1(out_sel[10]), 
	.A2(I10[5]), 
	.B1(out_sel[11]), 
	.B2(I11[5]), 
	.Z(O5[5])); 
	AO_CELL inst_6_5 ( 
	.A1(out_sel[12]), 
	.A2(I12[5]), 
	.B1(out_sel[13]), 
	.B2(I13[5]), 
	.Z(O6[5])); 
	AO_CELL inst_7_5 ( 
	.A1(out_sel[14]), 
	.A2(I14[5]), 
	.B1(out_sel[15]), 
	.B2(I15[5]), 
	.Z(O7[5])); 
	AO_CELL inst_8_5 ( 
	.A1(out_sel[16]), 
	.A2(I16[5]), 
	.B1(out_sel[17]), 
	.B2(I17[5]), 
	.Z(O8[5])); 
	AO_CELL inst_9_5 ( 
	.A1(out_sel[18]), 
	.A2(I18[5]), 
	.B1(out_sel[19]), 
	.B2(I19[5]), 
	.Z(O9[5])); 
	AO_CELL inst_10_5 ( 
	.A1(out_sel[20]), 
	.A2(I20[5]), 
	.B1(out_sel[21]), 
	.B2(I21[5]), 
	.Z(O10[5])); 
	AO_CELL inst_11_5 ( 
	.A1(out_sel[22]), 
	.A2(I22[5]), 
	.B1(out_sel[23]), 
	.B2(I23[5]), 
	.Z(O11[5])); 
	AO_CELL inst_12_5 ( 
	.A1(out_sel[24]), 
	.A2(I24[5]), 
	.B1(out_sel[25]), 
	.B2(I25[5]), 
	.Z(O12[5])); 
	AO_CELL inst_13_5 ( 
	.A1(out_sel[26]), 
	.A2(I26[5]), 
	.B1(out_sel[27]), 
	.B2(I27[5]), 
	.Z(O13[5])); 
	AO_CELL inst_14_5 ( 
	.A1(out_sel[28]), 
	.A2(I28[5]), 
	.B1(out_sel[29]), 
	.B2(I29[5]), 
	.Z(O14[5])); 
	AO_CELL inst_15_5 ( 
	.A1(out_sel[30]), 
	.A2(I30[5]), 
	.B1(out_sel[31]), 
	.B2(I31[5]), 
	.Z(O15[5])); 
	AO_CELL inst_16_5 ( 
	.A1(out_sel[32]), 
	.A2(I32[5]), 
	.B1(out_sel[33]), 
	.B2(I33[5]), 
	.Z(O16[5])); 
	AO_CELL inst_17_5 ( 
	.A1(out_sel[34]), 
	.A2(I34[5]), 
	.B1(out_sel[35]), 
	.B2(I35[5]), 
	.Z(O17[5])); 
	AO_CELL inst_18_5 ( 
	.A1(out_sel[36]), 
	.A2(I36[5]), 
	.B1(out_sel[37]), 
	.B2(I37[5]), 
	.Z(O18[5])); 
	AO_CELL inst_19_5 ( 
	.A1(out_sel[38]), 
	.A2(I38[5]), 
	.B1(out_sel[39]), 
	.B2(I39[5]), 
	.Z(O19[5])); 
	AO_CELL inst_20_5 ( 
	.A1(out_sel[40]), 
	.A2(I40[5]), 
	.B1(out_sel[41]), 
	.B2(I41[5]), 
	.Z(O20[5])); 
	AO_CELL inst_21_5 ( 
	.A1(out_sel[42]), 
	.A2(I42[5]), 
	.B1(out_sel[43]), 
	.B2(I43[5]), 
	.Z(O21[5])); 
	AO_CELL inst_22_5 ( 
	.A1(out_sel[44]), 
	.A2(I44[5]), 
	.B1(out_sel[45]), 
	.B2(I45[5]), 
	.Z(O22[5])); 
	AN_CELL inst_and_5 ( 
	.A1(out_sel[46]), 
	.A2(I46[5]), 
	.Z(O23[5])); 
	AO_CELL inst_0_6 ( 
	.A1(out_sel[0]), 
	.A2(I0[6]), 
	.B1(out_sel[1]), 
	.B2(I1[6]), 
	.Z(O0[6])); 
	AO_CELL inst_1_6 ( 
	.A1(out_sel[2]), 
	.A2(I2[6]), 
	.B1(out_sel[3]), 
	.B2(I3[6]), 
	.Z(O1[6])); 
	AO_CELL inst_2_6 ( 
	.A1(out_sel[4]), 
	.A2(I4[6]), 
	.B1(out_sel[5]), 
	.B2(I5[6]), 
	.Z(O2[6])); 
	AO_CELL inst_3_6 ( 
	.A1(out_sel[6]), 
	.A2(I6[6]), 
	.B1(out_sel[7]), 
	.B2(I7[6]), 
	.Z(O3[6])); 
	AO_CELL inst_4_6 ( 
	.A1(out_sel[8]), 
	.A2(I8[6]), 
	.B1(out_sel[9]), 
	.B2(I9[6]), 
	.Z(O4[6])); 
	AO_CELL inst_5_6 ( 
	.A1(out_sel[10]), 
	.A2(I10[6]), 
	.B1(out_sel[11]), 
	.B2(I11[6]), 
	.Z(O5[6])); 
	AO_CELL inst_6_6 ( 
	.A1(out_sel[12]), 
	.A2(I12[6]), 
	.B1(out_sel[13]), 
	.B2(I13[6]), 
	.Z(O6[6])); 
	AO_CELL inst_7_6 ( 
	.A1(out_sel[14]), 
	.A2(I14[6]), 
	.B1(out_sel[15]), 
	.B2(I15[6]), 
	.Z(O7[6])); 
	AO_CELL inst_8_6 ( 
	.A1(out_sel[16]), 
	.A2(I16[6]), 
	.B1(out_sel[17]), 
	.B2(I17[6]), 
	.Z(O8[6])); 
	AO_CELL inst_9_6 ( 
	.A1(out_sel[18]), 
	.A2(I18[6]), 
	.B1(out_sel[19]), 
	.B2(I19[6]), 
	.Z(O9[6])); 
	AO_CELL inst_10_6 ( 
	.A1(out_sel[20]), 
	.A2(I20[6]), 
	.B1(out_sel[21]), 
	.B2(I21[6]), 
	.Z(O10[6])); 
	AO_CELL inst_11_6 ( 
	.A1(out_sel[22]), 
	.A2(I22[6]), 
	.B1(out_sel[23]), 
	.B2(I23[6]), 
	.Z(O11[6])); 
	AO_CELL inst_12_6 ( 
	.A1(out_sel[24]), 
	.A2(I24[6]), 
	.B1(out_sel[25]), 
	.B2(I25[6]), 
	.Z(O12[6])); 
	AO_CELL inst_13_6 ( 
	.A1(out_sel[26]), 
	.A2(I26[6]), 
	.B1(out_sel[27]), 
	.B2(I27[6]), 
	.Z(O13[6])); 
	AO_CELL inst_14_6 ( 
	.A1(out_sel[28]), 
	.A2(I28[6]), 
	.B1(out_sel[29]), 
	.B2(I29[6]), 
	.Z(O14[6])); 
	AO_CELL inst_15_6 ( 
	.A1(out_sel[30]), 
	.A2(I30[6]), 
	.B1(out_sel[31]), 
	.B2(I31[6]), 
	.Z(O15[6])); 
	AO_CELL inst_16_6 ( 
	.A1(out_sel[32]), 
	.A2(I32[6]), 
	.B1(out_sel[33]), 
	.B2(I33[6]), 
	.Z(O16[6])); 
	AO_CELL inst_17_6 ( 
	.A1(out_sel[34]), 
	.A2(I34[6]), 
	.B1(out_sel[35]), 
	.B2(I35[6]), 
	.Z(O17[6])); 
	AO_CELL inst_18_6 ( 
	.A1(out_sel[36]), 
	.A2(I36[6]), 
	.B1(out_sel[37]), 
	.B2(I37[6]), 
	.Z(O18[6])); 
	AO_CELL inst_19_6 ( 
	.A1(out_sel[38]), 
	.A2(I38[6]), 
	.B1(out_sel[39]), 
	.B2(I39[6]), 
	.Z(O19[6])); 
	AO_CELL inst_20_6 ( 
	.A1(out_sel[40]), 
	.A2(I40[6]), 
	.B1(out_sel[41]), 
	.B2(I41[6]), 
	.Z(O20[6])); 
	AO_CELL inst_21_6 ( 
	.A1(out_sel[42]), 
	.A2(I42[6]), 
	.B1(out_sel[43]), 
	.B2(I43[6]), 
	.Z(O21[6])); 
	AO_CELL inst_22_6 ( 
	.A1(out_sel[44]), 
	.A2(I44[6]), 
	.B1(out_sel[45]), 
	.B2(I45[6]), 
	.Z(O22[6])); 
	AN_CELL inst_and_6 ( 
	.A1(out_sel[46]), 
	.A2(I46[6]), 
	.Z(O23[6])); 
	AO_CELL inst_0_7 ( 
	.A1(out_sel[0]), 
	.A2(I0[7]), 
	.B1(out_sel[1]), 
	.B2(I1[7]), 
	.Z(O0[7])); 
	AO_CELL inst_1_7 ( 
	.A1(out_sel[2]), 
	.A2(I2[7]), 
	.B1(out_sel[3]), 
	.B2(I3[7]), 
	.Z(O1[7])); 
	AO_CELL inst_2_7 ( 
	.A1(out_sel[4]), 
	.A2(I4[7]), 
	.B1(out_sel[5]), 
	.B2(I5[7]), 
	.Z(O2[7])); 
	AO_CELL inst_3_7 ( 
	.A1(out_sel[6]), 
	.A2(I6[7]), 
	.B1(out_sel[7]), 
	.B2(I7[7]), 
	.Z(O3[7])); 
	AO_CELL inst_4_7 ( 
	.A1(out_sel[8]), 
	.A2(I8[7]), 
	.B1(out_sel[9]), 
	.B2(I9[7]), 
	.Z(O4[7])); 
	AO_CELL inst_5_7 ( 
	.A1(out_sel[10]), 
	.A2(I10[7]), 
	.B1(out_sel[11]), 
	.B2(I11[7]), 
	.Z(O5[7])); 
	AO_CELL inst_6_7 ( 
	.A1(out_sel[12]), 
	.A2(I12[7]), 
	.B1(out_sel[13]), 
	.B2(I13[7]), 
	.Z(O6[7])); 
	AO_CELL inst_7_7 ( 
	.A1(out_sel[14]), 
	.A2(I14[7]), 
	.B1(out_sel[15]), 
	.B2(I15[7]), 
	.Z(O7[7])); 
	AO_CELL inst_8_7 ( 
	.A1(out_sel[16]), 
	.A2(I16[7]), 
	.B1(out_sel[17]), 
	.B2(I17[7]), 
	.Z(O8[7])); 
	AO_CELL inst_9_7 ( 
	.A1(out_sel[18]), 
	.A2(I18[7]), 
	.B1(out_sel[19]), 
	.B2(I19[7]), 
	.Z(O9[7])); 
	AO_CELL inst_10_7 ( 
	.A1(out_sel[20]), 
	.A2(I20[7]), 
	.B1(out_sel[21]), 
	.B2(I21[7]), 
	.Z(O10[7])); 
	AO_CELL inst_11_7 ( 
	.A1(out_sel[22]), 
	.A2(I22[7]), 
	.B1(out_sel[23]), 
	.B2(I23[7]), 
	.Z(O11[7])); 
	AO_CELL inst_12_7 ( 
	.A1(out_sel[24]), 
	.A2(I24[7]), 
	.B1(out_sel[25]), 
	.B2(I25[7]), 
	.Z(O12[7])); 
	AO_CELL inst_13_7 ( 
	.A1(out_sel[26]), 
	.A2(I26[7]), 
	.B1(out_sel[27]), 
	.B2(I27[7]), 
	.Z(O13[7])); 
	AO_CELL inst_14_7 ( 
	.A1(out_sel[28]), 
	.A2(I28[7]), 
	.B1(out_sel[29]), 
	.B2(I29[7]), 
	.Z(O14[7])); 
	AO_CELL inst_15_7 ( 
	.A1(out_sel[30]), 
	.A2(I30[7]), 
	.B1(out_sel[31]), 
	.B2(I31[7]), 
	.Z(O15[7])); 
	AO_CELL inst_16_7 ( 
	.A1(out_sel[32]), 
	.A2(I32[7]), 
	.B1(out_sel[33]), 
	.B2(I33[7]), 
	.Z(O16[7])); 
	AO_CELL inst_17_7 ( 
	.A1(out_sel[34]), 
	.A2(I34[7]), 
	.B1(out_sel[35]), 
	.B2(I35[7]), 
	.Z(O17[7])); 
	AO_CELL inst_18_7 ( 
	.A1(out_sel[36]), 
	.A2(I36[7]), 
	.B1(out_sel[37]), 
	.B2(I37[7]), 
	.Z(O18[7])); 
	AO_CELL inst_19_7 ( 
	.A1(out_sel[38]), 
	.A2(I38[7]), 
	.B1(out_sel[39]), 
	.B2(I39[7]), 
	.Z(O19[7])); 
	AO_CELL inst_20_7 ( 
	.A1(out_sel[40]), 
	.A2(I40[7]), 
	.B1(out_sel[41]), 
	.B2(I41[7]), 
	.Z(O20[7])); 
	AO_CELL inst_21_7 ( 
	.A1(out_sel[42]), 
	.A2(I42[7]), 
	.B1(out_sel[43]), 
	.B2(I43[7]), 
	.Z(O21[7])); 
	AO_CELL inst_22_7 ( 
	.A1(out_sel[44]), 
	.A2(I44[7]), 
	.B1(out_sel[45]), 
	.B2(I45[7]), 
	.Z(O22[7])); 
	AN_CELL inst_and_7 ( 
	.A1(out_sel[46]), 
	.A2(I46[7]), 
	.Z(O23[7])); 
	AO_CELL inst_0_8 ( 
	.A1(out_sel[0]), 
	.A2(I0[8]), 
	.B1(out_sel[1]), 
	.B2(I1[8]), 
	.Z(O0[8])); 
	AO_CELL inst_1_8 ( 
	.A1(out_sel[2]), 
	.A2(I2[8]), 
	.B1(out_sel[3]), 
	.B2(I3[8]), 
	.Z(O1[8])); 
	AO_CELL inst_2_8 ( 
	.A1(out_sel[4]), 
	.A2(I4[8]), 
	.B1(out_sel[5]), 
	.B2(I5[8]), 
	.Z(O2[8])); 
	AO_CELL inst_3_8 ( 
	.A1(out_sel[6]), 
	.A2(I6[8]), 
	.B1(out_sel[7]), 
	.B2(I7[8]), 
	.Z(O3[8])); 
	AO_CELL inst_4_8 ( 
	.A1(out_sel[8]), 
	.A2(I8[8]), 
	.B1(out_sel[9]), 
	.B2(I9[8]), 
	.Z(O4[8])); 
	AO_CELL inst_5_8 ( 
	.A1(out_sel[10]), 
	.A2(I10[8]), 
	.B1(out_sel[11]), 
	.B2(I11[8]), 
	.Z(O5[8])); 
	AO_CELL inst_6_8 ( 
	.A1(out_sel[12]), 
	.A2(I12[8]), 
	.B1(out_sel[13]), 
	.B2(I13[8]), 
	.Z(O6[8])); 
	AO_CELL inst_7_8 ( 
	.A1(out_sel[14]), 
	.A2(I14[8]), 
	.B1(out_sel[15]), 
	.B2(I15[8]), 
	.Z(O7[8])); 
	AO_CELL inst_8_8 ( 
	.A1(out_sel[16]), 
	.A2(I16[8]), 
	.B1(out_sel[17]), 
	.B2(I17[8]), 
	.Z(O8[8])); 
	AO_CELL inst_9_8 ( 
	.A1(out_sel[18]), 
	.A2(I18[8]), 
	.B1(out_sel[19]), 
	.B2(I19[8]), 
	.Z(O9[8])); 
	AO_CELL inst_10_8 ( 
	.A1(out_sel[20]), 
	.A2(I20[8]), 
	.B1(out_sel[21]), 
	.B2(I21[8]), 
	.Z(O10[8])); 
	AO_CELL inst_11_8 ( 
	.A1(out_sel[22]), 
	.A2(I22[8]), 
	.B1(out_sel[23]), 
	.B2(I23[8]), 
	.Z(O11[8])); 
	AO_CELL inst_12_8 ( 
	.A1(out_sel[24]), 
	.A2(I24[8]), 
	.B1(out_sel[25]), 
	.B2(I25[8]), 
	.Z(O12[8])); 
	AO_CELL inst_13_8 ( 
	.A1(out_sel[26]), 
	.A2(I26[8]), 
	.B1(out_sel[27]), 
	.B2(I27[8]), 
	.Z(O13[8])); 
	AO_CELL inst_14_8 ( 
	.A1(out_sel[28]), 
	.A2(I28[8]), 
	.B1(out_sel[29]), 
	.B2(I29[8]), 
	.Z(O14[8])); 
	AO_CELL inst_15_8 ( 
	.A1(out_sel[30]), 
	.A2(I30[8]), 
	.B1(out_sel[31]), 
	.B2(I31[8]), 
	.Z(O15[8])); 
	AO_CELL inst_16_8 ( 
	.A1(out_sel[32]), 
	.A2(I32[8]), 
	.B1(out_sel[33]), 
	.B2(I33[8]), 
	.Z(O16[8])); 
	AO_CELL inst_17_8 ( 
	.A1(out_sel[34]), 
	.A2(I34[8]), 
	.B1(out_sel[35]), 
	.B2(I35[8]), 
	.Z(O17[8])); 
	AO_CELL inst_18_8 ( 
	.A1(out_sel[36]), 
	.A2(I36[8]), 
	.B1(out_sel[37]), 
	.B2(I37[8]), 
	.Z(O18[8])); 
	AO_CELL inst_19_8 ( 
	.A1(out_sel[38]), 
	.A2(I38[8]), 
	.B1(out_sel[39]), 
	.B2(I39[8]), 
	.Z(O19[8])); 
	AO_CELL inst_20_8 ( 
	.A1(out_sel[40]), 
	.A2(I40[8]), 
	.B1(out_sel[41]), 
	.B2(I41[8]), 
	.Z(O20[8])); 
	AO_CELL inst_21_8 ( 
	.A1(out_sel[42]), 
	.A2(I42[8]), 
	.B1(out_sel[43]), 
	.B2(I43[8]), 
	.Z(O21[8])); 
	AO_CELL inst_22_8 ( 
	.A1(out_sel[44]), 
	.A2(I44[8]), 
	.B1(out_sel[45]), 
	.B2(I45[8]), 
	.Z(O22[8])); 
	AN_CELL inst_and_8 ( 
	.A1(out_sel[46]), 
	.A2(I46[8]), 
	.Z(O23[8])); 
	AO_CELL inst_0_9 ( 
	.A1(out_sel[0]), 
	.A2(I0[9]), 
	.B1(out_sel[1]), 
	.B2(I1[9]), 
	.Z(O0[9])); 
	AO_CELL inst_1_9 ( 
	.A1(out_sel[2]), 
	.A2(I2[9]), 
	.B1(out_sel[3]), 
	.B2(I3[9]), 
	.Z(O1[9])); 
	AO_CELL inst_2_9 ( 
	.A1(out_sel[4]), 
	.A2(I4[9]), 
	.B1(out_sel[5]), 
	.B2(I5[9]), 
	.Z(O2[9])); 
	AO_CELL inst_3_9 ( 
	.A1(out_sel[6]), 
	.A2(I6[9]), 
	.B1(out_sel[7]), 
	.B2(I7[9]), 
	.Z(O3[9])); 
	AO_CELL inst_4_9 ( 
	.A1(out_sel[8]), 
	.A2(I8[9]), 
	.B1(out_sel[9]), 
	.B2(I9[9]), 
	.Z(O4[9])); 
	AO_CELL inst_5_9 ( 
	.A1(out_sel[10]), 
	.A2(I10[9]), 
	.B1(out_sel[11]), 
	.B2(I11[9]), 
	.Z(O5[9])); 
	AO_CELL inst_6_9 ( 
	.A1(out_sel[12]), 
	.A2(I12[9]), 
	.B1(out_sel[13]), 
	.B2(I13[9]), 
	.Z(O6[9])); 
	AO_CELL inst_7_9 ( 
	.A1(out_sel[14]), 
	.A2(I14[9]), 
	.B1(out_sel[15]), 
	.B2(I15[9]), 
	.Z(O7[9])); 
	AO_CELL inst_8_9 ( 
	.A1(out_sel[16]), 
	.A2(I16[9]), 
	.B1(out_sel[17]), 
	.B2(I17[9]), 
	.Z(O8[9])); 
	AO_CELL inst_9_9 ( 
	.A1(out_sel[18]), 
	.A2(I18[9]), 
	.B1(out_sel[19]), 
	.B2(I19[9]), 
	.Z(O9[9])); 
	AO_CELL inst_10_9 ( 
	.A1(out_sel[20]), 
	.A2(I20[9]), 
	.B1(out_sel[21]), 
	.B2(I21[9]), 
	.Z(O10[9])); 
	AO_CELL inst_11_9 ( 
	.A1(out_sel[22]), 
	.A2(I22[9]), 
	.B1(out_sel[23]), 
	.B2(I23[9]), 
	.Z(O11[9])); 
	AO_CELL inst_12_9 ( 
	.A1(out_sel[24]), 
	.A2(I24[9]), 
	.B1(out_sel[25]), 
	.B2(I25[9]), 
	.Z(O12[9])); 
	AO_CELL inst_13_9 ( 
	.A1(out_sel[26]), 
	.A2(I26[9]), 
	.B1(out_sel[27]), 
	.B2(I27[9]), 
	.Z(O13[9])); 
	AO_CELL inst_14_9 ( 
	.A1(out_sel[28]), 
	.A2(I28[9]), 
	.B1(out_sel[29]), 
	.B2(I29[9]), 
	.Z(O14[9])); 
	AO_CELL inst_15_9 ( 
	.A1(out_sel[30]), 
	.A2(I30[9]), 
	.B1(out_sel[31]), 
	.B2(I31[9]), 
	.Z(O15[9])); 
	AO_CELL inst_16_9 ( 
	.A1(out_sel[32]), 
	.A2(I32[9]), 
	.B1(out_sel[33]), 
	.B2(I33[9]), 
	.Z(O16[9])); 
	AO_CELL inst_17_9 ( 
	.A1(out_sel[34]), 
	.A2(I34[9]), 
	.B1(out_sel[35]), 
	.B2(I35[9]), 
	.Z(O17[9])); 
	AO_CELL inst_18_9 ( 
	.A1(out_sel[36]), 
	.A2(I36[9]), 
	.B1(out_sel[37]), 
	.B2(I37[9]), 
	.Z(O18[9])); 
	AO_CELL inst_19_9 ( 
	.A1(out_sel[38]), 
	.A2(I38[9]), 
	.B1(out_sel[39]), 
	.B2(I39[9]), 
	.Z(O19[9])); 
	AO_CELL inst_20_9 ( 
	.A1(out_sel[40]), 
	.A2(I40[9]), 
	.B1(out_sel[41]), 
	.B2(I41[9]), 
	.Z(O20[9])); 
	AO_CELL inst_21_9 ( 
	.A1(out_sel[42]), 
	.A2(I42[9]), 
	.B1(out_sel[43]), 
	.B2(I43[9]), 
	.Z(O21[9])); 
	AO_CELL inst_22_9 ( 
	.A1(out_sel[44]), 
	.A2(I44[9]), 
	.B1(out_sel[45]), 
	.B2(I45[9]), 
	.Z(O22[9])); 
	AN_CELL inst_and_9 ( 
	.A1(out_sel[46]), 
	.A2(I46[9]), 
	.Z(O23[9])); 
	AO_CELL inst_0_10 ( 
	.A1(out_sel[0]), 
	.A2(I0[10]), 
	.B1(out_sel[1]), 
	.B2(I1[10]), 
	.Z(O0[10])); 
	AO_CELL inst_1_10 ( 
	.A1(out_sel[2]), 
	.A2(I2[10]), 
	.B1(out_sel[3]), 
	.B2(I3[10]), 
	.Z(O1[10])); 
	AO_CELL inst_2_10 ( 
	.A1(out_sel[4]), 
	.A2(I4[10]), 
	.B1(out_sel[5]), 
	.B2(I5[10]), 
	.Z(O2[10])); 
	AO_CELL inst_3_10 ( 
	.A1(out_sel[6]), 
	.A2(I6[10]), 
	.B1(out_sel[7]), 
	.B2(I7[10]), 
	.Z(O3[10])); 
	AO_CELL inst_4_10 ( 
	.A1(out_sel[8]), 
	.A2(I8[10]), 
	.B1(out_sel[9]), 
	.B2(I9[10]), 
	.Z(O4[10])); 
	AO_CELL inst_5_10 ( 
	.A1(out_sel[10]), 
	.A2(I10[10]), 
	.B1(out_sel[11]), 
	.B2(I11[10]), 
	.Z(O5[10])); 
	AO_CELL inst_6_10 ( 
	.A1(out_sel[12]), 
	.A2(I12[10]), 
	.B1(out_sel[13]), 
	.B2(I13[10]), 
	.Z(O6[10])); 
	AO_CELL inst_7_10 ( 
	.A1(out_sel[14]), 
	.A2(I14[10]), 
	.B1(out_sel[15]), 
	.B2(I15[10]), 
	.Z(O7[10])); 
	AO_CELL inst_8_10 ( 
	.A1(out_sel[16]), 
	.A2(I16[10]), 
	.B1(out_sel[17]), 
	.B2(I17[10]), 
	.Z(O8[10])); 
	AO_CELL inst_9_10 ( 
	.A1(out_sel[18]), 
	.A2(I18[10]), 
	.B1(out_sel[19]), 
	.B2(I19[10]), 
	.Z(O9[10])); 
	AO_CELL inst_10_10 ( 
	.A1(out_sel[20]), 
	.A2(I20[10]), 
	.B1(out_sel[21]), 
	.B2(I21[10]), 
	.Z(O10[10])); 
	AO_CELL inst_11_10 ( 
	.A1(out_sel[22]), 
	.A2(I22[10]), 
	.B1(out_sel[23]), 
	.B2(I23[10]), 
	.Z(O11[10])); 
	AO_CELL inst_12_10 ( 
	.A1(out_sel[24]), 
	.A2(I24[10]), 
	.B1(out_sel[25]), 
	.B2(I25[10]), 
	.Z(O12[10])); 
	AO_CELL inst_13_10 ( 
	.A1(out_sel[26]), 
	.A2(I26[10]), 
	.B1(out_sel[27]), 
	.B2(I27[10]), 
	.Z(O13[10])); 
	AO_CELL inst_14_10 ( 
	.A1(out_sel[28]), 
	.A2(I28[10]), 
	.B1(out_sel[29]), 
	.B2(I29[10]), 
	.Z(O14[10])); 
	AO_CELL inst_15_10 ( 
	.A1(out_sel[30]), 
	.A2(I30[10]), 
	.B1(out_sel[31]), 
	.B2(I31[10]), 
	.Z(O15[10])); 
	AO_CELL inst_16_10 ( 
	.A1(out_sel[32]), 
	.A2(I32[10]), 
	.B1(out_sel[33]), 
	.B2(I33[10]), 
	.Z(O16[10])); 
	AO_CELL inst_17_10 ( 
	.A1(out_sel[34]), 
	.A2(I34[10]), 
	.B1(out_sel[35]), 
	.B2(I35[10]), 
	.Z(O17[10])); 
	AO_CELL inst_18_10 ( 
	.A1(out_sel[36]), 
	.A2(I36[10]), 
	.B1(out_sel[37]), 
	.B2(I37[10]), 
	.Z(O18[10])); 
	AO_CELL inst_19_10 ( 
	.A1(out_sel[38]), 
	.A2(I38[10]), 
	.B1(out_sel[39]), 
	.B2(I39[10]), 
	.Z(O19[10])); 
	AO_CELL inst_20_10 ( 
	.A1(out_sel[40]), 
	.A2(I40[10]), 
	.B1(out_sel[41]), 
	.B2(I41[10]), 
	.Z(O20[10])); 
	AO_CELL inst_21_10 ( 
	.A1(out_sel[42]), 
	.A2(I42[10]), 
	.B1(out_sel[43]), 
	.B2(I43[10]), 
	.Z(O21[10])); 
	AO_CELL inst_22_10 ( 
	.A1(out_sel[44]), 
	.A2(I44[10]), 
	.B1(out_sel[45]), 
	.B2(I45[10]), 
	.Z(O22[10])); 
	AN_CELL inst_and_10 ( 
	.A1(out_sel[46]), 
	.A2(I46[10]), 
	.Z(O23[10])); 
	AO_CELL inst_0_11 ( 
	.A1(out_sel[0]), 
	.A2(I0[11]), 
	.B1(out_sel[1]), 
	.B2(I1[11]), 
	.Z(O0[11])); 
	AO_CELL inst_1_11 ( 
	.A1(out_sel[2]), 
	.A2(I2[11]), 
	.B1(out_sel[3]), 
	.B2(I3[11]), 
	.Z(O1[11])); 
	AO_CELL inst_2_11 ( 
	.A1(out_sel[4]), 
	.A2(I4[11]), 
	.B1(out_sel[5]), 
	.B2(I5[11]), 
	.Z(O2[11])); 
	AO_CELL inst_3_11 ( 
	.A1(out_sel[6]), 
	.A2(I6[11]), 
	.B1(out_sel[7]), 
	.B2(I7[11]), 
	.Z(O3[11])); 
	AO_CELL inst_4_11 ( 
	.A1(out_sel[8]), 
	.A2(I8[11]), 
	.B1(out_sel[9]), 
	.B2(I9[11]), 
	.Z(O4[11])); 
	AO_CELL inst_5_11 ( 
	.A1(out_sel[10]), 
	.A2(I10[11]), 
	.B1(out_sel[11]), 
	.B2(I11[11]), 
	.Z(O5[11])); 
	AO_CELL inst_6_11 ( 
	.A1(out_sel[12]), 
	.A2(I12[11]), 
	.B1(out_sel[13]), 
	.B2(I13[11]), 
	.Z(O6[11])); 
	AO_CELL inst_7_11 ( 
	.A1(out_sel[14]), 
	.A2(I14[11]), 
	.B1(out_sel[15]), 
	.B2(I15[11]), 
	.Z(O7[11])); 
	AO_CELL inst_8_11 ( 
	.A1(out_sel[16]), 
	.A2(I16[11]), 
	.B1(out_sel[17]), 
	.B2(I17[11]), 
	.Z(O8[11])); 
	AO_CELL inst_9_11 ( 
	.A1(out_sel[18]), 
	.A2(I18[11]), 
	.B1(out_sel[19]), 
	.B2(I19[11]), 
	.Z(O9[11])); 
	AO_CELL inst_10_11 ( 
	.A1(out_sel[20]), 
	.A2(I20[11]), 
	.B1(out_sel[21]), 
	.B2(I21[11]), 
	.Z(O10[11])); 
	AO_CELL inst_11_11 ( 
	.A1(out_sel[22]), 
	.A2(I22[11]), 
	.B1(out_sel[23]), 
	.B2(I23[11]), 
	.Z(O11[11])); 
	AO_CELL inst_12_11 ( 
	.A1(out_sel[24]), 
	.A2(I24[11]), 
	.B1(out_sel[25]), 
	.B2(I25[11]), 
	.Z(O12[11])); 
	AO_CELL inst_13_11 ( 
	.A1(out_sel[26]), 
	.A2(I26[11]), 
	.B1(out_sel[27]), 
	.B2(I27[11]), 
	.Z(O13[11])); 
	AO_CELL inst_14_11 ( 
	.A1(out_sel[28]), 
	.A2(I28[11]), 
	.B1(out_sel[29]), 
	.B2(I29[11]), 
	.Z(O14[11])); 
	AO_CELL inst_15_11 ( 
	.A1(out_sel[30]), 
	.A2(I30[11]), 
	.B1(out_sel[31]), 
	.B2(I31[11]), 
	.Z(O15[11])); 
	AO_CELL inst_16_11 ( 
	.A1(out_sel[32]), 
	.A2(I32[11]), 
	.B1(out_sel[33]), 
	.B2(I33[11]), 
	.Z(O16[11])); 
	AO_CELL inst_17_11 ( 
	.A1(out_sel[34]), 
	.A2(I34[11]), 
	.B1(out_sel[35]), 
	.B2(I35[11]), 
	.Z(O17[11])); 
	AO_CELL inst_18_11 ( 
	.A1(out_sel[36]), 
	.A2(I36[11]), 
	.B1(out_sel[37]), 
	.B2(I37[11]), 
	.Z(O18[11])); 
	AO_CELL inst_19_11 ( 
	.A1(out_sel[38]), 
	.A2(I38[11]), 
	.B1(out_sel[39]), 
	.B2(I39[11]), 
	.Z(O19[11])); 
	AO_CELL inst_20_11 ( 
	.A1(out_sel[40]), 
	.A2(I40[11]), 
	.B1(out_sel[41]), 
	.B2(I41[11]), 
	.Z(O20[11])); 
	AO_CELL inst_21_11 ( 
	.A1(out_sel[42]), 
	.A2(I42[11]), 
	.B1(out_sel[43]), 
	.B2(I43[11]), 
	.Z(O21[11])); 
	AO_CELL inst_22_11 ( 
	.A1(out_sel[44]), 
	.A2(I44[11]), 
	.B1(out_sel[45]), 
	.B2(I45[11]), 
	.Z(O22[11])); 
	AN_CELL inst_and_11 ( 
	.A1(out_sel[46]), 
	.A2(I46[11]), 
	.Z(O23[11])); 
	AO_CELL inst_0_12 ( 
	.A1(out_sel[0]), 
	.A2(I0[12]), 
	.B1(out_sel[1]), 
	.B2(I1[12]), 
	.Z(O0[12])); 
	AO_CELL inst_1_12 ( 
	.A1(out_sel[2]), 
	.A2(I2[12]), 
	.B1(out_sel[3]), 
	.B2(I3[12]), 
	.Z(O1[12])); 
	AO_CELL inst_2_12 ( 
	.A1(out_sel[4]), 
	.A2(I4[12]), 
	.B1(out_sel[5]), 
	.B2(I5[12]), 
	.Z(O2[12])); 
	AO_CELL inst_3_12 ( 
	.A1(out_sel[6]), 
	.A2(I6[12]), 
	.B1(out_sel[7]), 
	.B2(I7[12]), 
	.Z(O3[12])); 
	AO_CELL inst_4_12 ( 
	.A1(out_sel[8]), 
	.A2(I8[12]), 
	.B1(out_sel[9]), 
	.B2(I9[12]), 
	.Z(O4[12])); 
	AO_CELL inst_5_12 ( 
	.A1(out_sel[10]), 
	.A2(I10[12]), 
	.B1(out_sel[11]), 
	.B2(I11[12]), 
	.Z(O5[12])); 
	AO_CELL inst_6_12 ( 
	.A1(out_sel[12]), 
	.A2(I12[12]), 
	.B1(out_sel[13]), 
	.B2(I13[12]), 
	.Z(O6[12])); 
	AO_CELL inst_7_12 ( 
	.A1(out_sel[14]), 
	.A2(I14[12]), 
	.B1(out_sel[15]), 
	.B2(I15[12]), 
	.Z(O7[12])); 
	AO_CELL inst_8_12 ( 
	.A1(out_sel[16]), 
	.A2(I16[12]), 
	.B1(out_sel[17]), 
	.B2(I17[12]), 
	.Z(O8[12])); 
	AO_CELL inst_9_12 ( 
	.A1(out_sel[18]), 
	.A2(I18[12]), 
	.B1(out_sel[19]), 
	.B2(I19[12]), 
	.Z(O9[12])); 
	AO_CELL inst_10_12 ( 
	.A1(out_sel[20]), 
	.A2(I20[12]), 
	.B1(out_sel[21]), 
	.B2(I21[12]), 
	.Z(O10[12])); 
	AO_CELL inst_11_12 ( 
	.A1(out_sel[22]), 
	.A2(I22[12]), 
	.B1(out_sel[23]), 
	.B2(I23[12]), 
	.Z(O11[12])); 
	AO_CELL inst_12_12 ( 
	.A1(out_sel[24]), 
	.A2(I24[12]), 
	.B1(out_sel[25]), 
	.B2(I25[12]), 
	.Z(O12[12])); 
	AO_CELL inst_13_12 ( 
	.A1(out_sel[26]), 
	.A2(I26[12]), 
	.B1(out_sel[27]), 
	.B2(I27[12]), 
	.Z(O13[12])); 
	AO_CELL inst_14_12 ( 
	.A1(out_sel[28]), 
	.A2(I28[12]), 
	.B1(out_sel[29]), 
	.B2(I29[12]), 
	.Z(O14[12])); 
	AO_CELL inst_15_12 ( 
	.A1(out_sel[30]), 
	.A2(I30[12]), 
	.B1(out_sel[31]), 
	.B2(I31[12]), 
	.Z(O15[12])); 
	AO_CELL inst_16_12 ( 
	.A1(out_sel[32]), 
	.A2(I32[12]), 
	.B1(out_sel[33]), 
	.B2(I33[12]), 
	.Z(O16[12])); 
	AO_CELL inst_17_12 ( 
	.A1(out_sel[34]), 
	.A2(I34[12]), 
	.B1(out_sel[35]), 
	.B2(I35[12]), 
	.Z(O17[12])); 
	AO_CELL inst_18_12 ( 
	.A1(out_sel[36]), 
	.A2(I36[12]), 
	.B1(out_sel[37]), 
	.B2(I37[12]), 
	.Z(O18[12])); 
	AO_CELL inst_19_12 ( 
	.A1(out_sel[38]), 
	.A2(I38[12]), 
	.B1(out_sel[39]), 
	.B2(I39[12]), 
	.Z(O19[12])); 
	AO_CELL inst_20_12 ( 
	.A1(out_sel[40]), 
	.A2(I40[12]), 
	.B1(out_sel[41]), 
	.B2(I41[12]), 
	.Z(O20[12])); 
	AO_CELL inst_21_12 ( 
	.A1(out_sel[42]), 
	.A2(I42[12]), 
	.B1(out_sel[43]), 
	.B2(I43[12]), 
	.Z(O21[12])); 
	AO_CELL inst_22_12 ( 
	.A1(out_sel[44]), 
	.A2(I44[12]), 
	.B1(out_sel[45]), 
	.B2(I45[12]), 
	.Z(O22[12])); 
	AN_CELL inst_and_12 ( 
	.A1(out_sel[46]), 
	.A2(I46[12]), 
	.Z(O23[12])); 
	AO_CELL inst_0_13 ( 
	.A1(out_sel[0]), 
	.A2(I0[13]), 
	.B1(out_sel[1]), 
	.B2(I1[13]), 
	.Z(O0[13])); 
	AO_CELL inst_1_13 ( 
	.A1(out_sel[2]), 
	.A2(I2[13]), 
	.B1(out_sel[3]), 
	.B2(I3[13]), 
	.Z(O1[13])); 
	AO_CELL inst_2_13 ( 
	.A1(out_sel[4]), 
	.A2(I4[13]), 
	.B1(out_sel[5]), 
	.B2(I5[13]), 
	.Z(O2[13])); 
	AO_CELL inst_3_13 ( 
	.A1(out_sel[6]), 
	.A2(I6[13]), 
	.B1(out_sel[7]), 
	.B2(I7[13]), 
	.Z(O3[13])); 
	AO_CELL inst_4_13 ( 
	.A1(out_sel[8]), 
	.A2(I8[13]), 
	.B1(out_sel[9]), 
	.B2(I9[13]), 
	.Z(O4[13])); 
	AO_CELL inst_5_13 ( 
	.A1(out_sel[10]), 
	.A2(I10[13]), 
	.B1(out_sel[11]), 
	.B2(I11[13]), 
	.Z(O5[13])); 
	AO_CELL inst_6_13 ( 
	.A1(out_sel[12]), 
	.A2(I12[13]), 
	.B1(out_sel[13]), 
	.B2(I13[13]), 
	.Z(O6[13])); 
	AO_CELL inst_7_13 ( 
	.A1(out_sel[14]), 
	.A2(I14[13]), 
	.B1(out_sel[15]), 
	.B2(I15[13]), 
	.Z(O7[13])); 
	AO_CELL inst_8_13 ( 
	.A1(out_sel[16]), 
	.A2(I16[13]), 
	.B1(out_sel[17]), 
	.B2(I17[13]), 
	.Z(O8[13])); 
	AO_CELL inst_9_13 ( 
	.A1(out_sel[18]), 
	.A2(I18[13]), 
	.B1(out_sel[19]), 
	.B2(I19[13]), 
	.Z(O9[13])); 
	AO_CELL inst_10_13 ( 
	.A1(out_sel[20]), 
	.A2(I20[13]), 
	.B1(out_sel[21]), 
	.B2(I21[13]), 
	.Z(O10[13])); 
	AO_CELL inst_11_13 ( 
	.A1(out_sel[22]), 
	.A2(I22[13]), 
	.B1(out_sel[23]), 
	.B2(I23[13]), 
	.Z(O11[13])); 
	AO_CELL inst_12_13 ( 
	.A1(out_sel[24]), 
	.A2(I24[13]), 
	.B1(out_sel[25]), 
	.B2(I25[13]), 
	.Z(O12[13])); 
	AO_CELL inst_13_13 ( 
	.A1(out_sel[26]), 
	.A2(I26[13]), 
	.B1(out_sel[27]), 
	.B2(I27[13]), 
	.Z(O13[13])); 
	AO_CELL inst_14_13 ( 
	.A1(out_sel[28]), 
	.A2(I28[13]), 
	.B1(out_sel[29]), 
	.B2(I29[13]), 
	.Z(O14[13])); 
	AO_CELL inst_15_13 ( 
	.A1(out_sel[30]), 
	.A2(I30[13]), 
	.B1(out_sel[31]), 
	.B2(I31[13]), 
	.Z(O15[13])); 
	AO_CELL inst_16_13 ( 
	.A1(out_sel[32]), 
	.A2(I32[13]), 
	.B1(out_sel[33]), 
	.B2(I33[13]), 
	.Z(O16[13])); 
	AO_CELL inst_17_13 ( 
	.A1(out_sel[34]), 
	.A2(I34[13]), 
	.B1(out_sel[35]), 
	.B2(I35[13]), 
	.Z(O17[13])); 
	AO_CELL inst_18_13 ( 
	.A1(out_sel[36]), 
	.A2(I36[13]), 
	.B1(out_sel[37]), 
	.B2(I37[13]), 
	.Z(O18[13])); 
	AO_CELL inst_19_13 ( 
	.A1(out_sel[38]), 
	.A2(I38[13]), 
	.B1(out_sel[39]), 
	.B2(I39[13]), 
	.Z(O19[13])); 
	AO_CELL inst_20_13 ( 
	.A1(out_sel[40]), 
	.A2(I40[13]), 
	.B1(out_sel[41]), 
	.B2(I41[13]), 
	.Z(O20[13])); 
	AO_CELL inst_21_13 ( 
	.A1(out_sel[42]), 
	.A2(I42[13]), 
	.B1(out_sel[43]), 
	.B2(I43[13]), 
	.Z(O21[13])); 
	AO_CELL inst_22_13 ( 
	.A1(out_sel[44]), 
	.A2(I44[13]), 
	.B1(out_sel[45]), 
	.B2(I45[13]), 
	.Z(O22[13])); 
	AN_CELL inst_and_13 ( 
	.A1(out_sel[46]), 
	.A2(I46[13]), 
	.Z(O23[13])); 
	AO_CELL inst_0_14 ( 
	.A1(out_sel[0]), 
	.A2(I0[14]), 
	.B1(out_sel[1]), 
	.B2(I1[14]), 
	.Z(O0[14])); 
	AO_CELL inst_1_14 ( 
	.A1(out_sel[2]), 
	.A2(I2[14]), 
	.B1(out_sel[3]), 
	.B2(I3[14]), 
	.Z(O1[14])); 
	AO_CELL inst_2_14 ( 
	.A1(out_sel[4]), 
	.A2(I4[14]), 
	.B1(out_sel[5]), 
	.B2(I5[14]), 
	.Z(O2[14])); 
	AO_CELL inst_3_14 ( 
	.A1(out_sel[6]), 
	.A2(I6[14]), 
	.B1(out_sel[7]), 
	.B2(I7[14]), 
	.Z(O3[14])); 
	AO_CELL inst_4_14 ( 
	.A1(out_sel[8]), 
	.A2(I8[14]), 
	.B1(out_sel[9]), 
	.B2(I9[14]), 
	.Z(O4[14])); 
	AO_CELL inst_5_14 ( 
	.A1(out_sel[10]), 
	.A2(I10[14]), 
	.B1(out_sel[11]), 
	.B2(I11[14]), 
	.Z(O5[14])); 
	AO_CELL inst_6_14 ( 
	.A1(out_sel[12]), 
	.A2(I12[14]), 
	.B1(out_sel[13]), 
	.B2(I13[14]), 
	.Z(O6[14])); 
	AO_CELL inst_7_14 ( 
	.A1(out_sel[14]), 
	.A2(I14[14]), 
	.B1(out_sel[15]), 
	.B2(I15[14]), 
	.Z(O7[14])); 
	AO_CELL inst_8_14 ( 
	.A1(out_sel[16]), 
	.A2(I16[14]), 
	.B1(out_sel[17]), 
	.B2(I17[14]), 
	.Z(O8[14])); 
	AO_CELL inst_9_14 ( 
	.A1(out_sel[18]), 
	.A2(I18[14]), 
	.B1(out_sel[19]), 
	.B2(I19[14]), 
	.Z(O9[14])); 
	AO_CELL inst_10_14 ( 
	.A1(out_sel[20]), 
	.A2(I20[14]), 
	.B1(out_sel[21]), 
	.B2(I21[14]), 
	.Z(O10[14])); 
	AO_CELL inst_11_14 ( 
	.A1(out_sel[22]), 
	.A2(I22[14]), 
	.B1(out_sel[23]), 
	.B2(I23[14]), 
	.Z(O11[14])); 
	AO_CELL inst_12_14 ( 
	.A1(out_sel[24]), 
	.A2(I24[14]), 
	.B1(out_sel[25]), 
	.B2(I25[14]), 
	.Z(O12[14])); 
	AO_CELL inst_13_14 ( 
	.A1(out_sel[26]), 
	.A2(I26[14]), 
	.B1(out_sel[27]), 
	.B2(I27[14]), 
	.Z(O13[14])); 
	AO_CELL inst_14_14 ( 
	.A1(out_sel[28]), 
	.A2(I28[14]), 
	.B1(out_sel[29]), 
	.B2(I29[14]), 
	.Z(O14[14])); 
	AO_CELL inst_15_14 ( 
	.A1(out_sel[30]), 
	.A2(I30[14]), 
	.B1(out_sel[31]), 
	.B2(I31[14]), 
	.Z(O15[14])); 
	AO_CELL inst_16_14 ( 
	.A1(out_sel[32]), 
	.A2(I32[14]), 
	.B1(out_sel[33]), 
	.B2(I33[14]), 
	.Z(O16[14])); 
	AO_CELL inst_17_14 ( 
	.A1(out_sel[34]), 
	.A2(I34[14]), 
	.B1(out_sel[35]), 
	.B2(I35[14]), 
	.Z(O17[14])); 
	AO_CELL inst_18_14 ( 
	.A1(out_sel[36]), 
	.A2(I36[14]), 
	.B1(out_sel[37]), 
	.B2(I37[14]), 
	.Z(O18[14])); 
	AO_CELL inst_19_14 ( 
	.A1(out_sel[38]), 
	.A2(I38[14]), 
	.B1(out_sel[39]), 
	.B2(I39[14]), 
	.Z(O19[14])); 
	AO_CELL inst_20_14 ( 
	.A1(out_sel[40]), 
	.A2(I40[14]), 
	.B1(out_sel[41]), 
	.B2(I41[14]), 
	.Z(O20[14])); 
	AO_CELL inst_21_14 ( 
	.A1(out_sel[42]), 
	.A2(I42[14]), 
	.B1(out_sel[43]), 
	.B2(I43[14]), 
	.Z(O21[14])); 
	AO_CELL inst_22_14 ( 
	.A1(out_sel[44]), 
	.A2(I44[14]), 
	.B1(out_sel[45]), 
	.B2(I45[14]), 
	.Z(O22[14])); 
	AN_CELL inst_and_14 ( 
	.A1(out_sel[46]), 
	.A2(I46[14]), 
	.Z(O23[14])); 
	AO_CELL inst_0_15 ( 
	.A1(out_sel[0]), 
	.A2(I0[15]), 
	.B1(out_sel[1]), 
	.B2(I1[15]), 
	.Z(O0[15])); 
	AO_CELL inst_1_15 ( 
	.A1(out_sel[2]), 
	.A2(I2[15]), 
	.B1(out_sel[3]), 
	.B2(I3[15]), 
	.Z(O1[15])); 
	AO_CELL inst_2_15 ( 
	.A1(out_sel[4]), 
	.A2(I4[15]), 
	.B1(out_sel[5]), 
	.B2(I5[15]), 
	.Z(O2[15])); 
	AO_CELL inst_3_15 ( 
	.A1(out_sel[6]), 
	.A2(I6[15]), 
	.B1(out_sel[7]), 
	.B2(I7[15]), 
	.Z(O3[15])); 
	AO_CELL inst_4_15 ( 
	.A1(out_sel[8]), 
	.A2(I8[15]), 
	.B1(out_sel[9]), 
	.B2(I9[15]), 
	.Z(O4[15])); 
	AO_CELL inst_5_15 ( 
	.A1(out_sel[10]), 
	.A2(I10[15]), 
	.B1(out_sel[11]), 
	.B2(I11[15]), 
	.Z(O5[15])); 
	AO_CELL inst_6_15 ( 
	.A1(out_sel[12]), 
	.A2(I12[15]), 
	.B1(out_sel[13]), 
	.B2(I13[15]), 
	.Z(O6[15])); 
	AO_CELL inst_7_15 ( 
	.A1(out_sel[14]), 
	.A2(I14[15]), 
	.B1(out_sel[15]), 
	.B2(I15[15]), 
	.Z(O7[15])); 
	AO_CELL inst_8_15 ( 
	.A1(out_sel[16]), 
	.A2(I16[15]), 
	.B1(out_sel[17]), 
	.B2(I17[15]), 
	.Z(O8[15])); 
	AO_CELL inst_9_15 ( 
	.A1(out_sel[18]), 
	.A2(I18[15]), 
	.B1(out_sel[19]), 
	.B2(I19[15]), 
	.Z(O9[15])); 
	AO_CELL inst_10_15 ( 
	.A1(out_sel[20]), 
	.A2(I20[15]), 
	.B1(out_sel[21]), 
	.B2(I21[15]), 
	.Z(O10[15])); 
	AO_CELL inst_11_15 ( 
	.A1(out_sel[22]), 
	.A2(I22[15]), 
	.B1(out_sel[23]), 
	.B2(I23[15]), 
	.Z(O11[15])); 
	AO_CELL inst_12_15 ( 
	.A1(out_sel[24]), 
	.A2(I24[15]), 
	.B1(out_sel[25]), 
	.B2(I25[15]), 
	.Z(O12[15])); 
	AO_CELL inst_13_15 ( 
	.A1(out_sel[26]), 
	.A2(I26[15]), 
	.B1(out_sel[27]), 
	.B2(I27[15]), 
	.Z(O13[15])); 
	AO_CELL inst_14_15 ( 
	.A1(out_sel[28]), 
	.A2(I28[15]), 
	.B1(out_sel[29]), 
	.B2(I29[15]), 
	.Z(O14[15])); 
	AO_CELL inst_15_15 ( 
	.A1(out_sel[30]), 
	.A2(I30[15]), 
	.B1(out_sel[31]), 
	.B2(I31[15]), 
	.Z(O15[15])); 
	AO_CELL inst_16_15 ( 
	.A1(out_sel[32]), 
	.A2(I32[15]), 
	.B1(out_sel[33]), 
	.B2(I33[15]), 
	.Z(O16[15])); 
	AO_CELL inst_17_15 ( 
	.A1(out_sel[34]), 
	.A2(I34[15]), 
	.B1(out_sel[35]), 
	.B2(I35[15]), 
	.Z(O17[15])); 
	AO_CELL inst_18_15 ( 
	.A1(out_sel[36]), 
	.A2(I36[15]), 
	.B1(out_sel[37]), 
	.B2(I37[15]), 
	.Z(O18[15])); 
	AO_CELL inst_19_15 ( 
	.A1(out_sel[38]), 
	.A2(I38[15]), 
	.B1(out_sel[39]), 
	.B2(I39[15]), 
	.Z(O19[15])); 
	AO_CELL inst_20_15 ( 
	.A1(out_sel[40]), 
	.A2(I40[15]), 
	.B1(out_sel[41]), 
	.B2(I41[15]), 
	.Z(O20[15])); 
	AO_CELL inst_21_15 ( 
	.A1(out_sel[42]), 
	.A2(I42[15]), 
	.B1(out_sel[43]), 
	.B2(I43[15]), 
	.Z(O21[15])); 
	AO_CELL inst_22_15 ( 
	.A1(out_sel[44]), 
	.A2(I44[15]), 
	.B1(out_sel[45]), 
	.B2(I45[15]), 
	.Z(O22[15])); 
	AN_CELL inst_and_15 ( 
	.A1(out_sel[46]), 
	.A2(I46[15]), 
	.Z(O23[15])); 
	AO_CELL inst_0_16 ( 
	.A1(out_sel[0]), 
	.A2(I0[16]), 
	.B1(out_sel[1]), 
	.B2(I1[16]), 
	.Z(O0[16])); 
	AO_CELL inst_1_16 ( 
	.A1(out_sel[2]), 
	.A2(I2[16]), 
	.B1(out_sel[3]), 
	.B2(I3[16]), 
	.Z(O1[16])); 
	AO_CELL inst_2_16 ( 
	.A1(out_sel[4]), 
	.A2(I4[16]), 
	.B1(out_sel[5]), 
	.B2(I5[16]), 
	.Z(O2[16])); 
	AO_CELL inst_3_16 ( 
	.A1(out_sel[6]), 
	.A2(I6[16]), 
	.B1(out_sel[7]), 
	.B2(I7[16]), 
	.Z(O3[16])); 
	AO_CELL inst_4_16 ( 
	.A1(out_sel[8]), 
	.A2(I8[16]), 
	.B1(out_sel[9]), 
	.B2(I9[16]), 
	.Z(O4[16])); 
	AO_CELL inst_5_16 ( 
	.A1(out_sel[10]), 
	.A2(I10[16]), 
	.B1(out_sel[11]), 
	.B2(I11[16]), 
	.Z(O5[16])); 
	AO_CELL inst_6_16 ( 
	.A1(out_sel[12]), 
	.A2(I12[16]), 
	.B1(out_sel[13]), 
	.B2(I13[16]), 
	.Z(O6[16])); 
	AO_CELL inst_7_16 ( 
	.A1(out_sel[14]), 
	.A2(I14[16]), 
	.B1(out_sel[15]), 
	.B2(I15[16]), 
	.Z(O7[16])); 
	AO_CELL inst_8_16 ( 
	.A1(out_sel[16]), 
	.A2(I16[16]), 
	.B1(out_sel[17]), 
	.B2(I17[16]), 
	.Z(O8[16])); 
	AO_CELL inst_9_16 ( 
	.A1(out_sel[18]), 
	.A2(I18[16]), 
	.B1(out_sel[19]), 
	.B2(I19[16]), 
	.Z(O9[16])); 
	AO_CELL inst_10_16 ( 
	.A1(out_sel[20]), 
	.A2(I20[16]), 
	.B1(out_sel[21]), 
	.B2(I21[16]), 
	.Z(O10[16])); 
	AO_CELL inst_11_16 ( 
	.A1(out_sel[22]), 
	.A2(I22[16]), 
	.B1(out_sel[23]), 
	.B2(I23[16]), 
	.Z(O11[16])); 
	AO_CELL inst_12_16 ( 
	.A1(out_sel[24]), 
	.A2(I24[16]), 
	.B1(out_sel[25]), 
	.B2(I25[16]), 
	.Z(O12[16])); 
	AO_CELL inst_13_16 ( 
	.A1(out_sel[26]), 
	.A2(I26[16]), 
	.B1(out_sel[27]), 
	.B2(I27[16]), 
	.Z(O13[16])); 
	AO_CELL inst_14_16 ( 
	.A1(out_sel[28]), 
	.A2(I28[16]), 
	.B1(out_sel[29]), 
	.B2(I29[16]), 
	.Z(O14[16])); 
	AO_CELL inst_15_16 ( 
	.A1(out_sel[30]), 
	.A2(I30[16]), 
	.B1(out_sel[31]), 
	.B2(I31[16]), 
	.Z(O15[16])); 
	AO_CELL inst_16_16 ( 
	.A1(out_sel[32]), 
	.A2(I32[16]), 
	.B1(out_sel[33]), 
	.B2(I33[16]), 
	.Z(O16[16])); 
	AO_CELL inst_17_16 ( 
	.A1(out_sel[34]), 
	.A2(I34[16]), 
	.B1(out_sel[35]), 
	.B2(I35[16]), 
	.Z(O17[16])); 
	AO_CELL inst_18_16 ( 
	.A1(out_sel[36]), 
	.A2(I36[16]), 
	.B1(out_sel[37]), 
	.B2(I37[16]), 
	.Z(O18[16])); 
	AO_CELL inst_19_16 ( 
	.A1(out_sel[38]), 
	.A2(I38[16]), 
	.B1(out_sel[39]), 
	.B2(I39[16]), 
	.Z(O19[16])); 
	AO_CELL inst_20_16 ( 
	.A1(out_sel[40]), 
	.A2(I40[16]), 
	.B1(out_sel[41]), 
	.B2(I41[16]), 
	.Z(O20[16])); 
	AO_CELL inst_21_16 ( 
	.A1(out_sel[42]), 
	.A2(I42[16]), 
	.B1(out_sel[43]), 
	.B2(I43[16]), 
	.Z(O21[16])); 
	AO_CELL inst_22_16 ( 
	.A1(out_sel[44]), 
	.A2(I44[16]), 
	.B1(out_sel[45]), 
	.B2(I45[16]), 
	.Z(O22[16])); 
	AN_CELL inst_and_16 ( 
	.A1(out_sel[46]), 
	.A2(I46[16]), 
	.Z(O23[16])); 
	AO_CELL inst_0_17 ( 
	.A1(out_sel[0]), 
	.A2(I0[17]), 
	.B1(out_sel[1]), 
	.B2(I1[17]), 
	.Z(O0[17])); 
	AO_CELL inst_1_17 ( 
	.A1(out_sel[2]), 
	.A2(I2[17]), 
	.B1(out_sel[3]), 
	.B2(I3[17]), 
	.Z(O1[17])); 
	AO_CELL inst_2_17 ( 
	.A1(out_sel[4]), 
	.A2(I4[17]), 
	.B1(out_sel[5]), 
	.B2(I5[17]), 
	.Z(O2[17])); 
	AO_CELL inst_3_17 ( 
	.A1(out_sel[6]), 
	.A2(I6[17]), 
	.B1(out_sel[7]), 
	.B2(I7[17]), 
	.Z(O3[17])); 
	AO_CELL inst_4_17 ( 
	.A1(out_sel[8]), 
	.A2(I8[17]), 
	.B1(out_sel[9]), 
	.B2(I9[17]), 
	.Z(O4[17])); 
	AO_CELL inst_5_17 ( 
	.A1(out_sel[10]), 
	.A2(I10[17]), 
	.B1(out_sel[11]), 
	.B2(I11[17]), 
	.Z(O5[17])); 
	AO_CELL inst_6_17 ( 
	.A1(out_sel[12]), 
	.A2(I12[17]), 
	.B1(out_sel[13]), 
	.B2(I13[17]), 
	.Z(O6[17])); 
	AO_CELL inst_7_17 ( 
	.A1(out_sel[14]), 
	.A2(I14[17]), 
	.B1(out_sel[15]), 
	.B2(I15[17]), 
	.Z(O7[17])); 
	AO_CELL inst_8_17 ( 
	.A1(out_sel[16]), 
	.A2(I16[17]), 
	.B1(out_sel[17]), 
	.B2(I17[17]), 
	.Z(O8[17])); 
	AO_CELL inst_9_17 ( 
	.A1(out_sel[18]), 
	.A2(I18[17]), 
	.B1(out_sel[19]), 
	.B2(I19[17]), 
	.Z(O9[17])); 
	AO_CELL inst_10_17 ( 
	.A1(out_sel[20]), 
	.A2(I20[17]), 
	.B1(out_sel[21]), 
	.B2(I21[17]), 
	.Z(O10[17])); 
	AO_CELL inst_11_17 ( 
	.A1(out_sel[22]), 
	.A2(I22[17]), 
	.B1(out_sel[23]), 
	.B2(I23[17]), 
	.Z(O11[17])); 
	AO_CELL inst_12_17 ( 
	.A1(out_sel[24]), 
	.A2(I24[17]), 
	.B1(out_sel[25]), 
	.B2(I25[17]), 
	.Z(O12[17])); 
	AO_CELL inst_13_17 ( 
	.A1(out_sel[26]), 
	.A2(I26[17]), 
	.B1(out_sel[27]), 
	.B2(I27[17]), 
	.Z(O13[17])); 
	AO_CELL inst_14_17 ( 
	.A1(out_sel[28]), 
	.A2(I28[17]), 
	.B1(out_sel[29]), 
	.B2(I29[17]), 
	.Z(O14[17])); 
	AO_CELL inst_15_17 ( 
	.A1(out_sel[30]), 
	.A2(I30[17]), 
	.B1(out_sel[31]), 
	.B2(I31[17]), 
	.Z(O15[17])); 
	AO_CELL inst_16_17 ( 
	.A1(out_sel[32]), 
	.A2(I32[17]), 
	.B1(out_sel[33]), 
	.B2(I33[17]), 
	.Z(O16[17])); 
	AO_CELL inst_17_17 ( 
	.A1(out_sel[34]), 
	.A2(I34[17]), 
	.B1(out_sel[35]), 
	.B2(I35[17]), 
	.Z(O17[17])); 
	AO_CELL inst_18_17 ( 
	.A1(out_sel[36]), 
	.A2(I36[17]), 
	.B1(out_sel[37]), 
	.B2(I37[17]), 
	.Z(O18[17])); 
	AO_CELL inst_19_17 ( 
	.A1(out_sel[38]), 
	.A2(I38[17]), 
	.B1(out_sel[39]), 
	.B2(I39[17]), 
	.Z(O19[17])); 
	AO_CELL inst_20_17 ( 
	.A1(out_sel[40]), 
	.A2(I40[17]), 
	.B1(out_sel[41]), 
	.B2(I41[17]), 
	.Z(O20[17])); 
	AO_CELL inst_21_17 ( 
	.A1(out_sel[42]), 
	.A2(I42[17]), 
	.B1(out_sel[43]), 
	.B2(I43[17]), 
	.Z(O21[17])); 
	AO_CELL inst_22_17 ( 
	.A1(out_sel[44]), 
	.A2(I44[17]), 
	.B1(out_sel[45]), 
	.B2(I45[17]), 
	.Z(O22[17])); 
	AN_CELL inst_and_17 ( 
	.A1(out_sel[46]), 
	.A2(I46[17]), 
	.Z(O23[17])); 
	AO_CELL inst_0_18 ( 
	.A1(out_sel[0]), 
	.A2(I0[18]), 
	.B1(out_sel[1]), 
	.B2(I1[18]), 
	.Z(O0[18])); 
	AO_CELL inst_1_18 ( 
	.A1(out_sel[2]), 
	.A2(I2[18]), 
	.B1(out_sel[3]), 
	.B2(I3[18]), 
	.Z(O1[18])); 
	AO_CELL inst_2_18 ( 
	.A1(out_sel[4]), 
	.A2(I4[18]), 
	.B1(out_sel[5]), 
	.B2(I5[18]), 
	.Z(O2[18])); 
	AO_CELL inst_3_18 ( 
	.A1(out_sel[6]), 
	.A2(I6[18]), 
	.B1(out_sel[7]), 
	.B2(I7[18]), 
	.Z(O3[18])); 
	AO_CELL inst_4_18 ( 
	.A1(out_sel[8]), 
	.A2(I8[18]), 
	.B1(out_sel[9]), 
	.B2(I9[18]), 
	.Z(O4[18])); 
	AO_CELL inst_5_18 ( 
	.A1(out_sel[10]), 
	.A2(I10[18]), 
	.B1(out_sel[11]), 
	.B2(I11[18]), 
	.Z(O5[18])); 
	AO_CELL inst_6_18 ( 
	.A1(out_sel[12]), 
	.A2(I12[18]), 
	.B1(out_sel[13]), 
	.B2(I13[18]), 
	.Z(O6[18])); 
	AO_CELL inst_7_18 ( 
	.A1(out_sel[14]), 
	.A2(I14[18]), 
	.B1(out_sel[15]), 
	.B2(I15[18]), 
	.Z(O7[18])); 
	AO_CELL inst_8_18 ( 
	.A1(out_sel[16]), 
	.A2(I16[18]), 
	.B1(out_sel[17]), 
	.B2(I17[18]), 
	.Z(O8[18])); 
	AO_CELL inst_9_18 ( 
	.A1(out_sel[18]), 
	.A2(I18[18]), 
	.B1(out_sel[19]), 
	.B2(I19[18]), 
	.Z(O9[18])); 
	AO_CELL inst_10_18 ( 
	.A1(out_sel[20]), 
	.A2(I20[18]), 
	.B1(out_sel[21]), 
	.B2(I21[18]), 
	.Z(O10[18])); 
	AO_CELL inst_11_18 ( 
	.A1(out_sel[22]), 
	.A2(I22[18]), 
	.B1(out_sel[23]), 
	.B2(I23[18]), 
	.Z(O11[18])); 
	AO_CELL inst_12_18 ( 
	.A1(out_sel[24]), 
	.A2(I24[18]), 
	.B1(out_sel[25]), 
	.B2(I25[18]), 
	.Z(O12[18])); 
	AO_CELL inst_13_18 ( 
	.A1(out_sel[26]), 
	.A2(I26[18]), 
	.B1(out_sel[27]), 
	.B2(I27[18]), 
	.Z(O13[18])); 
	AO_CELL inst_14_18 ( 
	.A1(out_sel[28]), 
	.A2(I28[18]), 
	.B1(out_sel[29]), 
	.B2(I29[18]), 
	.Z(O14[18])); 
	AO_CELL inst_15_18 ( 
	.A1(out_sel[30]), 
	.A2(I30[18]), 
	.B1(out_sel[31]), 
	.B2(I31[18]), 
	.Z(O15[18])); 
	AO_CELL inst_16_18 ( 
	.A1(out_sel[32]), 
	.A2(I32[18]), 
	.B1(out_sel[33]), 
	.B2(I33[18]), 
	.Z(O16[18])); 
	AO_CELL inst_17_18 ( 
	.A1(out_sel[34]), 
	.A2(I34[18]), 
	.B1(out_sel[35]), 
	.B2(I35[18]), 
	.Z(O17[18])); 
	AO_CELL inst_18_18 ( 
	.A1(out_sel[36]), 
	.A2(I36[18]), 
	.B1(out_sel[37]), 
	.B2(I37[18]), 
	.Z(O18[18])); 
	AO_CELL inst_19_18 ( 
	.A1(out_sel[38]), 
	.A2(I38[18]), 
	.B1(out_sel[39]), 
	.B2(I39[18]), 
	.Z(O19[18])); 
	AO_CELL inst_20_18 ( 
	.A1(out_sel[40]), 
	.A2(I40[18]), 
	.B1(out_sel[41]), 
	.B2(I41[18]), 
	.Z(O20[18])); 
	AO_CELL inst_21_18 ( 
	.A1(out_sel[42]), 
	.A2(I42[18]), 
	.B1(out_sel[43]), 
	.B2(I43[18]), 
	.Z(O21[18])); 
	AO_CELL inst_22_18 ( 
	.A1(out_sel[44]), 
	.A2(I44[18]), 
	.B1(out_sel[45]), 
	.B2(I45[18]), 
	.Z(O22[18])); 
	AN_CELL inst_and_18 ( 
	.A1(out_sel[46]), 
	.A2(I46[18]), 
	.Z(O23[18])); 
	AO_CELL inst_0_19 ( 
	.A1(out_sel[0]), 
	.A2(I0[19]), 
	.B1(out_sel[1]), 
	.B2(I1[19]), 
	.Z(O0[19])); 
	AO_CELL inst_1_19 ( 
	.A1(out_sel[2]), 
	.A2(I2[19]), 
	.B1(out_sel[3]), 
	.B2(I3[19]), 
	.Z(O1[19])); 
	AO_CELL inst_2_19 ( 
	.A1(out_sel[4]), 
	.A2(I4[19]), 
	.B1(out_sel[5]), 
	.B2(I5[19]), 
	.Z(O2[19])); 
	AO_CELL inst_3_19 ( 
	.A1(out_sel[6]), 
	.A2(I6[19]), 
	.B1(out_sel[7]), 
	.B2(I7[19]), 
	.Z(O3[19])); 
	AO_CELL inst_4_19 ( 
	.A1(out_sel[8]), 
	.A2(I8[19]), 
	.B1(out_sel[9]), 
	.B2(I9[19]), 
	.Z(O4[19])); 
	AO_CELL inst_5_19 ( 
	.A1(out_sel[10]), 
	.A2(I10[19]), 
	.B1(out_sel[11]), 
	.B2(I11[19]), 
	.Z(O5[19])); 
	AO_CELL inst_6_19 ( 
	.A1(out_sel[12]), 
	.A2(I12[19]), 
	.B1(out_sel[13]), 
	.B2(I13[19]), 
	.Z(O6[19])); 
	AO_CELL inst_7_19 ( 
	.A1(out_sel[14]), 
	.A2(I14[19]), 
	.B1(out_sel[15]), 
	.B2(I15[19]), 
	.Z(O7[19])); 
	AO_CELL inst_8_19 ( 
	.A1(out_sel[16]), 
	.A2(I16[19]), 
	.B1(out_sel[17]), 
	.B2(I17[19]), 
	.Z(O8[19])); 
	AO_CELL inst_9_19 ( 
	.A1(out_sel[18]), 
	.A2(I18[19]), 
	.B1(out_sel[19]), 
	.B2(I19[19]), 
	.Z(O9[19])); 
	AO_CELL inst_10_19 ( 
	.A1(out_sel[20]), 
	.A2(I20[19]), 
	.B1(out_sel[21]), 
	.B2(I21[19]), 
	.Z(O10[19])); 
	AO_CELL inst_11_19 ( 
	.A1(out_sel[22]), 
	.A2(I22[19]), 
	.B1(out_sel[23]), 
	.B2(I23[19]), 
	.Z(O11[19])); 
	AO_CELL inst_12_19 ( 
	.A1(out_sel[24]), 
	.A2(I24[19]), 
	.B1(out_sel[25]), 
	.B2(I25[19]), 
	.Z(O12[19])); 
	AO_CELL inst_13_19 ( 
	.A1(out_sel[26]), 
	.A2(I26[19]), 
	.B1(out_sel[27]), 
	.B2(I27[19]), 
	.Z(O13[19])); 
	AO_CELL inst_14_19 ( 
	.A1(out_sel[28]), 
	.A2(I28[19]), 
	.B1(out_sel[29]), 
	.B2(I29[19]), 
	.Z(O14[19])); 
	AO_CELL inst_15_19 ( 
	.A1(out_sel[30]), 
	.A2(I30[19]), 
	.B1(out_sel[31]), 
	.B2(I31[19]), 
	.Z(O15[19])); 
	AO_CELL inst_16_19 ( 
	.A1(out_sel[32]), 
	.A2(I32[19]), 
	.B1(out_sel[33]), 
	.B2(I33[19]), 
	.Z(O16[19])); 
	AO_CELL inst_17_19 ( 
	.A1(out_sel[34]), 
	.A2(I34[19]), 
	.B1(out_sel[35]), 
	.B2(I35[19]), 
	.Z(O17[19])); 
	AO_CELL inst_18_19 ( 
	.A1(out_sel[36]), 
	.A2(I36[19]), 
	.B1(out_sel[37]), 
	.B2(I37[19]), 
	.Z(O18[19])); 
	AO_CELL inst_19_19 ( 
	.A1(out_sel[38]), 
	.A2(I38[19]), 
	.B1(out_sel[39]), 
	.B2(I39[19]), 
	.Z(O19[19])); 
	AO_CELL inst_20_19 ( 
	.A1(out_sel[40]), 
	.A2(I40[19]), 
	.B1(out_sel[41]), 
	.B2(I41[19]), 
	.Z(O20[19])); 
	AO_CELL inst_21_19 ( 
	.A1(out_sel[42]), 
	.A2(I42[19]), 
	.B1(out_sel[43]), 
	.B2(I43[19]), 
	.Z(O21[19])); 
	AO_CELL inst_22_19 ( 
	.A1(out_sel[44]), 
	.A2(I44[19]), 
	.B1(out_sel[45]), 
	.B2(I45[19]), 
	.Z(O22[19])); 
	AN_CELL inst_and_19 ( 
	.A1(out_sel[46]), 
	.A2(I46[19]), 
	.Z(O23[19])); 
	AO_CELL inst_0_20 ( 
	.A1(out_sel[0]), 
	.A2(I0[20]), 
	.B1(out_sel[1]), 
	.B2(I1[20]), 
	.Z(O0[20])); 
	AO_CELL inst_1_20 ( 
	.A1(out_sel[2]), 
	.A2(I2[20]), 
	.B1(out_sel[3]), 
	.B2(I3[20]), 
	.Z(O1[20])); 
	AO_CELL inst_2_20 ( 
	.A1(out_sel[4]), 
	.A2(I4[20]), 
	.B1(out_sel[5]), 
	.B2(I5[20]), 
	.Z(O2[20])); 
	AO_CELL inst_3_20 ( 
	.A1(out_sel[6]), 
	.A2(I6[20]), 
	.B1(out_sel[7]), 
	.B2(I7[20]), 
	.Z(O3[20])); 
	AO_CELL inst_4_20 ( 
	.A1(out_sel[8]), 
	.A2(I8[20]), 
	.B1(out_sel[9]), 
	.B2(I9[20]), 
	.Z(O4[20])); 
	AO_CELL inst_5_20 ( 
	.A1(out_sel[10]), 
	.A2(I10[20]), 
	.B1(out_sel[11]), 
	.B2(I11[20]), 
	.Z(O5[20])); 
	AO_CELL inst_6_20 ( 
	.A1(out_sel[12]), 
	.A2(I12[20]), 
	.B1(out_sel[13]), 
	.B2(I13[20]), 
	.Z(O6[20])); 
	AO_CELL inst_7_20 ( 
	.A1(out_sel[14]), 
	.A2(I14[20]), 
	.B1(out_sel[15]), 
	.B2(I15[20]), 
	.Z(O7[20])); 
	AO_CELL inst_8_20 ( 
	.A1(out_sel[16]), 
	.A2(I16[20]), 
	.B1(out_sel[17]), 
	.B2(I17[20]), 
	.Z(O8[20])); 
	AO_CELL inst_9_20 ( 
	.A1(out_sel[18]), 
	.A2(I18[20]), 
	.B1(out_sel[19]), 
	.B2(I19[20]), 
	.Z(O9[20])); 
	AO_CELL inst_10_20 ( 
	.A1(out_sel[20]), 
	.A2(I20[20]), 
	.B1(out_sel[21]), 
	.B2(I21[20]), 
	.Z(O10[20])); 
	AO_CELL inst_11_20 ( 
	.A1(out_sel[22]), 
	.A2(I22[20]), 
	.B1(out_sel[23]), 
	.B2(I23[20]), 
	.Z(O11[20])); 
	AO_CELL inst_12_20 ( 
	.A1(out_sel[24]), 
	.A2(I24[20]), 
	.B1(out_sel[25]), 
	.B2(I25[20]), 
	.Z(O12[20])); 
	AO_CELL inst_13_20 ( 
	.A1(out_sel[26]), 
	.A2(I26[20]), 
	.B1(out_sel[27]), 
	.B2(I27[20]), 
	.Z(O13[20])); 
	AO_CELL inst_14_20 ( 
	.A1(out_sel[28]), 
	.A2(I28[20]), 
	.B1(out_sel[29]), 
	.B2(I29[20]), 
	.Z(O14[20])); 
	AO_CELL inst_15_20 ( 
	.A1(out_sel[30]), 
	.A2(I30[20]), 
	.B1(out_sel[31]), 
	.B2(I31[20]), 
	.Z(O15[20])); 
	AO_CELL inst_16_20 ( 
	.A1(out_sel[32]), 
	.A2(I32[20]), 
	.B1(out_sel[33]), 
	.B2(I33[20]), 
	.Z(O16[20])); 
	AO_CELL inst_17_20 ( 
	.A1(out_sel[34]), 
	.A2(I34[20]), 
	.B1(out_sel[35]), 
	.B2(I35[20]), 
	.Z(O17[20])); 
	AO_CELL inst_18_20 ( 
	.A1(out_sel[36]), 
	.A2(I36[20]), 
	.B1(out_sel[37]), 
	.B2(I37[20]), 
	.Z(O18[20])); 
	AO_CELL inst_19_20 ( 
	.A1(out_sel[38]), 
	.A2(I38[20]), 
	.B1(out_sel[39]), 
	.B2(I39[20]), 
	.Z(O19[20])); 
	AO_CELL inst_20_20 ( 
	.A1(out_sel[40]), 
	.A2(I40[20]), 
	.B1(out_sel[41]), 
	.B2(I41[20]), 
	.Z(O20[20])); 
	AO_CELL inst_21_20 ( 
	.A1(out_sel[42]), 
	.A2(I42[20]), 
	.B1(out_sel[43]), 
	.B2(I43[20]), 
	.Z(O21[20])); 
	AO_CELL inst_22_20 ( 
	.A1(out_sel[44]), 
	.A2(I44[20]), 
	.B1(out_sel[45]), 
	.B2(I45[20]), 
	.Z(O22[20])); 
	AN_CELL inst_and_20 ( 
	.A1(out_sel[46]), 
	.A2(I46[20]), 
	.Z(O23[20])); 
	AO_CELL inst_0_21 ( 
	.A1(out_sel[0]), 
	.A2(I0[21]), 
	.B1(out_sel[1]), 
	.B2(I1[21]), 
	.Z(O0[21])); 
	AO_CELL inst_1_21 ( 
	.A1(out_sel[2]), 
	.A2(I2[21]), 
	.B1(out_sel[3]), 
	.B2(I3[21]), 
	.Z(O1[21])); 
	AO_CELL inst_2_21 ( 
	.A1(out_sel[4]), 
	.A2(I4[21]), 
	.B1(out_sel[5]), 
	.B2(I5[21]), 
	.Z(O2[21])); 
	AO_CELL inst_3_21 ( 
	.A1(out_sel[6]), 
	.A2(I6[21]), 
	.B1(out_sel[7]), 
	.B2(I7[21]), 
	.Z(O3[21])); 
	AO_CELL inst_4_21 ( 
	.A1(out_sel[8]), 
	.A2(I8[21]), 
	.B1(out_sel[9]), 
	.B2(I9[21]), 
	.Z(O4[21])); 
	AO_CELL inst_5_21 ( 
	.A1(out_sel[10]), 
	.A2(I10[21]), 
	.B1(out_sel[11]), 
	.B2(I11[21]), 
	.Z(O5[21])); 
	AO_CELL inst_6_21 ( 
	.A1(out_sel[12]), 
	.A2(I12[21]), 
	.B1(out_sel[13]), 
	.B2(I13[21]), 
	.Z(O6[21])); 
	AO_CELL inst_7_21 ( 
	.A1(out_sel[14]), 
	.A2(I14[21]), 
	.B1(out_sel[15]), 
	.B2(I15[21]), 
	.Z(O7[21])); 
	AO_CELL inst_8_21 ( 
	.A1(out_sel[16]), 
	.A2(I16[21]), 
	.B1(out_sel[17]), 
	.B2(I17[21]), 
	.Z(O8[21])); 
	AO_CELL inst_9_21 ( 
	.A1(out_sel[18]), 
	.A2(I18[21]), 
	.B1(out_sel[19]), 
	.B2(I19[21]), 
	.Z(O9[21])); 
	AO_CELL inst_10_21 ( 
	.A1(out_sel[20]), 
	.A2(I20[21]), 
	.B1(out_sel[21]), 
	.B2(I21[21]), 
	.Z(O10[21])); 
	AO_CELL inst_11_21 ( 
	.A1(out_sel[22]), 
	.A2(I22[21]), 
	.B1(out_sel[23]), 
	.B2(I23[21]), 
	.Z(O11[21])); 
	AO_CELL inst_12_21 ( 
	.A1(out_sel[24]), 
	.A2(I24[21]), 
	.B1(out_sel[25]), 
	.B2(I25[21]), 
	.Z(O12[21])); 
	AO_CELL inst_13_21 ( 
	.A1(out_sel[26]), 
	.A2(I26[21]), 
	.B1(out_sel[27]), 
	.B2(I27[21]), 
	.Z(O13[21])); 
	AO_CELL inst_14_21 ( 
	.A1(out_sel[28]), 
	.A2(I28[21]), 
	.B1(out_sel[29]), 
	.B2(I29[21]), 
	.Z(O14[21])); 
	AO_CELL inst_15_21 ( 
	.A1(out_sel[30]), 
	.A2(I30[21]), 
	.B1(out_sel[31]), 
	.B2(I31[21]), 
	.Z(O15[21])); 
	AO_CELL inst_16_21 ( 
	.A1(out_sel[32]), 
	.A2(I32[21]), 
	.B1(out_sel[33]), 
	.B2(I33[21]), 
	.Z(O16[21])); 
	AO_CELL inst_17_21 ( 
	.A1(out_sel[34]), 
	.A2(I34[21]), 
	.B1(out_sel[35]), 
	.B2(I35[21]), 
	.Z(O17[21])); 
	AO_CELL inst_18_21 ( 
	.A1(out_sel[36]), 
	.A2(I36[21]), 
	.B1(out_sel[37]), 
	.B2(I37[21]), 
	.Z(O18[21])); 
	AO_CELL inst_19_21 ( 
	.A1(out_sel[38]), 
	.A2(I38[21]), 
	.B1(out_sel[39]), 
	.B2(I39[21]), 
	.Z(O19[21])); 
	AO_CELL inst_20_21 ( 
	.A1(out_sel[40]), 
	.A2(I40[21]), 
	.B1(out_sel[41]), 
	.B2(I41[21]), 
	.Z(O20[21])); 
	AO_CELL inst_21_21 ( 
	.A1(out_sel[42]), 
	.A2(I42[21]), 
	.B1(out_sel[43]), 
	.B2(I43[21]), 
	.Z(O21[21])); 
	AO_CELL inst_22_21 ( 
	.A1(out_sel[44]), 
	.A2(I44[21]), 
	.B1(out_sel[45]), 
	.B2(I45[21]), 
	.Z(O22[21])); 
	AN_CELL inst_and_21 ( 
	.A1(out_sel[46]), 
	.A2(I46[21]), 
	.Z(O23[21])); 
	AO_CELL inst_0_22 ( 
	.A1(out_sel[0]), 
	.A2(I0[22]), 
	.B1(out_sel[1]), 
	.B2(I1[22]), 
	.Z(O0[22])); 
	AO_CELL inst_1_22 ( 
	.A1(out_sel[2]), 
	.A2(I2[22]), 
	.B1(out_sel[3]), 
	.B2(I3[22]), 
	.Z(O1[22])); 
	AO_CELL inst_2_22 ( 
	.A1(out_sel[4]), 
	.A2(I4[22]), 
	.B1(out_sel[5]), 
	.B2(I5[22]), 
	.Z(O2[22])); 
	AO_CELL inst_3_22 ( 
	.A1(out_sel[6]), 
	.A2(I6[22]), 
	.B1(out_sel[7]), 
	.B2(I7[22]), 
	.Z(O3[22])); 
	AO_CELL inst_4_22 ( 
	.A1(out_sel[8]), 
	.A2(I8[22]), 
	.B1(out_sel[9]), 
	.B2(I9[22]), 
	.Z(O4[22])); 
	AO_CELL inst_5_22 ( 
	.A1(out_sel[10]), 
	.A2(I10[22]), 
	.B1(out_sel[11]), 
	.B2(I11[22]), 
	.Z(O5[22])); 
	AO_CELL inst_6_22 ( 
	.A1(out_sel[12]), 
	.A2(I12[22]), 
	.B1(out_sel[13]), 
	.B2(I13[22]), 
	.Z(O6[22])); 
	AO_CELL inst_7_22 ( 
	.A1(out_sel[14]), 
	.A2(I14[22]), 
	.B1(out_sel[15]), 
	.B2(I15[22]), 
	.Z(O7[22])); 
	AO_CELL inst_8_22 ( 
	.A1(out_sel[16]), 
	.A2(I16[22]), 
	.B1(out_sel[17]), 
	.B2(I17[22]), 
	.Z(O8[22])); 
	AO_CELL inst_9_22 ( 
	.A1(out_sel[18]), 
	.A2(I18[22]), 
	.B1(out_sel[19]), 
	.B2(I19[22]), 
	.Z(O9[22])); 
	AO_CELL inst_10_22 ( 
	.A1(out_sel[20]), 
	.A2(I20[22]), 
	.B1(out_sel[21]), 
	.B2(I21[22]), 
	.Z(O10[22])); 
	AO_CELL inst_11_22 ( 
	.A1(out_sel[22]), 
	.A2(I22[22]), 
	.B1(out_sel[23]), 
	.B2(I23[22]), 
	.Z(O11[22])); 
	AO_CELL inst_12_22 ( 
	.A1(out_sel[24]), 
	.A2(I24[22]), 
	.B1(out_sel[25]), 
	.B2(I25[22]), 
	.Z(O12[22])); 
	AO_CELL inst_13_22 ( 
	.A1(out_sel[26]), 
	.A2(I26[22]), 
	.B1(out_sel[27]), 
	.B2(I27[22]), 
	.Z(O13[22])); 
	AO_CELL inst_14_22 ( 
	.A1(out_sel[28]), 
	.A2(I28[22]), 
	.B1(out_sel[29]), 
	.B2(I29[22]), 
	.Z(O14[22])); 
	AO_CELL inst_15_22 ( 
	.A1(out_sel[30]), 
	.A2(I30[22]), 
	.B1(out_sel[31]), 
	.B2(I31[22]), 
	.Z(O15[22])); 
	AO_CELL inst_16_22 ( 
	.A1(out_sel[32]), 
	.A2(I32[22]), 
	.B1(out_sel[33]), 
	.B2(I33[22]), 
	.Z(O16[22])); 
	AO_CELL inst_17_22 ( 
	.A1(out_sel[34]), 
	.A2(I34[22]), 
	.B1(out_sel[35]), 
	.B2(I35[22]), 
	.Z(O17[22])); 
	AO_CELL inst_18_22 ( 
	.A1(out_sel[36]), 
	.A2(I36[22]), 
	.B1(out_sel[37]), 
	.B2(I37[22]), 
	.Z(O18[22])); 
	AO_CELL inst_19_22 ( 
	.A1(out_sel[38]), 
	.A2(I38[22]), 
	.B1(out_sel[39]), 
	.B2(I39[22]), 
	.Z(O19[22])); 
	AO_CELL inst_20_22 ( 
	.A1(out_sel[40]), 
	.A2(I40[22]), 
	.B1(out_sel[41]), 
	.B2(I41[22]), 
	.Z(O20[22])); 
	AO_CELL inst_21_22 ( 
	.A1(out_sel[42]), 
	.A2(I42[22]), 
	.B1(out_sel[43]), 
	.B2(I43[22]), 
	.Z(O21[22])); 
	AO_CELL inst_22_22 ( 
	.A1(out_sel[44]), 
	.A2(I44[22]), 
	.B1(out_sel[45]), 
	.B2(I45[22]), 
	.Z(O22[22])); 
	AN_CELL inst_and_22 ( 
	.A1(out_sel[46]), 
	.A2(I46[22]), 
	.Z(O23[22])); 
	AO_CELL inst_0_23 ( 
	.A1(out_sel[0]), 
	.A2(I0[23]), 
	.B1(out_sel[1]), 
	.B2(I1[23]), 
	.Z(O0[23])); 
	AO_CELL inst_1_23 ( 
	.A1(out_sel[2]), 
	.A2(I2[23]), 
	.B1(out_sel[3]), 
	.B2(I3[23]), 
	.Z(O1[23])); 
	AO_CELL inst_2_23 ( 
	.A1(out_sel[4]), 
	.A2(I4[23]), 
	.B1(out_sel[5]), 
	.B2(I5[23]), 
	.Z(O2[23])); 
	AO_CELL inst_3_23 ( 
	.A1(out_sel[6]), 
	.A2(I6[23]), 
	.B1(out_sel[7]), 
	.B2(I7[23]), 
	.Z(O3[23])); 
	AO_CELL inst_4_23 ( 
	.A1(out_sel[8]), 
	.A2(I8[23]), 
	.B1(out_sel[9]), 
	.B2(I9[23]), 
	.Z(O4[23])); 
	AO_CELL inst_5_23 ( 
	.A1(out_sel[10]), 
	.A2(I10[23]), 
	.B1(out_sel[11]), 
	.B2(I11[23]), 
	.Z(O5[23])); 
	AO_CELL inst_6_23 ( 
	.A1(out_sel[12]), 
	.A2(I12[23]), 
	.B1(out_sel[13]), 
	.B2(I13[23]), 
	.Z(O6[23])); 
	AO_CELL inst_7_23 ( 
	.A1(out_sel[14]), 
	.A2(I14[23]), 
	.B1(out_sel[15]), 
	.B2(I15[23]), 
	.Z(O7[23])); 
	AO_CELL inst_8_23 ( 
	.A1(out_sel[16]), 
	.A2(I16[23]), 
	.B1(out_sel[17]), 
	.B2(I17[23]), 
	.Z(O8[23])); 
	AO_CELL inst_9_23 ( 
	.A1(out_sel[18]), 
	.A2(I18[23]), 
	.B1(out_sel[19]), 
	.B2(I19[23]), 
	.Z(O9[23])); 
	AO_CELL inst_10_23 ( 
	.A1(out_sel[20]), 
	.A2(I20[23]), 
	.B1(out_sel[21]), 
	.B2(I21[23]), 
	.Z(O10[23])); 
	AO_CELL inst_11_23 ( 
	.A1(out_sel[22]), 
	.A2(I22[23]), 
	.B1(out_sel[23]), 
	.B2(I23[23]), 
	.Z(O11[23])); 
	AO_CELL inst_12_23 ( 
	.A1(out_sel[24]), 
	.A2(I24[23]), 
	.B1(out_sel[25]), 
	.B2(I25[23]), 
	.Z(O12[23])); 
	AO_CELL inst_13_23 ( 
	.A1(out_sel[26]), 
	.A2(I26[23]), 
	.B1(out_sel[27]), 
	.B2(I27[23]), 
	.Z(O13[23])); 
	AO_CELL inst_14_23 ( 
	.A1(out_sel[28]), 
	.A2(I28[23]), 
	.B1(out_sel[29]), 
	.B2(I29[23]), 
	.Z(O14[23])); 
	AO_CELL inst_15_23 ( 
	.A1(out_sel[30]), 
	.A2(I30[23]), 
	.B1(out_sel[31]), 
	.B2(I31[23]), 
	.Z(O15[23])); 
	AO_CELL inst_16_23 ( 
	.A1(out_sel[32]), 
	.A2(I32[23]), 
	.B1(out_sel[33]), 
	.B2(I33[23]), 
	.Z(O16[23])); 
	AO_CELL inst_17_23 ( 
	.A1(out_sel[34]), 
	.A2(I34[23]), 
	.B1(out_sel[35]), 
	.B2(I35[23]), 
	.Z(O17[23])); 
	AO_CELL inst_18_23 ( 
	.A1(out_sel[36]), 
	.A2(I36[23]), 
	.B1(out_sel[37]), 
	.B2(I37[23]), 
	.Z(O18[23])); 
	AO_CELL inst_19_23 ( 
	.A1(out_sel[38]), 
	.A2(I38[23]), 
	.B1(out_sel[39]), 
	.B2(I39[23]), 
	.Z(O19[23])); 
	AO_CELL inst_20_23 ( 
	.A1(out_sel[40]), 
	.A2(I40[23]), 
	.B1(out_sel[41]), 
	.B2(I41[23]), 
	.Z(O20[23])); 
	AO_CELL inst_21_23 ( 
	.A1(out_sel[42]), 
	.A2(I42[23]), 
	.B1(out_sel[43]), 
	.B2(I43[23]), 
	.Z(O21[23])); 
	AO_CELL inst_22_23 ( 
	.A1(out_sel[44]), 
	.A2(I44[23]), 
	.B1(out_sel[45]), 
	.B2(I45[23]), 
	.Z(O22[23])); 
	AN_CELL inst_and_23 ( 
	.A1(out_sel[46]), 
	.A2(I46[23]), 
	.Z(O23[23])); 
	AO_CELL inst_0_24 ( 
	.A1(out_sel[0]), 
	.A2(I0[24]), 
	.B1(out_sel[1]), 
	.B2(I1[24]), 
	.Z(O0[24])); 
	AO_CELL inst_1_24 ( 
	.A1(out_sel[2]), 
	.A2(I2[24]), 
	.B1(out_sel[3]), 
	.B2(I3[24]), 
	.Z(O1[24])); 
	AO_CELL inst_2_24 ( 
	.A1(out_sel[4]), 
	.A2(I4[24]), 
	.B1(out_sel[5]), 
	.B2(I5[24]), 
	.Z(O2[24])); 
	AO_CELL inst_3_24 ( 
	.A1(out_sel[6]), 
	.A2(I6[24]), 
	.B1(out_sel[7]), 
	.B2(I7[24]), 
	.Z(O3[24])); 
	AO_CELL inst_4_24 ( 
	.A1(out_sel[8]), 
	.A2(I8[24]), 
	.B1(out_sel[9]), 
	.B2(I9[24]), 
	.Z(O4[24])); 
	AO_CELL inst_5_24 ( 
	.A1(out_sel[10]), 
	.A2(I10[24]), 
	.B1(out_sel[11]), 
	.B2(I11[24]), 
	.Z(O5[24])); 
	AO_CELL inst_6_24 ( 
	.A1(out_sel[12]), 
	.A2(I12[24]), 
	.B1(out_sel[13]), 
	.B2(I13[24]), 
	.Z(O6[24])); 
	AO_CELL inst_7_24 ( 
	.A1(out_sel[14]), 
	.A2(I14[24]), 
	.B1(out_sel[15]), 
	.B2(I15[24]), 
	.Z(O7[24])); 
	AO_CELL inst_8_24 ( 
	.A1(out_sel[16]), 
	.A2(I16[24]), 
	.B1(out_sel[17]), 
	.B2(I17[24]), 
	.Z(O8[24])); 
	AO_CELL inst_9_24 ( 
	.A1(out_sel[18]), 
	.A2(I18[24]), 
	.B1(out_sel[19]), 
	.B2(I19[24]), 
	.Z(O9[24])); 
	AO_CELL inst_10_24 ( 
	.A1(out_sel[20]), 
	.A2(I20[24]), 
	.B1(out_sel[21]), 
	.B2(I21[24]), 
	.Z(O10[24])); 
	AO_CELL inst_11_24 ( 
	.A1(out_sel[22]), 
	.A2(I22[24]), 
	.B1(out_sel[23]), 
	.B2(I23[24]), 
	.Z(O11[24])); 
	AO_CELL inst_12_24 ( 
	.A1(out_sel[24]), 
	.A2(I24[24]), 
	.B1(out_sel[25]), 
	.B2(I25[24]), 
	.Z(O12[24])); 
	AO_CELL inst_13_24 ( 
	.A1(out_sel[26]), 
	.A2(I26[24]), 
	.B1(out_sel[27]), 
	.B2(I27[24]), 
	.Z(O13[24])); 
	AO_CELL inst_14_24 ( 
	.A1(out_sel[28]), 
	.A2(I28[24]), 
	.B1(out_sel[29]), 
	.B2(I29[24]), 
	.Z(O14[24])); 
	AO_CELL inst_15_24 ( 
	.A1(out_sel[30]), 
	.A2(I30[24]), 
	.B1(out_sel[31]), 
	.B2(I31[24]), 
	.Z(O15[24])); 
	AO_CELL inst_16_24 ( 
	.A1(out_sel[32]), 
	.A2(I32[24]), 
	.B1(out_sel[33]), 
	.B2(I33[24]), 
	.Z(O16[24])); 
	AO_CELL inst_17_24 ( 
	.A1(out_sel[34]), 
	.A2(I34[24]), 
	.B1(out_sel[35]), 
	.B2(I35[24]), 
	.Z(O17[24])); 
	AO_CELL inst_18_24 ( 
	.A1(out_sel[36]), 
	.A2(I36[24]), 
	.B1(out_sel[37]), 
	.B2(I37[24]), 
	.Z(O18[24])); 
	AO_CELL inst_19_24 ( 
	.A1(out_sel[38]), 
	.A2(I38[24]), 
	.B1(out_sel[39]), 
	.B2(I39[24]), 
	.Z(O19[24])); 
	AO_CELL inst_20_24 ( 
	.A1(out_sel[40]), 
	.A2(I40[24]), 
	.B1(out_sel[41]), 
	.B2(I41[24]), 
	.Z(O20[24])); 
	AO_CELL inst_21_24 ( 
	.A1(out_sel[42]), 
	.A2(I42[24]), 
	.B1(out_sel[43]), 
	.B2(I43[24]), 
	.Z(O21[24])); 
	AO_CELL inst_22_24 ( 
	.A1(out_sel[44]), 
	.A2(I44[24]), 
	.B1(out_sel[45]), 
	.B2(I45[24]), 
	.Z(O22[24])); 
	AN_CELL inst_and_24 ( 
	.A1(out_sel[46]), 
	.A2(I46[24]), 
	.Z(O23[24])); 
	AO_CELL inst_0_25 ( 
	.A1(out_sel[0]), 
	.A2(I0[25]), 
	.B1(out_sel[1]), 
	.B2(I1[25]), 
	.Z(O0[25])); 
	AO_CELL inst_1_25 ( 
	.A1(out_sel[2]), 
	.A2(I2[25]), 
	.B1(out_sel[3]), 
	.B2(I3[25]), 
	.Z(O1[25])); 
	AO_CELL inst_2_25 ( 
	.A1(out_sel[4]), 
	.A2(I4[25]), 
	.B1(out_sel[5]), 
	.B2(I5[25]), 
	.Z(O2[25])); 
	AO_CELL inst_3_25 ( 
	.A1(out_sel[6]), 
	.A2(I6[25]), 
	.B1(out_sel[7]), 
	.B2(I7[25]), 
	.Z(O3[25])); 
	AO_CELL inst_4_25 ( 
	.A1(out_sel[8]), 
	.A2(I8[25]), 
	.B1(out_sel[9]), 
	.B2(I9[25]), 
	.Z(O4[25])); 
	AO_CELL inst_5_25 ( 
	.A1(out_sel[10]), 
	.A2(I10[25]), 
	.B1(out_sel[11]), 
	.B2(I11[25]), 
	.Z(O5[25])); 
	AO_CELL inst_6_25 ( 
	.A1(out_sel[12]), 
	.A2(I12[25]), 
	.B1(out_sel[13]), 
	.B2(I13[25]), 
	.Z(O6[25])); 
	AO_CELL inst_7_25 ( 
	.A1(out_sel[14]), 
	.A2(I14[25]), 
	.B1(out_sel[15]), 
	.B2(I15[25]), 
	.Z(O7[25])); 
	AO_CELL inst_8_25 ( 
	.A1(out_sel[16]), 
	.A2(I16[25]), 
	.B1(out_sel[17]), 
	.B2(I17[25]), 
	.Z(O8[25])); 
	AO_CELL inst_9_25 ( 
	.A1(out_sel[18]), 
	.A2(I18[25]), 
	.B1(out_sel[19]), 
	.B2(I19[25]), 
	.Z(O9[25])); 
	AO_CELL inst_10_25 ( 
	.A1(out_sel[20]), 
	.A2(I20[25]), 
	.B1(out_sel[21]), 
	.B2(I21[25]), 
	.Z(O10[25])); 
	AO_CELL inst_11_25 ( 
	.A1(out_sel[22]), 
	.A2(I22[25]), 
	.B1(out_sel[23]), 
	.B2(I23[25]), 
	.Z(O11[25])); 
	AO_CELL inst_12_25 ( 
	.A1(out_sel[24]), 
	.A2(I24[25]), 
	.B1(out_sel[25]), 
	.B2(I25[25]), 
	.Z(O12[25])); 
	AO_CELL inst_13_25 ( 
	.A1(out_sel[26]), 
	.A2(I26[25]), 
	.B1(out_sel[27]), 
	.B2(I27[25]), 
	.Z(O13[25])); 
	AO_CELL inst_14_25 ( 
	.A1(out_sel[28]), 
	.A2(I28[25]), 
	.B1(out_sel[29]), 
	.B2(I29[25]), 
	.Z(O14[25])); 
	AO_CELL inst_15_25 ( 
	.A1(out_sel[30]), 
	.A2(I30[25]), 
	.B1(out_sel[31]), 
	.B2(I31[25]), 
	.Z(O15[25])); 
	AO_CELL inst_16_25 ( 
	.A1(out_sel[32]), 
	.A2(I32[25]), 
	.B1(out_sel[33]), 
	.B2(I33[25]), 
	.Z(O16[25])); 
	AO_CELL inst_17_25 ( 
	.A1(out_sel[34]), 
	.A2(I34[25]), 
	.B1(out_sel[35]), 
	.B2(I35[25]), 
	.Z(O17[25])); 
	AO_CELL inst_18_25 ( 
	.A1(out_sel[36]), 
	.A2(I36[25]), 
	.B1(out_sel[37]), 
	.B2(I37[25]), 
	.Z(O18[25])); 
	AO_CELL inst_19_25 ( 
	.A1(out_sel[38]), 
	.A2(I38[25]), 
	.B1(out_sel[39]), 
	.B2(I39[25]), 
	.Z(O19[25])); 
	AO_CELL inst_20_25 ( 
	.A1(out_sel[40]), 
	.A2(I40[25]), 
	.B1(out_sel[41]), 
	.B2(I41[25]), 
	.Z(O20[25])); 
	AO_CELL inst_21_25 ( 
	.A1(out_sel[42]), 
	.A2(I42[25]), 
	.B1(out_sel[43]), 
	.B2(I43[25]), 
	.Z(O21[25])); 
	AO_CELL inst_22_25 ( 
	.A1(out_sel[44]), 
	.A2(I44[25]), 
	.B1(out_sel[45]), 
	.B2(I45[25]), 
	.Z(O22[25])); 
	AN_CELL inst_and_25 ( 
	.A1(out_sel[46]), 
	.A2(I46[25]), 
	.Z(O23[25])); 
	AO_CELL inst_0_26 ( 
	.A1(out_sel[0]), 
	.A2(I0[26]), 
	.B1(out_sel[1]), 
	.B2(I1[26]), 
	.Z(O0[26])); 
	AO_CELL inst_1_26 ( 
	.A1(out_sel[2]), 
	.A2(I2[26]), 
	.B1(out_sel[3]), 
	.B2(I3[26]), 
	.Z(O1[26])); 
	AO_CELL inst_2_26 ( 
	.A1(out_sel[4]), 
	.A2(I4[26]), 
	.B1(out_sel[5]), 
	.B2(I5[26]), 
	.Z(O2[26])); 
	AO_CELL inst_3_26 ( 
	.A1(out_sel[6]), 
	.A2(I6[26]), 
	.B1(out_sel[7]), 
	.B2(I7[26]), 
	.Z(O3[26])); 
	AO_CELL inst_4_26 ( 
	.A1(out_sel[8]), 
	.A2(I8[26]), 
	.B1(out_sel[9]), 
	.B2(I9[26]), 
	.Z(O4[26])); 
	AO_CELL inst_5_26 ( 
	.A1(out_sel[10]), 
	.A2(I10[26]), 
	.B1(out_sel[11]), 
	.B2(I11[26]), 
	.Z(O5[26])); 
	AO_CELL inst_6_26 ( 
	.A1(out_sel[12]), 
	.A2(I12[26]), 
	.B1(out_sel[13]), 
	.B2(I13[26]), 
	.Z(O6[26])); 
	AO_CELL inst_7_26 ( 
	.A1(out_sel[14]), 
	.A2(I14[26]), 
	.B1(out_sel[15]), 
	.B2(I15[26]), 
	.Z(O7[26])); 
	AO_CELL inst_8_26 ( 
	.A1(out_sel[16]), 
	.A2(I16[26]), 
	.B1(out_sel[17]), 
	.B2(I17[26]), 
	.Z(O8[26])); 
	AO_CELL inst_9_26 ( 
	.A1(out_sel[18]), 
	.A2(I18[26]), 
	.B1(out_sel[19]), 
	.B2(I19[26]), 
	.Z(O9[26])); 
	AO_CELL inst_10_26 ( 
	.A1(out_sel[20]), 
	.A2(I20[26]), 
	.B1(out_sel[21]), 
	.B2(I21[26]), 
	.Z(O10[26])); 
	AO_CELL inst_11_26 ( 
	.A1(out_sel[22]), 
	.A2(I22[26]), 
	.B1(out_sel[23]), 
	.B2(I23[26]), 
	.Z(O11[26])); 
	AO_CELL inst_12_26 ( 
	.A1(out_sel[24]), 
	.A2(I24[26]), 
	.B1(out_sel[25]), 
	.B2(I25[26]), 
	.Z(O12[26])); 
	AO_CELL inst_13_26 ( 
	.A1(out_sel[26]), 
	.A2(I26[26]), 
	.B1(out_sel[27]), 
	.B2(I27[26]), 
	.Z(O13[26])); 
	AO_CELL inst_14_26 ( 
	.A1(out_sel[28]), 
	.A2(I28[26]), 
	.B1(out_sel[29]), 
	.B2(I29[26]), 
	.Z(O14[26])); 
	AO_CELL inst_15_26 ( 
	.A1(out_sel[30]), 
	.A2(I30[26]), 
	.B1(out_sel[31]), 
	.B2(I31[26]), 
	.Z(O15[26])); 
	AO_CELL inst_16_26 ( 
	.A1(out_sel[32]), 
	.A2(I32[26]), 
	.B1(out_sel[33]), 
	.B2(I33[26]), 
	.Z(O16[26])); 
	AO_CELL inst_17_26 ( 
	.A1(out_sel[34]), 
	.A2(I34[26]), 
	.B1(out_sel[35]), 
	.B2(I35[26]), 
	.Z(O17[26])); 
	AO_CELL inst_18_26 ( 
	.A1(out_sel[36]), 
	.A2(I36[26]), 
	.B1(out_sel[37]), 
	.B2(I37[26]), 
	.Z(O18[26])); 
	AO_CELL inst_19_26 ( 
	.A1(out_sel[38]), 
	.A2(I38[26]), 
	.B1(out_sel[39]), 
	.B2(I39[26]), 
	.Z(O19[26])); 
	AO_CELL inst_20_26 ( 
	.A1(out_sel[40]), 
	.A2(I40[26]), 
	.B1(out_sel[41]), 
	.B2(I41[26]), 
	.Z(O20[26])); 
	AO_CELL inst_21_26 ( 
	.A1(out_sel[42]), 
	.A2(I42[26]), 
	.B1(out_sel[43]), 
	.B2(I43[26]), 
	.Z(O21[26])); 
	AO_CELL inst_22_26 ( 
	.A1(out_sel[44]), 
	.A2(I44[26]), 
	.B1(out_sel[45]), 
	.B2(I45[26]), 
	.Z(O22[26])); 
	AN_CELL inst_and_26 ( 
	.A1(out_sel[46]), 
	.A2(I46[26]), 
	.Z(O23[26])); 
	AO_CELL inst_0_27 ( 
	.A1(out_sel[0]), 
	.A2(I0[27]), 
	.B1(out_sel[1]), 
	.B2(I1[27]), 
	.Z(O0[27])); 
	AO_CELL inst_1_27 ( 
	.A1(out_sel[2]), 
	.A2(I2[27]), 
	.B1(out_sel[3]), 
	.B2(I3[27]), 
	.Z(O1[27])); 
	AO_CELL inst_2_27 ( 
	.A1(out_sel[4]), 
	.A2(I4[27]), 
	.B1(out_sel[5]), 
	.B2(I5[27]), 
	.Z(O2[27])); 
	AO_CELL inst_3_27 ( 
	.A1(out_sel[6]), 
	.A2(I6[27]), 
	.B1(out_sel[7]), 
	.B2(I7[27]), 
	.Z(O3[27])); 
	AO_CELL inst_4_27 ( 
	.A1(out_sel[8]), 
	.A2(I8[27]), 
	.B1(out_sel[9]), 
	.B2(I9[27]), 
	.Z(O4[27])); 
	AO_CELL inst_5_27 ( 
	.A1(out_sel[10]), 
	.A2(I10[27]), 
	.B1(out_sel[11]), 
	.B2(I11[27]), 
	.Z(O5[27])); 
	AO_CELL inst_6_27 ( 
	.A1(out_sel[12]), 
	.A2(I12[27]), 
	.B1(out_sel[13]), 
	.B2(I13[27]), 
	.Z(O6[27])); 
	AO_CELL inst_7_27 ( 
	.A1(out_sel[14]), 
	.A2(I14[27]), 
	.B1(out_sel[15]), 
	.B2(I15[27]), 
	.Z(O7[27])); 
	AO_CELL inst_8_27 ( 
	.A1(out_sel[16]), 
	.A2(I16[27]), 
	.B1(out_sel[17]), 
	.B2(I17[27]), 
	.Z(O8[27])); 
	AO_CELL inst_9_27 ( 
	.A1(out_sel[18]), 
	.A2(I18[27]), 
	.B1(out_sel[19]), 
	.B2(I19[27]), 
	.Z(O9[27])); 
	AO_CELL inst_10_27 ( 
	.A1(out_sel[20]), 
	.A2(I20[27]), 
	.B1(out_sel[21]), 
	.B2(I21[27]), 
	.Z(O10[27])); 
	AO_CELL inst_11_27 ( 
	.A1(out_sel[22]), 
	.A2(I22[27]), 
	.B1(out_sel[23]), 
	.B2(I23[27]), 
	.Z(O11[27])); 
	AO_CELL inst_12_27 ( 
	.A1(out_sel[24]), 
	.A2(I24[27]), 
	.B1(out_sel[25]), 
	.B2(I25[27]), 
	.Z(O12[27])); 
	AO_CELL inst_13_27 ( 
	.A1(out_sel[26]), 
	.A2(I26[27]), 
	.B1(out_sel[27]), 
	.B2(I27[27]), 
	.Z(O13[27])); 
	AO_CELL inst_14_27 ( 
	.A1(out_sel[28]), 
	.A2(I28[27]), 
	.B1(out_sel[29]), 
	.B2(I29[27]), 
	.Z(O14[27])); 
	AO_CELL inst_15_27 ( 
	.A1(out_sel[30]), 
	.A2(I30[27]), 
	.B1(out_sel[31]), 
	.B2(I31[27]), 
	.Z(O15[27])); 
	AO_CELL inst_16_27 ( 
	.A1(out_sel[32]), 
	.A2(I32[27]), 
	.B1(out_sel[33]), 
	.B2(I33[27]), 
	.Z(O16[27])); 
	AO_CELL inst_17_27 ( 
	.A1(out_sel[34]), 
	.A2(I34[27]), 
	.B1(out_sel[35]), 
	.B2(I35[27]), 
	.Z(O17[27])); 
	AO_CELL inst_18_27 ( 
	.A1(out_sel[36]), 
	.A2(I36[27]), 
	.B1(out_sel[37]), 
	.B2(I37[27]), 
	.Z(O18[27])); 
	AO_CELL inst_19_27 ( 
	.A1(out_sel[38]), 
	.A2(I38[27]), 
	.B1(out_sel[39]), 
	.B2(I39[27]), 
	.Z(O19[27])); 
	AO_CELL inst_20_27 ( 
	.A1(out_sel[40]), 
	.A2(I40[27]), 
	.B1(out_sel[41]), 
	.B2(I41[27]), 
	.Z(O20[27])); 
	AO_CELL inst_21_27 ( 
	.A1(out_sel[42]), 
	.A2(I42[27]), 
	.B1(out_sel[43]), 
	.B2(I43[27]), 
	.Z(O21[27])); 
	AO_CELL inst_22_27 ( 
	.A1(out_sel[44]), 
	.A2(I44[27]), 
	.B1(out_sel[45]), 
	.B2(I45[27]), 
	.Z(O22[27])); 
	AN_CELL inst_and_27 ( 
	.A1(out_sel[46]), 
	.A2(I46[27]), 
	.Z(O23[27])); 
	AO_CELL inst_0_28 ( 
	.A1(out_sel[0]), 
	.A2(I0[28]), 
	.B1(out_sel[1]), 
	.B2(I1[28]), 
	.Z(O0[28])); 
	AO_CELL inst_1_28 ( 
	.A1(out_sel[2]), 
	.A2(I2[28]), 
	.B1(out_sel[3]), 
	.B2(I3[28]), 
	.Z(O1[28])); 
	AO_CELL inst_2_28 ( 
	.A1(out_sel[4]), 
	.A2(I4[28]), 
	.B1(out_sel[5]), 
	.B2(I5[28]), 
	.Z(O2[28])); 
	AO_CELL inst_3_28 ( 
	.A1(out_sel[6]), 
	.A2(I6[28]), 
	.B1(out_sel[7]), 
	.B2(I7[28]), 
	.Z(O3[28])); 
	AO_CELL inst_4_28 ( 
	.A1(out_sel[8]), 
	.A2(I8[28]), 
	.B1(out_sel[9]), 
	.B2(I9[28]), 
	.Z(O4[28])); 
	AO_CELL inst_5_28 ( 
	.A1(out_sel[10]), 
	.A2(I10[28]), 
	.B1(out_sel[11]), 
	.B2(I11[28]), 
	.Z(O5[28])); 
	AO_CELL inst_6_28 ( 
	.A1(out_sel[12]), 
	.A2(I12[28]), 
	.B1(out_sel[13]), 
	.B2(I13[28]), 
	.Z(O6[28])); 
	AO_CELL inst_7_28 ( 
	.A1(out_sel[14]), 
	.A2(I14[28]), 
	.B1(out_sel[15]), 
	.B2(I15[28]), 
	.Z(O7[28])); 
	AO_CELL inst_8_28 ( 
	.A1(out_sel[16]), 
	.A2(I16[28]), 
	.B1(out_sel[17]), 
	.B2(I17[28]), 
	.Z(O8[28])); 
	AO_CELL inst_9_28 ( 
	.A1(out_sel[18]), 
	.A2(I18[28]), 
	.B1(out_sel[19]), 
	.B2(I19[28]), 
	.Z(O9[28])); 
	AO_CELL inst_10_28 ( 
	.A1(out_sel[20]), 
	.A2(I20[28]), 
	.B1(out_sel[21]), 
	.B2(I21[28]), 
	.Z(O10[28])); 
	AO_CELL inst_11_28 ( 
	.A1(out_sel[22]), 
	.A2(I22[28]), 
	.B1(out_sel[23]), 
	.B2(I23[28]), 
	.Z(O11[28])); 
	AO_CELL inst_12_28 ( 
	.A1(out_sel[24]), 
	.A2(I24[28]), 
	.B1(out_sel[25]), 
	.B2(I25[28]), 
	.Z(O12[28])); 
	AO_CELL inst_13_28 ( 
	.A1(out_sel[26]), 
	.A2(I26[28]), 
	.B1(out_sel[27]), 
	.B2(I27[28]), 
	.Z(O13[28])); 
	AO_CELL inst_14_28 ( 
	.A1(out_sel[28]), 
	.A2(I28[28]), 
	.B1(out_sel[29]), 
	.B2(I29[28]), 
	.Z(O14[28])); 
	AO_CELL inst_15_28 ( 
	.A1(out_sel[30]), 
	.A2(I30[28]), 
	.B1(out_sel[31]), 
	.B2(I31[28]), 
	.Z(O15[28])); 
	AO_CELL inst_16_28 ( 
	.A1(out_sel[32]), 
	.A2(I32[28]), 
	.B1(out_sel[33]), 
	.B2(I33[28]), 
	.Z(O16[28])); 
	AO_CELL inst_17_28 ( 
	.A1(out_sel[34]), 
	.A2(I34[28]), 
	.B1(out_sel[35]), 
	.B2(I35[28]), 
	.Z(O17[28])); 
	AO_CELL inst_18_28 ( 
	.A1(out_sel[36]), 
	.A2(I36[28]), 
	.B1(out_sel[37]), 
	.B2(I37[28]), 
	.Z(O18[28])); 
	AO_CELL inst_19_28 ( 
	.A1(out_sel[38]), 
	.A2(I38[28]), 
	.B1(out_sel[39]), 
	.B2(I39[28]), 
	.Z(O19[28])); 
	AO_CELL inst_20_28 ( 
	.A1(out_sel[40]), 
	.A2(I40[28]), 
	.B1(out_sel[41]), 
	.B2(I41[28]), 
	.Z(O20[28])); 
	AO_CELL inst_21_28 ( 
	.A1(out_sel[42]), 
	.A2(I42[28]), 
	.B1(out_sel[43]), 
	.B2(I43[28]), 
	.Z(O21[28])); 
	AO_CELL inst_22_28 ( 
	.A1(out_sel[44]), 
	.A2(I44[28]), 
	.B1(out_sel[45]), 
	.B2(I45[28]), 
	.Z(O22[28])); 
	AN_CELL inst_and_28 ( 
	.A1(out_sel[46]), 
	.A2(I46[28]), 
	.Z(O23[28])); 
	AO_CELL inst_0_29 ( 
	.A1(out_sel[0]), 
	.A2(I0[29]), 
	.B1(out_sel[1]), 
	.B2(I1[29]), 
	.Z(O0[29])); 
	AO_CELL inst_1_29 ( 
	.A1(out_sel[2]), 
	.A2(I2[29]), 
	.B1(out_sel[3]), 
	.B2(I3[29]), 
	.Z(O1[29])); 
	AO_CELL inst_2_29 ( 
	.A1(out_sel[4]), 
	.A2(I4[29]), 
	.B1(out_sel[5]), 
	.B2(I5[29]), 
	.Z(O2[29])); 
	AO_CELL inst_3_29 ( 
	.A1(out_sel[6]), 
	.A2(I6[29]), 
	.B1(out_sel[7]), 
	.B2(I7[29]), 
	.Z(O3[29])); 
	AO_CELL inst_4_29 ( 
	.A1(out_sel[8]), 
	.A2(I8[29]), 
	.B1(out_sel[9]), 
	.B2(I9[29]), 
	.Z(O4[29])); 
	AO_CELL inst_5_29 ( 
	.A1(out_sel[10]), 
	.A2(I10[29]), 
	.B1(out_sel[11]), 
	.B2(I11[29]), 
	.Z(O5[29])); 
	AO_CELL inst_6_29 ( 
	.A1(out_sel[12]), 
	.A2(I12[29]), 
	.B1(out_sel[13]), 
	.B2(I13[29]), 
	.Z(O6[29])); 
	AO_CELL inst_7_29 ( 
	.A1(out_sel[14]), 
	.A2(I14[29]), 
	.B1(out_sel[15]), 
	.B2(I15[29]), 
	.Z(O7[29])); 
	AO_CELL inst_8_29 ( 
	.A1(out_sel[16]), 
	.A2(I16[29]), 
	.B1(out_sel[17]), 
	.B2(I17[29]), 
	.Z(O8[29])); 
	AO_CELL inst_9_29 ( 
	.A1(out_sel[18]), 
	.A2(I18[29]), 
	.B1(out_sel[19]), 
	.B2(I19[29]), 
	.Z(O9[29])); 
	AO_CELL inst_10_29 ( 
	.A1(out_sel[20]), 
	.A2(I20[29]), 
	.B1(out_sel[21]), 
	.B2(I21[29]), 
	.Z(O10[29])); 
	AO_CELL inst_11_29 ( 
	.A1(out_sel[22]), 
	.A2(I22[29]), 
	.B1(out_sel[23]), 
	.B2(I23[29]), 
	.Z(O11[29])); 
	AO_CELL inst_12_29 ( 
	.A1(out_sel[24]), 
	.A2(I24[29]), 
	.B1(out_sel[25]), 
	.B2(I25[29]), 
	.Z(O12[29])); 
	AO_CELL inst_13_29 ( 
	.A1(out_sel[26]), 
	.A2(I26[29]), 
	.B1(out_sel[27]), 
	.B2(I27[29]), 
	.Z(O13[29])); 
	AO_CELL inst_14_29 ( 
	.A1(out_sel[28]), 
	.A2(I28[29]), 
	.B1(out_sel[29]), 
	.B2(I29[29]), 
	.Z(O14[29])); 
	AO_CELL inst_15_29 ( 
	.A1(out_sel[30]), 
	.A2(I30[29]), 
	.B1(out_sel[31]), 
	.B2(I31[29]), 
	.Z(O15[29])); 
	AO_CELL inst_16_29 ( 
	.A1(out_sel[32]), 
	.A2(I32[29]), 
	.B1(out_sel[33]), 
	.B2(I33[29]), 
	.Z(O16[29])); 
	AO_CELL inst_17_29 ( 
	.A1(out_sel[34]), 
	.A2(I34[29]), 
	.B1(out_sel[35]), 
	.B2(I35[29]), 
	.Z(O17[29])); 
	AO_CELL inst_18_29 ( 
	.A1(out_sel[36]), 
	.A2(I36[29]), 
	.B1(out_sel[37]), 
	.B2(I37[29]), 
	.Z(O18[29])); 
	AO_CELL inst_19_29 ( 
	.A1(out_sel[38]), 
	.A2(I38[29]), 
	.B1(out_sel[39]), 
	.B2(I39[29]), 
	.Z(O19[29])); 
	AO_CELL inst_20_29 ( 
	.A1(out_sel[40]), 
	.A2(I40[29]), 
	.B1(out_sel[41]), 
	.B2(I41[29]), 
	.Z(O20[29])); 
	AO_CELL inst_21_29 ( 
	.A1(out_sel[42]), 
	.A2(I42[29]), 
	.B1(out_sel[43]), 
	.B2(I43[29]), 
	.Z(O21[29])); 
	AO_CELL inst_22_29 ( 
	.A1(out_sel[44]), 
	.A2(I44[29]), 
	.B1(out_sel[45]), 
	.B2(I45[29]), 
	.Z(O22[29])); 
	AN_CELL inst_and_29 ( 
	.A1(out_sel[46]), 
	.A2(I46[29]), 
	.Z(O23[29])); 
	AO_CELL inst_0_30 ( 
	.A1(out_sel[0]), 
	.A2(I0[30]), 
	.B1(out_sel[1]), 
	.B2(I1[30]), 
	.Z(O0[30])); 
	AO_CELL inst_1_30 ( 
	.A1(out_sel[2]), 
	.A2(I2[30]), 
	.B1(out_sel[3]), 
	.B2(I3[30]), 
	.Z(O1[30])); 
	AO_CELL inst_2_30 ( 
	.A1(out_sel[4]), 
	.A2(I4[30]), 
	.B1(out_sel[5]), 
	.B2(I5[30]), 
	.Z(O2[30])); 
	AO_CELL inst_3_30 ( 
	.A1(out_sel[6]), 
	.A2(I6[30]), 
	.B1(out_sel[7]), 
	.B2(I7[30]), 
	.Z(O3[30])); 
	AO_CELL inst_4_30 ( 
	.A1(out_sel[8]), 
	.A2(I8[30]), 
	.B1(out_sel[9]), 
	.B2(I9[30]), 
	.Z(O4[30])); 
	AO_CELL inst_5_30 ( 
	.A1(out_sel[10]), 
	.A2(I10[30]), 
	.B1(out_sel[11]), 
	.B2(I11[30]), 
	.Z(O5[30])); 
	AO_CELL inst_6_30 ( 
	.A1(out_sel[12]), 
	.A2(I12[30]), 
	.B1(out_sel[13]), 
	.B2(I13[30]), 
	.Z(O6[30])); 
	AO_CELL inst_7_30 ( 
	.A1(out_sel[14]), 
	.A2(I14[30]), 
	.B1(out_sel[15]), 
	.B2(I15[30]), 
	.Z(O7[30])); 
	AO_CELL inst_8_30 ( 
	.A1(out_sel[16]), 
	.A2(I16[30]), 
	.B1(out_sel[17]), 
	.B2(I17[30]), 
	.Z(O8[30])); 
	AO_CELL inst_9_30 ( 
	.A1(out_sel[18]), 
	.A2(I18[30]), 
	.B1(out_sel[19]), 
	.B2(I19[30]), 
	.Z(O9[30])); 
	AO_CELL inst_10_30 ( 
	.A1(out_sel[20]), 
	.A2(I20[30]), 
	.B1(out_sel[21]), 
	.B2(I21[30]), 
	.Z(O10[30])); 
	AO_CELL inst_11_30 ( 
	.A1(out_sel[22]), 
	.A2(I22[30]), 
	.B1(out_sel[23]), 
	.B2(I23[30]), 
	.Z(O11[30])); 
	AO_CELL inst_12_30 ( 
	.A1(out_sel[24]), 
	.A2(I24[30]), 
	.B1(out_sel[25]), 
	.B2(I25[30]), 
	.Z(O12[30])); 
	AO_CELL inst_13_30 ( 
	.A1(out_sel[26]), 
	.A2(I26[30]), 
	.B1(out_sel[27]), 
	.B2(I27[30]), 
	.Z(O13[30])); 
	AO_CELL inst_14_30 ( 
	.A1(out_sel[28]), 
	.A2(I28[30]), 
	.B1(out_sel[29]), 
	.B2(I29[30]), 
	.Z(O14[30])); 
	AO_CELL inst_15_30 ( 
	.A1(out_sel[30]), 
	.A2(I30[30]), 
	.B1(out_sel[31]), 
	.B2(I31[30]), 
	.Z(O15[30])); 
	AO_CELL inst_16_30 ( 
	.A1(out_sel[32]), 
	.A2(I32[30]), 
	.B1(out_sel[33]), 
	.B2(I33[30]), 
	.Z(O16[30])); 
	AO_CELL inst_17_30 ( 
	.A1(out_sel[34]), 
	.A2(I34[30]), 
	.B1(out_sel[35]), 
	.B2(I35[30]), 
	.Z(O17[30])); 
	AO_CELL inst_18_30 ( 
	.A1(out_sel[36]), 
	.A2(I36[30]), 
	.B1(out_sel[37]), 
	.B2(I37[30]), 
	.Z(O18[30])); 
	AO_CELL inst_19_30 ( 
	.A1(out_sel[38]), 
	.A2(I38[30]), 
	.B1(out_sel[39]), 
	.B2(I39[30]), 
	.Z(O19[30])); 
	AO_CELL inst_20_30 ( 
	.A1(out_sel[40]), 
	.A2(I40[30]), 
	.B1(out_sel[41]), 
	.B2(I41[30]), 
	.Z(O20[30])); 
	AO_CELL inst_21_30 ( 
	.A1(out_sel[42]), 
	.A2(I42[30]), 
	.B1(out_sel[43]), 
	.B2(I43[30]), 
	.Z(O21[30])); 
	AO_CELL inst_22_30 ( 
	.A1(out_sel[44]), 
	.A2(I44[30]), 
	.B1(out_sel[45]), 
	.B2(I45[30]), 
	.Z(O22[30])); 
	AN_CELL inst_and_30 ( 
	.A1(out_sel[46]), 
	.A2(I46[30]), 
	.Z(O23[30])); 
	AO_CELL inst_0_31 ( 
	.A1(out_sel[0]), 
	.A2(I0[31]), 
	.B1(out_sel[1]), 
	.B2(I1[31]), 
	.Z(O0[31])); 
	AO_CELL inst_1_31 ( 
	.A1(out_sel[2]), 
	.A2(I2[31]), 
	.B1(out_sel[3]), 
	.B2(I3[31]), 
	.Z(O1[31])); 
	AO_CELL inst_2_31 ( 
	.A1(out_sel[4]), 
	.A2(I4[31]), 
	.B1(out_sel[5]), 
	.B2(I5[31]), 
	.Z(O2[31])); 
	AO_CELL inst_3_31 ( 
	.A1(out_sel[6]), 
	.A2(I6[31]), 
	.B1(out_sel[7]), 
	.B2(I7[31]), 
	.Z(O3[31])); 
	AO_CELL inst_4_31 ( 
	.A1(out_sel[8]), 
	.A2(I8[31]), 
	.B1(out_sel[9]), 
	.B2(I9[31]), 
	.Z(O4[31])); 
	AO_CELL inst_5_31 ( 
	.A1(out_sel[10]), 
	.A2(I10[31]), 
	.B1(out_sel[11]), 
	.B2(I11[31]), 
	.Z(O5[31])); 
	AO_CELL inst_6_31 ( 
	.A1(out_sel[12]), 
	.A2(I12[31]), 
	.B1(out_sel[13]), 
	.B2(I13[31]), 
	.Z(O6[31])); 
	AO_CELL inst_7_31 ( 
	.A1(out_sel[14]), 
	.A2(I14[31]), 
	.B1(out_sel[15]), 
	.B2(I15[31]), 
	.Z(O7[31])); 
	AO_CELL inst_8_31 ( 
	.A1(out_sel[16]), 
	.A2(I16[31]), 
	.B1(out_sel[17]), 
	.B2(I17[31]), 
	.Z(O8[31])); 
	AO_CELL inst_9_31 ( 
	.A1(out_sel[18]), 
	.A2(I18[31]), 
	.B1(out_sel[19]), 
	.B2(I19[31]), 
	.Z(O9[31])); 
	AO_CELL inst_10_31 ( 
	.A1(out_sel[20]), 
	.A2(I20[31]), 
	.B1(out_sel[21]), 
	.B2(I21[31]), 
	.Z(O10[31])); 
	AO_CELL inst_11_31 ( 
	.A1(out_sel[22]), 
	.A2(I22[31]), 
	.B1(out_sel[23]), 
	.B2(I23[31]), 
	.Z(O11[31])); 
	AO_CELL inst_12_31 ( 
	.A1(out_sel[24]), 
	.A2(I24[31]), 
	.B1(out_sel[25]), 
	.B2(I25[31]), 
	.Z(O12[31])); 
	AO_CELL inst_13_31 ( 
	.A1(out_sel[26]), 
	.A2(I26[31]), 
	.B1(out_sel[27]), 
	.B2(I27[31]), 
	.Z(O13[31])); 
	AO_CELL inst_14_31 ( 
	.A1(out_sel[28]), 
	.A2(I28[31]), 
	.B1(out_sel[29]), 
	.B2(I29[31]), 
	.Z(O14[31])); 
	AO_CELL inst_15_31 ( 
	.A1(out_sel[30]), 
	.A2(I30[31]), 
	.B1(out_sel[31]), 
	.B2(I31[31]), 
	.Z(O15[31])); 
	AO_CELL inst_16_31 ( 
	.A1(out_sel[32]), 
	.A2(I32[31]), 
	.B1(out_sel[33]), 
	.B2(I33[31]), 
	.Z(O16[31])); 
	AO_CELL inst_17_31 ( 
	.A1(out_sel[34]), 
	.A2(I34[31]), 
	.B1(out_sel[35]), 
	.B2(I35[31]), 
	.Z(O17[31])); 
	AO_CELL inst_18_31 ( 
	.A1(out_sel[36]), 
	.A2(I36[31]), 
	.B1(out_sel[37]), 
	.B2(I37[31]), 
	.Z(O18[31])); 
	AO_CELL inst_19_31 ( 
	.A1(out_sel[38]), 
	.A2(I38[31]), 
	.B1(out_sel[39]), 
	.B2(I39[31]), 
	.Z(O19[31])); 
	AO_CELL inst_20_31 ( 
	.A1(out_sel[40]), 
	.A2(I40[31]), 
	.B1(out_sel[41]), 
	.B2(I41[31]), 
	.Z(O20[31])); 
	AO_CELL inst_21_31 ( 
	.A1(out_sel[42]), 
	.A2(I42[31]), 
	.B1(out_sel[43]), 
	.B2(I43[31]), 
	.Z(O21[31])); 
	AO_CELL inst_22_31 ( 
	.A1(out_sel[44]), 
	.A2(I44[31]), 
	.B1(out_sel[45]), 
	.B2(I45[31]), 
	.Z(O22[31])); 
	AN_CELL inst_and_31 ( 
	.A1(out_sel[46]), 
	.A2(I46[31]), 
	.Z(O23[31])); 
endmodule 

module mux_aoi_2_32 ( 
	input logic  [31 : 0] I[1:0], 
input logic S, 
	output logic  [1 : 0] out_sel,
	output logic [31 : 0] O); 
	logic  [31 : 0] O_int0;

precoder_32_2 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_32_2 u_mux_logic ( 
	.I0 (I[0]),
	.I1 (I[1]),
	.out_sel(out_sel), 
	.O0(O_int0)); 
	assign O = (  	O_int0 	); 

endmodule 

module precoder_32_2 (
	input logic  [0 : 0] S ,
	output logic  [1 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		1'd0    :   out_sel = 2'b01;
		1'd1    :   out_sel = 2'b10;
		default :   out_sel = 2'b0;
	endcase 
end 

endmodule 

module mux_logic_32_2 ( 
	input logic  [1 : 0] out_sel,
	input logic  [31 : 0] I0, 
	input logic  [31 : 0] I1, 
	output logic  [31 : 0] O0); 
	AO_CELL inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	AO_CELL inst_0_1 ( 
	.A1(out_sel[0]), 
	.A2(I0[1]), 
	.B1(out_sel[1]), 
	.B2(I1[1]), 
	.Z(O0[1])); 
	AO_CELL inst_0_2 ( 
	.A1(out_sel[0]), 
	.A2(I0[2]), 
	.B1(out_sel[1]), 
	.B2(I1[2]), 
	.Z(O0[2])); 
	AO_CELL inst_0_3 ( 
	.A1(out_sel[0]), 
	.A2(I0[3]), 
	.B1(out_sel[1]), 
	.B2(I1[3]), 
	.Z(O0[3])); 
	AO_CELL inst_0_4 ( 
	.A1(out_sel[0]), 
	.A2(I0[4]), 
	.B1(out_sel[1]), 
	.B2(I1[4]), 
	.Z(O0[4])); 
	AO_CELL inst_0_5 ( 
	.A1(out_sel[0]), 
	.A2(I0[5]), 
	.B1(out_sel[1]), 
	.B2(I1[5]), 
	.Z(O0[5])); 
	AO_CELL inst_0_6 ( 
	.A1(out_sel[0]), 
	.A2(I0[6]), 
	.B1(out_sel[1]), 
	.B2(I1[6]), 
	.Z(O0[6])); 
	AO_CELL inst_0_7 ( 
	.A1(out_sel[0]), 
	.A2(I0[7]), 
	.B1(out_sel[1]), 
	.B2(I1[7]), 
	.Z(O0[7])); 
	AO_CELL inst_0_8 ( 
	.A1(out_sel[0]), 
	.A2(I0[8]), 
	.B1(out_sel[1]), 
	.B2(I1[8]), 
	.Z(O0[8])); 
	AO_CELL inst_0_9 ( 
	.A1(out_sel[0]), 
	.A2(I0[9]), 
	.B1(out_sel[1]), 
	.B2(I1[9]), 
	.Z(O0[9])); 
	AO_CELL inst_0_10 ( 
	.A1(out_sel[0]), 
	.A2(I0[10]), 
	.B1(out_sel[1]), 
	.B2(I1[10]), 
	.Z(O0[10])); 
	AO_CELL inst_0_11 ( 
	.A1(out_sel[0]), 
	.A2(I0[11]), 
	.B1(out_sel[1]), 
	.B2(I1[11]), 
	.Z(O0[11])); 
	AO_CELL inst_0_12 ( 
	.A1(out_sel[0]), 
	.A2(I0[12]), 
	.B1(out_sel[1]), 
	.B2(I1[12]), 
	.Z(O0[12])); 
	AO_CELL inst_0_13 ( 
	.A1(out_sel[0]), 
	.A2(I0[13]), 
	.B1(out_sel[1]), 
	.B2(I1[13]), 
	.Z(O0[13])); 
	AO_CELL inst_0_14 ( 
	.A1(out_sel[0]), 
	.A2(I0[14]), 
	.B1(out_sel[1]), 
	.B2(I1[14]), 
	.Z(O0[14])); 
	AO_CELL inst_0_15 ( 
	.A1(out_sel[0]), 
	.A2(I0[15]), 
	.B1(out_sel[1]), 
	.B2(I1[15]), 
	.Z(O0[15])); 
	AO_CELL inst_0_16 ( 
	.A1(out_sel[0]), 
	.A2(I0[16]), 
	.B1(out_sel[1]), 
	.B2(I1[16]), 
	.Z(O0[16])); 
	AO_CELL inst_0_17 ( 
	.A1(out_sel[0]), 
	.A2(I0[17]), 
	.B1(out_sel[1]), 
	.B2(I1[17]), 
	.Z(O0[17])); 
	AO_CELL inst_0_18 ( 
	.A1(out_sel[0]), 
	.A2(I0[18]), 
	.B1(out_sel[1]), 
	.B2(I1[18]), 
	.Z(O0[18])); 
	AO_CELL inst_0_19 ( 
	.A1(out_sel[0]), 
	.A2(I0[19]), 
	.B1(out_sel[1]), 
	.B2(I1[19]), 
	.Z(O0[19])); 
	AO_CELL inst_0_20 ( 
	.A1(out_sel[0]), 
	.A2(I0[20]), 
	.B1(out_sel[1]), 
	.B2(I1[20]), 
	.Z(O0[20])); 
	AO_CELL inst_0_21 ( 
	.A1(out_sel[0]), 
	.A2(I0[21]), 
	.B1(out_sel[1]), 
	.B2(I1[21]), 
	.Z(O0[21])); 
	AO_CELL inst_0_22 ( 
	.A1(out_sel[0]), 
	.A2(I0[22]), 
	.B1(out_sel[1]), 
	.B2(I1[22]), 
	.Z(O0[22])); 
	AO_CELL inst_0_23 ( 
	.A1(out_sel[0]), 
	.A2(I0[23]), 
	.B1(out_sel[1]), 
	.B2(I1[23]), 
	.Z(O0[23])); 
	AO_CELL inst_0_24 ( 
	.A1(out_sel[0]), 
	.A2(I0[24]), 
	.B1(out_sel[1]), 
	.B2(I1[24]), 
	.Z(O0[24])); 
	AO_CELL inst_0_25 ( 
	.A1(out_sel[0]), 
	.A2(I0[25]), 
	.B1(out_sel[1]), 
	.B2(I1[25]), 
	.Z(O0[25])); 
	AO_CELL inst_0_26 ( 
	.A1(out_sel[0]), 
	.A2(I0[26]), 
	.B1(out_sel[1]), 
	.B2(I1[26]), 
	.Z(O0[26])); 
	AO_CELL inst_0_27 ( 
	.A1(out_sel[0]), 
	.A2(I0[27]), 
	.B1(out_sel[1]), 
	.B2(I1[27]), 
	.Z(O0[27])); 
	AO_CELL inst_0_28 ( 
	.A1(out_sel[0]), 
	.A2(I0[28]), 
	.B1(out_sel[1]), 
	.B2(I1[28]), 
	.Z(O0[28])); 
	AO_CELL inst_0_29 ( 
	.A1(out_sel[0]), 
	.A2(I0[29]), 
	.B1(out_sel[1]), 
	.B2(I1[29]), 
	.Z(O0[29])); 
	AO_CELL inst_0_30 ( 
	.A1(out_sel[0]), 
	.A2(I0[30]), 
	.B1(out_sel[1]), 
	.B2(I1[30]), 
	.Z(O0[30])); 
	AO_CELL inst_0_31 ( 
	.A1(out_sel[0]), 
	.A2(I0[31]), 
	.B1(out_sel[1]), 
	.B2(I1[31]), 
	.Z(O0[31])); 
endmodule 

module mux_aoi_18_32 ( 
	input logic  [31 : 0] I[17:0], 
	input logic  [4 : 0] S ,
	output logic  [31 : 0] out_sel,
	output logic [31 : 0] O); 
	logic  [31 : 0] O_int0;
	logic  [31 : 0] O_int1;
	logic  [31 : 0] O_int2;
	logic  [31 : 0] O_int3;
	logic  [31 : 0] O_int4;
	logic  [31 : 0] O_int5;
	logic  [31 : 0] O_int6;
	logic  [31 : 0] O_int7;
	logic  [31 : 0] O_int8;

precoder_32_18 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_32_18 u_mux_logic ( 
	.I0 (I[0]),
	.I1 (I[1]),
	.I2 (I[2]),
	.I3 (I[3]),
	.I4 (I[4]),
	.I5 (I[5]),
	.I6 (I[6]),
	.I7 (I[7]),
	.I8 (I[8]),
	.I9 (I[9]),
	.I10 (I[10]),
	.I11 (I[11]),
	.I12 (I[12]),
	.I13 (I[13]),
	.I14 (I[14]),
	.I15 (I[15]),
	.I16 (I[16]),
	.I17 (I[17]),
	.out_sel(out_sel), 
	.O0(O_int0), 
	.O1(O_int1), 
	.O2(O_int2), 
	.O3(O_int3), 
	.O4(O_int4), 
	.O5(O_int5), 
	.O6(O_int6), 
	.O7(O_int7), 
	.O8(O_int8)); 
	assign O = (  	O_int0 | 	O_int1 | 	O_int2 | 	O_int3 | 	O_int4 | 	O_int5 | 	O_int6 | 	O_int7 | 	O_int8 	); 

endmodule 

module precoder_32_18 (
	input logic  [4 : 0] S ,
	output logic  [31 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		5'd0    :   out_sel = 32'b00000000000000000000000000000001;
		5'd1    :   out_sel = 32'b00000000000000000000000000000010;
		5'd2    :   out_sel = 32'b00000000000000000000000000000100;
		5'd3    :   out_sel = 32'b00000000000000000000000000001000;
		5'd4    :   out_sel = 32'b00000000000000000000000000010000;
		5'd5    :   out_sel = 32'b00000000000000000000000000100000;
		5'd6    :   out_sel = 32'b00000000000000000000000001000000;
		5'd7    :   out_sel = 32'b00000000000000000000000010000000;
		5'd8    :   out_sel = 32'b00000000000000000000000100000000;
		5'd9    :   out_sel = 32'b00000000000000000000001000000000;
		5'd10    :   out_sel = 32'b00000000000000000000010000000000;
		5'd11    :   out_sel = 32'b00000000000000000000100000000000;
		5'd12    :   out_sel = 32'b00000000000000000001000000000000;
		5'd13    :   out_sel = 32'b00000000000000000010000000000000;
		5'd14    :   out_sel = 32'b00000000000000000100000000000000;
		5'd15    :   out_sel = 32'b00000000000000001000000000000000;
		5'd16    :   out_sel = 32'b00000000000000010000000000000000;
		5'd17    :   out_sel = 32'b00000000000000100000000000000000;
		default :   out_sel = 32'b0;
	endcase 
end 

endmodule 

module mux_logic_32_18 ( 
	input logic  [31 : 0] out_sel,
	input logic  [31 : 0] I0, 
	input logic  [31 : 0] I1, 
	input logic  [31 : 0] I2, 
	input logic  [31 : 0] I3, 
	input logic  [31 : 0] I4, 
	input logic  [31 : 0] I5, 
	input logic  [31 : 0] I6, 
	input logic  [31 : 0] I7, 
	input logic  [31 : 0] I8, 
	input logic  [31 : 0] I9, 
	input logic  [31 : 0] I10, 
	input logic  [31 : 0] I11, 
	input logic  [31 : 0] I12, 
	input logic  [31 : 0] I13, 
	input logic  [31 : 0] I14, 
	input logic  [31 : 0] I15, 
	input logic  [31 : 0] I16, 
	input logic  [31 : 0] I17, 
	output logic  [31 : 0] O0, 
	output logic  [31 : 0] O1, 
	output logic  [31 : 0] O2, 
	output logic  [31 : 0] O3, 
	output logic  [31 : 0] O4, 
	output logic  [31 : 0] O5, 
	output logic  [31 : 0] O6, 
	output logic  [31 : 0] O7, 
	output logic  [31 : 0] O8); 
	AO_CELL inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	AO_CELL inst_1_0 ( 
	.A1(out_sel[2]), 
	.A2(I2[0]), 
	.B1(out_sel[3]), 
	.B2(I3[0]), 
	.Z(O1[0])); 
	AO_CELL inst_2_0 ( 
	.A1(out_sel[4]), 
	.A2(I4[0]), 
	.B1(out_sel[5]), 
	.B2(I5[0]), 
	.Z(O2[0])); 
	AO_CELL inst_3_0 ( 
	.A1(out_sel[6]), 
	.A2(I6[0]), 
	.B1(out_sel[7]), 
	.B2(I7[0]), 
	.Z(O3[0])); 
	AO_CELL inst_4_0 ( 
	.A1(out_sel[8]), 
	.A2(I8[0]), 
	.B1(out_sel[9]), 
	.B2(I9[0]), 
	.Z(O4[0])); 
	AO_CELL inst_5_0 ( 
	.A1(out_sel[10]), 
	.A2(I10[0]), 
	.B1(out_sel[11]), 
	.B2(I11[0]), 
	.Z(O5[0])); 
	AO_CELL inst_6_0 ( 
	.A1(out_sel[12]), 
	.A2(I12[0]), 
	.B1(out_sel[13]), 
	.B2(I13[0]), 
	.Z(O6[0])); 
	AO_CELL inst_7_0 ( 
	.A1(out_sel[14]), 
	.A2(I14[0]), 
	.B1(out_sel[15]), 
	.B2(I15[0]), 
	.Z(O7[0])); 
	AO_CELL inst_8_0 ( 
	.A1(out_sel[16]), 
	.A2(I16[0]), 
	.B1(out_sel[17]), 
	.B2(I17[0]), 
	.Z(O8[0])); 
	AO_CELL inst_0_1 ( 
	.A1(out_sel[0]), 
	.A2(I0[1]), 
	.B1(out_sel[1]), 
	.B2(I1[1]), 
	.Z(O0[1])); 
	AO_CELL inst_1_1 ( 
	.A1(out_sel[2]), 
	.A2(I2[1]), 
	.B1(out_sel[3]), 
	.B2(I3[1]), 
	.Z(O1[1])); 
	AO_CELL inst_2_1 ( 
	.A1(out_sel[4]), 
	.A2(I4[1]), 
	.B1(out_sel[5]), 
	.B2(I5[1]), 
	.Z(O2[1])); 
	AO_CELL inst_3_1 ( 
	.A1(out_sel[6]), 
	.A2(I6[1]), 
	.B1(out_sel[7]), 
	.B2(I7[1]), 
	.Z(O3[1])); 
	AO_CELL inst_4_1 ( 
	.A1(out_sel[8]), 
	.A2(I8[1]), 
	.B1(out_sel[9]), 
	.B2(I9[1]), 
	.Z(O4[1])); 
	AO_CELL inst_5_1 ( 
	.A1(out_sel[10]), 
	.A2(I10[1]), 
	.B1(out_sel[11]), 
	.B2(I11[1]), 
	.Z(O5[1])); 
	AO_CELL inst_6_1 ( 
	.A1(out_sel[12]), 
	.A2(I12[1]), 
	.B1(out_sel[13]), 
	.B2(I13[1]), 
	.Z(O6[1])); 
	AO_CELL inst_7_1 ( 
	.A1(out_sel[14]), 
	.A2(I14[1]), 
	.B1(out_sel[15]), 
	.B2(I15[1]), 
	.Z(O7[1])); 
	AO_CELL inst_8_1 ( 
	.A1(out_sel[16]), 
	.A2(I16[1]), 
	.B1(out_sel[17]), 
	.B2(I17[1]), 
	.Z(O8[1])); 
	AO_CELL inst_0_2 ( 
	.A1(out_sel[0]), 
	.A2(I0[2]), 
	.B1(out_sel[1]), 
	.B2(I1[2]), 
	.Z(O0[2])); 
	AO_CELL inst_1_2 ( 
	.A1(out_sel[2]), 
	.A2(I2[2]), 
	.B1(out_sel[3]), 
	.B2(I3[2]), 
	.Z(O1[2])); 
	AO_CELL inst_2_2 ( 
	.A1(out_sel[4]), 
	.A2(I4[2]), 
	.B1(out_sel[5]), 
	.B2(I5[2]), 
	.Z(O2[2])); 
	AO_CELL inst_3_2 ( 
	.A1(out_sel[6]), 
	.A2(I6[2]), 
	.B1(out_sel[7]), 
	.B2(I7[2]), 
	.Z(O3[2])); 
	AO_CELL inst_4_2 ( 
	.A1(out_sel[8]), 
	.A2(I8[2]), 
	.B1(out_sel[9]), 
	.B2(I9[2]), 
	.Z(O4[2])); 
	AO_CELL inst_5_2 ( 
	.A1(out_sel[10]), 
	.A2(I10[2]), 
	.B1(out_sel[11]), 
	.B2(I11[2]), 
	.Z(O5[2])); 
	AO_CELL inst_6_2 ( 
	.A1(out_sel[12]), 
	.A2(I12[2]), 
	.B1(out_sel[13]), 
	.B2(I13[2]), 
	.Z(O6[2])); 
	AO_CELL inst_7_2 ( 
	.A1(out_sel[14]), 
	.A2(I14[2]), 
	.B1(out_sel[15]), 
	.B2(I15[2]), 
	.Z(O7[2])); 
	AO_CELL inst_8_2 ( 
	.A1(out_sel[16]), 
	.A2(I16[2]), 
	.B1(out_sel[17]), 
	.B2(I17[2]), 
	.Z(O8[2])); 
	AO_CELL inst_0_3 ( 
	.A1(out_sel[0]), 
	.A2(I0[3]), 
	.B1(out_sel[1]), 
	.B2(I1[3]), 
	.Z(O0[3])); 
	AO_CELL inst_1_3 ( 
	.A1(out_sel[2]), 
	.A2(I2[3]), 
	.B1(out_sel[3]), 
	.B2(I3[3]), 
	.Z(O1[3])); 
	AO_CELL inst_2_3 ( 
	.A1(out_sel[4]), 
	.A2(I4[3]), 
	.B1(out_sel[5]), 
	.B2(I5[3]), 
	.Z(O2[3])); 
	AO_CELL inst_3_3 ( 
	.A1(out_sel[6]), 
	.A2(I6[3]), 
	.B1(out_sel[7]), 
	.B2(I7[3]), 
	.Z(O3[3])); 
	AO_CELL inst_4_3 ( 
	.A1(out_sel[8]), 
	.A2(I8[3]), 
	.B1(out_sel[9]), 
	.B2(I9[3]), 
	.Z(O4[3])); 
	AO_CELL inst_5_3 ( 
	.A1(out_sel[10]), 
	.A2(I10[3]), 
	.B1(out_sel[11]), 
	.B2(I11[3]), 
	.Z(O5[3])); 
	AO_CELL inst_6_3 ( 
	.A1(out_sel[12]), 
	.A2(I12[3]), 
	.B1(out_sel[13]), 
	.B2(I13[3]), 
	.Z(O6[3])); 
	AO_CELL inst_7_3 ( 
	.A1(out_sel[14]), 
	.A2(I14[3]), 
	.B1(out_sel[15]), 
	.B2(I15[3]), 
	.Z(O7[3])); 
	AO_CELL inst_8_3 ( 
	.A1(out_sel[16]), 
	.A2(I16[3]), 
	.B1(out_sel[17]), 
	.B2(I17[3]), 
	.Z(O8[3])); 
	AO_CELL inst_0_4 ( 
	.A1(out_sel[0]), 
	.A2(I0[4]), 
	.B1(out_sel[1]), 
	.B2(I1[4]), 
	.Z(O0[4])); 
	AO_CELL inst_1_4 ( 
	.A1(out_sel[2]), 
	.A2(I2[4]), 
	.B1(out_sel[3]), 
	.B2(I3[4]), 
	.Z(O1[4])); 
	AO_CELL inst_2_4 ( 
	.A1(out_sel[4]), 
	.A2(I4[4]), 
	.B1(out_sel[5]), 
	.B2(I5[4]), 
	.Z(O2[4])); 
	AO_CELL inst_3_4 ( 
	.A1(out_sel[6]), 
	.A2(I6[4]), 
	.B1(out_sel[7]), 
	.B2(I7[4]), 
	.Z(O3[4])); 
	AO_CELL inst_4_4 ( 
	.A1(out_sel[8]), 
	.A2(I8[4]), 
	.B1(out_sel[9]), 
	.B2(I9[4]), 
	.Z(O4[4])); 
	AO_CELL inst_5_4 ( 
	.A1(out_sel[10]), 
	.A2(I10[4]), 
	.B1(out_sel[11]), 
	.B2(I11[4]), 
	.Z(O5[4])); 
	AO_CELL inst_6_4 ( 
	.A1(out_sel[12]), 
	.A2(I12[4]), 
	.B1(out_sel[13]), 
	.B2(I13[4]), 
	.Z(O6[4])); 
	AO_CELL inst_7_4 ( 
	.A1(out_sel[14]), 
	.A2(I14[4]), 
	.B1(out_sel[15]), 
	.B2(I15[4]), 
	.Z(O7[4])); 
	AO_CELL inst_8_4 ( 
	.A1(out_sel[16]), 
	.A2(I16[4]), 
	.B1(out_sel[17]), 
	.B2(I17[4]), 
	.Z(O8[4])); 
	AO_CELL inst_0_5 ( 
	.A1(out_sel[0]), 
	.A2(I0[5]), 
	.B1(out_sel[1]), 
	.B2(I1[5]), 
	.Z(O0[5])); 
	AO_CELL inst_1_5 ( 
	.A1(out_sel[2]), 
	.A2(I2[5]), 
	.B1(out_sel[3]), 
	.B2(I3[5]), 
	.Z(O1[5])); 
	AO_CELL inst_2_5 ( 
	.A1(out_sel[4]), 
	.A2(I4[5]), 
	.B1(out_sel[5]), 
	.B2(I5[5]), 
	.Z(O2[5])); 
	AO_CELL inst_3_5 ( 
	.A1(out_sel[6]), 
	.A2(I6[5]), 
	.B1(out_sel[7]), 
	.B2(I7[5]), 
	.Z(O3[5])); 
	AO_CELL inst_4_5 ( 
	.A1(out_sel[8]), 
	.A2(I8[5]), 
	.B1(out_sel[9]), 
	.B2(I9[5]), 
	.Z(O4[5])); 
	AO_CELL inst_5_5 ( 
	.A1(out_sel[10]), 
	.A2(I10[5]), 
	.B1(out_sel[11]), 
	.B2(I11[5]), 
	.Z(O5[5])); 
	AO_CELL inst_6_5 ( 
	.A1(out_sel[12]), 
	.A2(I12[5]), 
	.B1(out_sel[13]), 
	.B2(I13[5]), 
	.Z(O6[5])); 
	AO_CELL inst_7_5 ( 
	.A1(out_sel[14]), 
	.A2(I14[5]), 
	.B1(out_sel[15]), 
	.B2(I15[5]), 
	.Z(O7[5])); 
	AO_CELL inst_8_5 ( 
	.A1(out_sel[16]), 
	.A2(I16[5]), 
	.B1(out_sel[17]), 
	.B2(I17[5]), 
	.Z(O8[5])); 
	AO_CELL inst_0_6 ( 
	.A1(out_sel[0]), 
	.A2(I0[6]), 
	.B1(out_sel[1]), 
	.B2(I1[6]), 
	.Z(O0[6])); 
	AO_CELL inst_1_6 ( 
	.A1(out_sel[2]), 
	.A2(I2[6]), 
	.B1(out_sel[3]), 
	.B2(I3[6]), 
	.Z(O1[6])); 
	AO_CELL inst_2_6 ( 
	.A1(out_sel[4]), 
	.A2(I4[6]), 
	.B1(out_sel[5]), 
	.B2(I5[6]), 
	.Z(O2[6])); 
	AO_CELL inst_3_6 ( 
	.A1(out_sel[6]), 
	.A2(I6[6]), 
	.B1(out_sel[7]), 
	.B2(I7[6]), 
	.Z(O3[6])); 
	AO_CELL inst_4_6 ( 
	.A1(out_sel[8]), 
	.A2(I8[6]), 
	.B1(out_sel[9]), 
	.B2(I9[6]), 
	.Z(O4[6])); 
	AO_CELL inst_5_6 ( 
	.A1(out_sel[10]), 
	.A2(I10[6]), 
	.B1(out_sel[11]), 
	.B2(I11[6]), 
	.Z(O5[6])); 
	AO_CELL inst_6_6 ( 
	.A1(out_sel[12]), 
	.A2(I12[6]), 
	.B1(out_sel[13]), 
	.B2(I13[6]), 
	.Z(O6[6])); 
	AO_CELL inst_7_6 ( 
	.A1(out_sel[14]), 
	.A2(I14[6]), 
	.B1(out_sel[15]), 
	.B2(I15[6]), 
	.Z(O7[6])); 
	AO_CELL inst_8_6 ( 
	.A1(out_sel[16]), 
	.A2(I16[6]), 
	.B1(out_sel[17]), 
	.B2(I17[6]), 
	.Z(O8[6])); 
	AO_CELL inst_0_7 ( 
	.A1(out_sel[0]), 
	.A2(I0[7]), 
	.B1(out_sel[1]), 
	.B2(I1[7]), 
	.Z(O0[7])); 
	AO_CELL inst_1_7 ( 
	.A1(out_sel[2]), 
	.A2(I2[7]), 
	.B1(out_sel[3]), 
	.B2(I3[7]), 
	.Z(O1[7])); 
	AO_CELL inst_2_7 ( 
	.A1(out_sel[4]), 
	.A2(I4[7]), 
	.B1(out_sel[5]), 
	.B2(I5[7]), 
	.Z(O2[7])); 
	AO_CELL inst_3_7 ( 
	.A1(out_sel[6]), 
	.A2(I6[7]), 
	.B1(out_sel[7]), 
	.B2(I7[7]), 
	.Z(O3[7])); 
	AO_CELL inst_4_7 ( 
	.A1(out_sel[8]), 
	.A2(I8[7]), 
	.B1(out_sel[9]), 
	.B2(I9[7]), 
	.Z(O4[7])); 
	AO_CELL inst_5_7 ( 
	.A1(out_sel[10]), 
	.A2(I10[7]), 
	.B1(out_sel[11]), 
	.B2(I11[7]), 
	.Z(O5[7])); 
	AO_CELL inst_6_7 ( 
	.A1(out_sel[12]), 
	.A2(I12[7]), 
	.B1(out_sel[13]), 
	.B2(I13[7]), 
	.Z(O6[7])); 
	AO_CELL inst_7_7 ( 
	.A1(out_sel[14]), 
	.A2(I14[7]), 
	.B1(out_sel[15]), 
	.B2(I15[7]), 
	.Z(O7[7])); 
	AO_CELL inst_8_7 ( 
	.A1(out_sel[16]), 
	.A2(I16[7]), 
	.B1(out_sel[17]), 
	.B2(I17[7]), 
	.Z(O8[7])); 
	AO_CELL inst_0_8 ( 
	.A1(out_sel[0]), 
	.A2(I0[8]), 
	.B1(out_sel[1]), 
	.B2(I1[8]), 
	.Z(O0[8])); 
	AO_CELL inst_1_8 ( 
	.A1(out_sel[2]), 
	.A2(I2[8]), 
	.B1(out_sel[3]), 
	.B2(I3[8]), 
	.Z(O1[8])); 
	AO_CELL inst_2_8 ( 
	.A1(out_sel[4]), 
	.A2(I4[8]), 
	.B1(out_sel[5]), 
	.B2(I5[8]), 
	.Z(O2[8])); 
	AO_CELL inst_3_8 ( 
	.A1(out_sel[6]), 
	.A2(I6[8]), 
	.B1(out_sel[7]), 
	.B2(I7[8]), 
	.Z(O3[8])); 
	AO_CELL inst_4_8 ( 
	.A1(out_sel[8]), 
	.A2(I8[8]), 
	.B1(out_sel[9]), 
	.B2(I9[8]), 
	.Z(O4[8])); 
	AO_CELL inst_5_8 ( 
	.A1(out_sel[10]), 
	.A2(I10[8]), 
	.B1(out_sel[11]), 
	.B2(I11[8]), 
	.Z(O5[8])); 
	AO_CELL inst_6_8 ( 
	.A1(out_sel[12]), 
	.A2(I12[8]), 
	.B1(out_sel[13]), 
	.B2(I13[8]), 
	.Z(O6[8])); 
	AO_CELL inst_7_8 ( 
	.A1(out_sel[14]), 
	.A2(I14[8]), 
	.B1(out_sel[15]), 
	.B2(I15[8]), 
	.Z(O7[8])); 
	AO_CELL inst_8_8 ( 
	.A1(out_sel[16]), 
	.A2(I16[8]), 
	.B1(out_sel[17]), 
	.B2(I17[8]), 
	.Z(O8[8])); 
	AO_CELL inst_0_9 ( 
	.A1(out_sel[0]), 
	.A2(I0[9]), 
	.B1(out_sel[1]), 
	.B2(I1[9]), 
	.Z(O0[9])); 
	AO_CELL inst_1_9 ( 
	.A1(out_sel[2]), 
	.A2(I2[9]), 
	.B1(out_sel[3]), 
	.B2(I3[9]), 
	.Z(O1[9])); 
	AO_CELL inst_2_9 ( 
	.A1(out_sel[4]), 
	.A2(I4[9]), 
	.B1(out_sel[5]), 
	.B2(I5[9]), 
	.Z(O2[9])); 
	AO_CELL inst_3_9 ( 
	.A1(out_sel[6]), 
	.A2(I6[9]), 
	.B1(out_sel[7]), 
	.B2(I7[9]), 
	.Z(O3[9])); 
	AO_CELL inst_4_9 ( 
	.A1(out_sel[8]), 
	.A2(I8[9]), 
	.B1(out_sel[9]), 
	.B2(I9[9]), 
	.Z(O4[9])); 
	AO_CELL inst_5_9 ( 
	.A1(out_sel[10]), 
	.A2(I10[9]), 
	.B1(out_sel[11]), 
	.B2(I11[9]), 
	.Z(O5[9])); 
	AO_CELL inst_6_9 ( 
	.A1(out_sel[12]), 
	.A2(I12[9]), 
	.B1(out_sel[13]), 
	.B2(I13[9]), 
	.Z(O6[9])); 
	AO_CELL inst_7_9 ( 
	.A1(out_sel[14]), 
	.A2(I14[9]), 
	.B1(out_sel[15]), 
	.B2(I15[9]), 
	.Z(O7[9])); 
	AO_CELL inst_8_9 ( 
	.A1(out_sel[16]), 
	.A2(I16[9]), 
	.B1(out_sel[17]), 
	.B2(I17[9]), 
	.Z(O8[9])); 
	AO_CELL inst_0_10 ( 
	.A1(out_sel[0]), 
	.A2(I0[10]), 
	.B1(out_sel[1]), 
	.B2(I1[10]), 
	.Z(O0[10])); 
	AO_CELL inst_1_10 ( 
	.A1(out_sel[2]), 
	.A2(I2[10]), 
	.B1(out_sel[3]), 
	.B2(I3[10]), 
	.Z(O1[10])); 
	AO_CELL inst_2_10 ( 
	.A1(out_sel[4]), 
	.A2(I4[10]), 
	.B1(out_sel[5]), 
	.B2(I5[10]), 
	.Z(O2[10])); 
	AO_CELL inst_3_10 ( 
	.A1(out_sel[6]), 
	.A2(I6[10]), 
	.B1(out_sel[7]), 
	.B2(I7[10]), 
	.Z(O3[10])); 
	AO_CELL inst_4_10 ( 
	.A1(out_sel[8]), 
	.A2(I8[10]), 
	.B1(out_sel[9]), 
	.B2(I9[10]), 
	.Z(O4[10])); 
	AO_CELL inst_5_10 ( 
	.A1(out_sel[10]), 
	.A2(I10[10]), 
	.B1(out_sel[11]), 
	.B2(I11[10]), 
	.Z(O5[10])); 
	AO_CELL inst_6_10 ( 
	.A1(out_sel[12]), 
	.A2(I12[10]), 
	.B1(out_sel[13]), 
	.B2(I13[10]), 
	.Z(O6[10])); 
	AO_CELL inst_7_10 ( 
	.A1(out_sel[14]), 
	.A2(I14[10]), 
	.B1(out_sel[15]), 
	.B2(I15[10]), 
	.Z(O7[10])); 
	AO_CELL inst_8_10 ( 
	.A1(out_sel[16]), 
	.A2(I16[10]), 
	.B1(out_sel[17]), 
	.B2(I17[10]), 
	.Z(O8[10])); 
	AO_CELL inst_0_11 ( 
	.A1(out_sel[0]), 
	.A2(I0[11]), 
	.B1(out_sel[1]), 
	.B2(I1[11]), 
	.Z(O0[11])); 
	AO_CELL inst_1_11 ( 
	.A1(out_sel[2]), 
	.A2(I2[11]), 
	.B1(out_sel[3]), 
	.B2(I3[11]), 
	.Z(O1[11])); 
	AO_CELL inst_2_11 ( 
	.A1(out_sel[4]), 
	.A2(I4[11]), 
	.B1(out_sel[5]), 
	.B2(I5[11]), 
	.Z(O2[11])); 
	AO_CELL inst_3_11 ( 
	.A1(out_sel[6]), 
	.A2(I6[11]), 
	.B1(out_sel[7]), 
	.B2(I7[11]), 
	.Z(O3[11])); 
	AO_CELL inst_4_11 ( 
	.A1(out_sel[8]), 
	.A2(I8[11]), 
	.B1(out_sel[9]), 
	.B2(I9[11]), 
	.Z(O4[11])); 
	AO_CELL inst_5_11 ( 
	.A1(out_sel[10]), 
	.A2(I10[11]), 
	.B1(out_sel[11]), 
	.B2(I11[11]), 
	.Z(O5[11])); 
	AO_CELL inst_6_11 ( 
	.A1(out_sel[12]), 
	.A2(I12[11]), 
	.B1(out_sel[13]), 
	.B2(I13[11]), 
	.Z(O6[11])); 
	AO_CELL inst_7_11 ( 
	.A1(out_sel[14]), 
	.A2(I14[11]), 
	.B1(out_sel[15]), 
	.B2(I15[11]), 
	.Z(O7[11])); 
	AO_CELL inst_8_11 ( 
	.A1(out_sel[16]), 
	.A2(I16[11]), 
	.B1(out_sel[17]), 
	.B2(I17[11]), 
	.Z(O8[11])); 
	AO_CELL inst_0_12 ( 
	.A1(out_sel[0]), 
	.A2(I0[12]), 
	.B1(out_sel[1]), 
	.B2(I1[12]), 
	.Z(O0[12])); 
	AO_CELL inst_1_12 ( 
	.A1(out_sel[2]), 
	.A2(I2[12]), 
	.B1(out_sel[3]), 
	.B2(I3[12]), 
	.Z(O1[12])); 
	AO_CELL inst_2_12 ( 
	.A1(out_sel[4]), 
	.A2(I4[12]), 
	.B1(out_sel[5]), 
	.B2(I5[12]), 
	.Z(O2[12])); 
	AO_CELL inst_3_12 ( 
	.A1(out_sel[6]), 
	.A2(I6[12]), 
	.B1(out_sel[7]), 
	.B2(I7[12]), 
	.Z(O3[12])); 
	AO_CELL inst_4_12 ( 
	.A1(out_sel[8]), 
	.A2(I8[12]), 
	.B1(out_sel[9]), 
	.B2(I9[12]), 
	.Z(O4[12])); 
	AO_CELL inst_5_12 ( 
	.A1(out_sel[10]), 
	.A2(I10[12]), 
	.B1(out_sel[11]), 
	.B2(I11[12]), 
	.Z(O5[12])); 
	AO_CELL inst_6_12 ( 
	.A1(out_sel[12]), 
	.A2(I12[12]), 
	.B1(out_sel[13]), 
	.B2(I13[12]), 
	.Z(O6[12])); 
	AO_CELL inst_7_12 ( 
	.A1(out_sel[14]), 
	.A2(I14[12]), 
	.B1(out_sel[15]), 
	.B2(I15[12]), 
	.Z(O7[12])); 
	AO_CELL inst_8_12 ( 
	.A1(out_sel[16]), 
	.A2(I16[12]), 
	.B1(out_sel[17]), 
	.B2(I17[12]), 
	.Z(O8[12])); 
	AO_CELL inst_0_13 ( 
	.A1(out_sel[0]), 
	.A2(I0[13]), 
	.B1(out_sel[1]), 
	.B2(I1[13]), 
	.Z(O0[13])); 
	AO_CELL inst_1_13 ( 
	.A1(out_sel[2]), 
	.A2(I2[13]), 
	.B1(out_sel[3]), 
	.B2(I3[13]), 
	.Z(O1[13])); 
	AO_CELL inst_2_13 ( 
	.A1(out_sel[4]), 
	.A2(I4[13]), 
	.B1(out_sel[5]), 
	.B2(I5[13]), 
	.Z(O2[13])); 
	AO_CELL inst_3_13 ( 
	.A1(out_sel[6]), 
	.A2(I6[13]), 
	.B1(out_sel[7]), 
	.B2(I7[13]), 
	.Z(O3[13])); 
	AO_CELL inst_4_13 ( 
	.A1(out_sel[8]), 
	.A2(I8[13]), 
	.B1(out_sel[9]), 
	.B2(I9[13]), 
	.Z(O4[13])); 
	AO_CELL inst_5_13 ( 
	.A1(out_sel[10]), 
	.A2(I10[13]), 
	.B1(out_sel[11]), 
	.B2(I11[13]), 
	.Z(O5[13])); 
	AO_CELL inst_6_13 ( 
	.A1(out_sel[12]), 
	.A2(I12[13]), 
	.B1(out_sel[13]), 
	.B2(I13[13]), 
	.Z(O6[13])); 
	AO_CELL inst_7_13 ( 
	.A1(out_sel[14]), 
	.A2(I14[13]), 
	.B1(out_sel[15]), 
	.B2(I15[13]), 
	.Z(O7[13])); 
	AO_CELL inst_8_13 ( 
	.A1(out_sel[16]), 
	.A2(I16[13]), 
	.B1(out_sel[17]), 
	.B2(I17[13]), 
	.Z(O8[13])); 
	AO_CELL inst_0_14 ( 
	.A1(out_sel[0]), 
	.A2(I0[14]), 
	.B1(out_sel[1]), 
	.B2(I1[14]), 
	.Z(O0[14])); 
	AO_CELL inst_1_14 ( 
	.A1(out_sel[2]), 
	.A2(I2[14]), 
	.B1(out_sel[3]), 
	.B2(I3[14]), 
	.Z(O1[14])); 
	AO_CELL inst_2_14 ( 
	.A1(out_sel[4]), 
	.A2(I4[14]), 
	.B1(out_sel[5]), 
	.B2(I5[14]), 
	.Z(O2[14])); 
	AO_CELL inst_3_14 ( 
	.A1(out_sel[6]), 
	.A2(I6[14]), 
	.B1(out_sel[7]), 
	.B2(I7[14]), 
	.Z(O3[14])); 
	AO_CELL inst_4_14 ( 
	.A1(out_sel[8]), 
	.A2(I8[14]), 
	.B1(out_sel[9]), 
	.B2(I9[14]), 
	.Z(O4[14])); 
	AO_CELL inst_5_14 ( 
	.A1(out_sel[10]), 
	.A2(I10[14]), 
	.B1(out_sel[11]), 
	.B2(I11[14]), 
	.Z(O5[14])); 
	AO_CELL inst_6_14 ( 
	.A1(out_sel[12]), 
	.A2(I12[14]), 
	.B1(out_sel[13]), 
	.B2(I13[14]), 
	.Z(O6[14])); 
	AO_CELL inst_7_14 ( 
	.A1(out_sel[14]), 
	.A2(I14[14]), 
	.B1(out_sel[15]), 
	.B2(I15[14]), 
	.Z(O7[14])); 
	AO_CELL inst_8_14 ( 
	.A1(out_sel[16]), 
	.A2(I16[14]), 
	.B1(out_sel[17]), 
	.B2(I17[14]), 
	.Z(O8[14])); 
	AO_CELL inst_0_15 ( 
	.A1(out_sel[0]), 
	.A2(I0[15]), 
	.B1(out_sel[1]), 
	.B2(I1[15]), 
	.Z(O0[15])); 
	AO_CELL inst_1_15 ( 
	.A1(out_sel[2]), 
	.A2(I2[15]), 
	.B1(out_sel[3]), 
	.B2(I3[15]), 
	.Z(O1[15])); 
	AO_CELL inst_2_15 ( 
	.A1(out_sel[4]), 
	.A2(I4[15]), 
	.B1(out_sel[5]), 
	.B2(I5[15]), 
	.Z(O2[15])); 
	AO_CELL inst_3_15 ( 
	.A1(out_sel[6]), 
	.A2(I6[15]), 
	.B1(out_sel[7]), 
	.B2(I7[15]), 
	.Z(O3[15])); 
	AO_CELL inst_4_15 ( 
	.A1(out_sel[8]), 
	.A2(I8[15]), 
	.B1(out_sel[9]), 
	.B2(I9[15]), 
	.Z(O4[15])); 
	AO_CELL inst_5_15 ( 
	.A1(out_sel[10]), 
	.A2(I10[15]), 
	.B1(out_sel[11]), 
	.B2(I11[15]), 
	.Z(O5[15])); 
	AO_CELL inst_6_15 ( 
	.A1(out_sel[12]), 
	.A2(I12[15]), 
	.B1(out_sel[13]), 
	.B2(I13[15]), 
	.Z(O6[15])); 
	AO_CELL inst_7_15 ( 
	.A1(out_sel[14]), 
	.A2(I14[15]), 
	.B1(out_sel[15]), 
	.B2(I15[15]), 
	.Z(O7[15])); 
	AO_CELL inst_8_15 ( 
	.A1(out_sel[16]), 
	.A2(I16[15]), 
	.B1(out_sel[17]), 
	.B2(I17[15]), 
	.Z(O8[15])); 
	AO_CELL inst_0_16 ( 
	.A1(out_sel[0]), 
	.A2(I0[16]), 
	.B1(out_sel[1]), 
	.B2(I1[16]), 
	.Z(O0[16])); 
	AO_CELL inst_1_16 ( 
	.A1(out_sel[2]), 
	.A2(I2[16]), 
	.B1(out_sel[3]), 
	.B2(I3[16]), 
	.Z(O1[16])); 
	AO_CELL inst_2_16 ( 
	.A1(out_sel[4]), 
	.A2(I4[16]), 
	.B1(out_sel[5]), 
	.B2(I5[16]), 
	.Z(O2[16])); 
	AO_CELL inst_3_16 ( 
	.A1(out_sel[6]), 
	.A2(I6[16]), 
	.B1(out_sel[7]), 
	.B2(I7[16]), 
	.Z(O3[16])); 
	AO_CELL inst_4_16 ( 
	.A1(out_sel[8]), 
	.A2(I8[16]), 
	.B1(out_sel[9]), 
	.B2(I9[16]), 
	.Z(O4[16])); 
	AO_CELL inst_5_16 ( 
	.A1(out_sel[10]), 
	.A2(I10[16]), 
	.B1(out_sel[11]), 
	.B2(I11[16]), 
	.Z(O5[16])); 
	AO_CELL inst_6_16 ( 
	.A1(out_sel[12]), 
	.A2(I12[16]), 
	.B1(out_sel[13]), 
	.B2(I13[16]), 
	.Z(O6[16])); 
	AO_CELL inst_7_16 ( 
	.A1(out_sel[14]), 
	.A2(I14[16]), 
	.B1(out_sel[15]), 
	.B2(I15[16]), 
	.Z(O7[16])); 
	AO_CELL inst_8_16 ( 
	.A1(out_sel[16]), 
	.A2(I16[16]), 
	.B1(out_sel[17]), 
	.B2(I17[16]), 
	.Z(O8[16])); 
	AO_CELL inst_0_17 ( 
	.A1(out_sel[0]), 
	.A2(I0[17]), 
	.B1(out_sel[1]), 
	.B2(I1[17]), 
	.Z(O0[17])); 
	AO_CELL inst_1_17 ( 
	.A1(out_sel[2]), 
	.A2(I2[17]), 
	.B1(out_sel[3]), 
	.B2(I3[17]), 
	.Z(O1[17])); 
	AO_CELL inst_2_17 ( 
	.A1(out_sel[4]), 
	.A2(I4[17]), 
	.B1(out_sel[5]), 
	.B2(I5[17]), 
	.Z(O2[17])); 
	AO_CELL inst_3_17 ( 
	.A1(out_sel[6]), 
	.A2(I6[17]), 
	.B1(out_sel[7]), 
	.B2(I7[17]), 
	.Z(O3[17])); 
	AO_CELL inst_4_17 ( 
	.A1(out_sel[8]), 
	.A2(I8[17]), 
	.B1(out_sel[9]), 
	.B2(I9[17]), 
	.Z(O4[17])); 
	AO_CELL inst_5_17 ( 
	.A1(out_sel[10]), 
	.A2(I10[17]), 
	.B1(out_sel[11]), 
	.B2(I11[17]), 
	.Z(O5[17])); 
	AO_CELL inst_6_17 ( 
	.A1(out_sel[12]), 
	.A2(I12[17]), 
	.B1(out_sel[13]), 
	.B2(I13[17]), 
	.Z(O6[17])); 
	AO_CELL inst_7_17 ( 
	.A1(out_sel[14]), 
	.A2(I14[17]), 
	.B1(out_sel[15]), 
	.B2(I15[17]), 
	.Z(O7[17])); 
	AO_CELL inst_8_17 ( 
	.A1(out_sel[16]), 
	.A2(I16[17]), 
	.B1(out_sel[17]), 
	.B2(I17[17]), 
	.Z(O8[17])); 
	AO_CELL inst_0_18 ( 
	.A1(out_sel[0]), 
	.A2(I0[18]), 
	.B1(out_sel[1]), 
	.B2(I1[18]), 
	.Z(O0[18])); 
	AO_CELL inst_1_18 ( 
	.A1(out_sel[2]), 
	.A2(I2[18]), 
	.B1(out_sel[3]), 
	.B2(I3[18]), 
	.Z(O1[18])); 
	AO_CELL inst_2_18 ( 
	.A1(out_sel[4]), 
	.A2(I4[18]), 
	.B1(out_sel[5]), 
	.B2(I5[18]), 
	.Z(O2[18])); 
	AO_CELL inst_3_18 ( 
	.A1(out_sel[6]), 
	.A2(I6[18]), 
	.B1(out_sel[7]), 
	.B2(I7[18]), 
	.Z(O3[18])); 
	AO_CELL inst_4_18 ( 
	.A1(out_sel[8]), 
	.A2(I8[18]), 
	.B1(out_sel[9]), 
	.B2(I9[18]), 
	.Z(O4[18])); 
	AO_CELL inst_5_18 ( 
	.A1(out_sel[10]), 
	.A2(I10[18]), 
	.B1(out_sel[11]), 
	.B2(I11[18]), 
	.Z(O5[18])); 
	AO_CELL inst_6_18 ( 
	.A1(out_sel[12]), 
	.A2(I12[18]), 
	.B1(out_sel[13]), 
	.B2(I13[18]), 
	.Z(O6[18])); 
	AO_CELL inst_7_18 ( 
	.A1(out_sel[14]), 
	.A2(I14[18]), 
	.B1(out_sel[15]), 
	.B2(I15[18]), 
	.Z(O7[18])); 
	AO_CELL inst_8_18 ( 
	.A1(out_sel[16]), 
	.A2(I16[18]), 
	.B1(out_sel[17]), 
	.B2(I17[18]), 
	.Z(O8[18])); 
	AO_CELL inst_0_19 ( 
	.A1(out_sel[0]), 
	.A2(I0[19]), 
	.B1(out_sel[1]), 
	.B2(I1[19]), 
	.Z(O0[19])); 
	AO_CELL inst_1_19 ( 
	.A1(out_sel[2]), 
	.A2(I2[19]), 
	.B1(out_sel[3]), 
	.B2(I3[19]), 
	.Z(O1[19])); 
	AO_CELL inst_2_19 ( 
	.A1(out_sel[4]), 
	.A2(I4[19]), 
	.B1(out_sel[5]), 
	.B2(I5[19]), 
	.Z(O2[19])); 
	AO_CELL inst_3_19 ( 
	.A1(out_sel[6]), 
	.A2(I6[19]), 
	.B1(out_sel[7]), 
	.B2(I7[19]), 
	.Z(O3[19])); 
	AO_CELL inst_4_19 ( 
	.A1(out_sel[8]), 
	.A2(I8[19]), 
	.B1(out_sel[9]), 
	.B2(I9[19]), 
	.Z(O4[19])); 
	AO_CELL inst_5_19 ( 
	.A1(out_sel[10]), 
	.A2(I10[19]), 
	.B1(out_sel[11]), 
	.B2(I11[19]), 
	.Z(O5[19])); 
	AO_CELL inst_6_19 ( 
	.A1(out_sel[12]), 
	.A2(I12[19]), 
	.B1(out_sel[13]), 
	.B2(I13[19]), 
	.Z(O6[19])); 
	AO_CELL inst_7_19 ( 
	.A1(out_sel[14]), 
	.A2(I14[19]), 
	.B1(out_sel[15]), 
	.B2(I15[19]), 
	.Z(O7[19])); 
	AO_CELL inst_8_19 ( 
	.A1(out_sel[16]), 
	.A2(I16[19]), 
	.B1(out_sel[17]), 
	.B2(I17[19]), 
	.Z(O8[19])); 
	AO_CELL inst_0_20 ( 
	.A1(out_sel[0]), 
	.A2(I0[20]), 
	.B1(out_sel[1]), 
	.B2(I1[20]), 
	.Z(O0[20])); 
	AO_CELL inst_1_20 ( 
	.A1(out_sel[2]), 
	.A2(I2[20]), 
	.B1(out_sel[3]), 
	.B2(I3[20]), 
	.Z(O1[20])); 
	AO_CELL inst_2_20 ( 
	.A1(out_sel[4]), 
	.A2(I4[20]), 
	.B1(out_sel[5]), 
	.B2(I5[20]), 
	.Z(O2[20])); 
	AO_CELL inst_3_20 ( 
	.A1(out_sel[6]), 
	.A2(I6[20]), 
	.B1(out_sel[7]), 
	.B2(I7[20]), 
	.Z(O3[20])); 
	AO_CELL inst_4_20 ( 
	.A1(out_sel[8]), 
	.A2(I8[20]), 
	.B1(out_sel[9]), 
	.B2(I9[20]), 
	.Z(O4[20])); 
	AO_CELL inst_5_20 ( 
	.A1(out_sel[10]), 
	.A2(I10[20]), 
	.B1(out_sel[11]), 
	.B2(I11[20]), 
	.Z(O5[20])); 
	AO_CELL inst_6_20 ( 
	.A1(out_sel[12]), 
	.A2(I12[20]), 
	.B1(out_sel[13]), 
	.B2(I13[20]), 
	.Z(O6[20])); 
	AO_CELL inst_7_20 ( 
	.A1(out_sel[14]), 
	.A2(I14[20]), 
	.B1(out_sel[15]), 
	.B2(I15[20]), 
	.Z(O7[20])); 
	AO_CELL inst_8_20 ( 
	.A1(out_sel[16]), 
	.A2(I16[20]), 
	.B1(out_sel[17]), 
	.B2(I17[20]), 
	.Z(O8[20])); 
	AO_CELL inst_0_21 ( 
	.A1(out_sel[0]), 
	.A2(I0[21]), 
	.B1(out_sel[1]), 
	.B2(I1[21]), 
	.Z(O0[21])); 
	AO_CELL inst_1_21 ( 
	.A1(out_sel[2]), 
	.A2(I2[21]), 
	.B1(out_sel[3]), 
	.B2(I3[21]), 
	.Z(O1[21])); 
	AO_CELL inst_2_21 ( 
	.A1(out_sel[4]), 
	.A2(I4[21]), 
	.B1(out_sel[5]), 
	.B2(I5[21]), 
	.Z(O2[21])); 
	AO_CELL inst_3_21 ( 
	.A1(out_sel[6]), 
	.A2(I6[21]), 
	.B1(out_sel[7]), 
	.B2(I7[21]), 
	.Z(O3[21])); 
	AO_CELL inst_4_21 ( 
	.A1(out_sel[8]), 
	.A2(I8[21]), 
	.B1(out_sel[9]), 
	.B2(I9[21]), 
	.Z(O4[21])); 
	AO_CELL inst_5_21 ( 
	.A1(out_sel[10]), 
	.A2(I10[21]), 
	.B1(out_sel[11]), 
	.B2(I11[21]), 
	.Z(O5[21])); 
	AO_CELL inst_6_21 ( 
	.A1(out_sel[12]), 
	.A2(I12[21]), 
	.B1(out_sel[13]), 
	.B2(I13[21]), 
	.Z(O6[21])); 
	AO_CELL inst_7_21 ( 
	.A1(out_sel[14]), 
	.A2(I14[21]), 
	.B1(out_sel[15]), 
	.B2(I15[21]), 
	.Z(O7[21])); 
	AO_CELL inst_8_21 ( 
	.A1(out_sel[16]), 
	.A2(I16[21]), 
	.B1(out_sel[17]), 
	.B2(I17[21]), 
	.Z(O8[21])); 
	AO_CELL inst_0_22 ( 
	.A1(out_sel[0]), 
	.A2(I0[22]), 
	.B1(out_sel[1]), 
	.B2(I1[22]), 
	.Z(O0[22])); 
	AO_CELL inst_1_22 ( 
	.A1(out_sel[2]), 
	.A2(I2[22]), 
	.B1(out_sel[3]), 
	.B2(I3[22]), 
	.Z(O1[22])); 
	AO_CELL inst_2_22 ( 
	.A1(out_sel[4]), 
	.A2(I4[22]), 
	.B1(out_sel[5]), 
	.B2(I5[22]), 
	.Z(O2[22])); 
	AO_CELL inst_3_22 ( 
	.A1(out_sel[6]), 
	.A2(I6[22]), 
	.B1(out_sel[7]), 
	.B2(I7[22]), 
	.Z(O3[22])); 
	AO_CELL inst_4_22 ( 
	.A1(out_sel[8]), 
	.A2(I8[22]), 
	.B1(out_sel[9]), 
	.B2(I9[22]), 
	.Z(O4[22])); 
	AO_CELL inst_5_22 ( 
	.A1(out_sel[10]), 
	.A2(I10[22]), 
	.B1(out_sel[11]), 
	.B2(I11[22]), 
	.Z(O5[22])); 
	AO_CELL inst_6_22 ( 
	.A1(out_sel[12]), 
	.A2(I12[22]), 
	.B1(out_sel[13]), 
	.B2(I13[22]), 
	.Z(O6[22])); 
	AO_CELL inst_7_22 ( 
	.A1(out_sel[14]), 
	.A2(I14[22]), 
	.B1(out_sel[15]), 
	.B2(I15[22]), 
	.Z(O7[22])); 
	AO_CELL inst_8_22 ( 
	.A1(out_sel[16]), 
	.A2(I16[22]), 
	.B1(out_sel[17]), 
	.B2(I17[22]), 
	.Z(O8[22])); 
	AO_CELL inst_0_23 ( 
	.A1(out_sel[0]), 
	.A2(I0[23]), 
	.B1(out_sel[1]), 
	.B2(I1[23]), 
	.Z(O0[23])); 
	AO_CELL inst_1_23 ( 
	.A1(out_sel[2]), 
	.A2(I2[23]), 
	.B1(out_sel[3]), 
	.B2(I3[23]), 
	.Z(O1[23])); 
	AO_CELL inst_2_23 ( 
	.A1(out_sel[4]), 
	.A2(I4[23]), 
	.B1(out_sel[5]), 
	.B2(I5[23]), 
	.Z(O2[23])); 
	AO_CELL inst_3_23 ( 
	.A1(out_sel[6]), 
	.A2(I6[23]), 
	.B1(out_sel[7]), 
	.B2(I7[23]), 
	.Z(O3[23])); 
	AO_CELL inst_4_23 ( 
	.A1(out_sel[8]), 
	.A2(I8[23]), 
	.B1(out_sel[9]), 
	.B2(I9[23]), 
	.Z(O4[23])); 
	AO_CELL inst_5_23 ( 
	.A1(out_sel[10]), 
	.A2(I10[23]), 
	.B1(out_sel[11]), 
	.B2(I11[23]), 
	.Z(O5[23])); 
	AO_CELL inst_6_23 ( 
	.A1(out_sel[12]), 
	.A2(I12[23]), 
	.B1(out_sel[13]), 
	.B2(I13[23]), 
	.Z(O6[23])); 
	AO_CELL inst_7_23 ( 
	.A1(out_sel[14]), 
	.A2(I14[23]), 
	.B1(out_sel[15]), 
	.B2(I15[23]), 
	.Z(O7[23])); 
	AO_CELL inst_8_23 ( 
	.A1(out_sel[16]), 
	.A2(I16[23]), 
	.B1(out_sel[17]), 
	.B2(I17[23]), 
	.Z(O8[23])); 
	AO_CELL inst_0_24 ( 
	.A1(out_sel[0]), 
	.A2(I0[24]), 
	.B1(out_sel[1]), 
	.B2(I1[24]), 
	.Z(O0[24])); 
	AO_CELL inst_1_24 ( 
	.A1(out_sel[2]), 
	.A2(I2[24]), 
	.B1(out_sel[3]), 
	.B2(I3[24]), 
	.Z(O1[24])); 
	AO_CELL inst_2_24 ( 
	.A1(out_sel[4]), 
	.A2(I4[24]), 
	.B1(out_sel[5]), 
	.B2(I5[24]), 
	.Z(O2[24])); 
	AO_CELL inst_3_24 ( 
	.A1(out_sel[6]), 
	.A2(I6[24]), 
	.B1(out_sel[7]), 
	.B2(I7[24]), 
	.Z(O3[24])); 
	AO_CELL inst_4_24 ( 
	.A1(out_sel[8]), 
	.A2(I8[24]), 
	.B1(out_sel[9]), 
	.B2(I9[24]), 
	.Z(O4[24])); 
	AO_CELL inst_5_24 ( 
	.A1(out_sel[10]), 
	.A2(I10[24]), 
	.B1(out_sel[11]), 
	.B2(I11[24]), 
	.Z(O5[24])); 
	AO_CELL inst_6_24 ( 
	.A1(out_sel[12]), 
	.A2(I12[24]), 
	.B1(out_sel[13]), 
	.B2(I13[24]), 
	.Z(O6[24])); 
	AO_CELL inst_7_24 ( 
	.A1(out_sel[14]), 
	.A2(I14[24]), 
	.B1(out_sel[15]), 
	.B2(I15[24]), 
	.Z(O7[24])); 
	AO_CELL inst_8_24 ( 
	.A1(out_sel[16]), 
	.A2(I16[24]), 
	.B1(out_sel[17]), 
	.B2(I17[24]), 
	.Z(O8[24])); 
	AO_CELL inst_0_25 ( 
	.A1(out_sel[0]), 
	.A2(I0[25]), 
	.B1(out_sel[1]), 
	.B2(I1[25]), 
	.Z(O0[25])); 
	AO_CELL inst_1_25 ( 
	.A1(out_sel[2]), 
	.A2(I2[25]), 
	.B1(out_sel[3]), 
	.B2(I3[25]), 
	.Z(O1[25])); 
	AO_CELL inst_2_25 ( 
	.A1(out_sel[4]), 
	.A2(I4[25]), 
	.B1(out_sel[5]), 
	.B2(I5[25]), 
	.Z(O2[25])); 
	AO_CELL inst_3_25 ( 
	.A1(out_sel[6]), 
	.A2(I6[25]), 
	.B1(out_sel[7]), 
	.B2(I7[25]), 
	.Z(O3[25])); 
	AO_CELL inst_4_25 ( 
	.A1(out_sel[8]), 
	.A2(I8[25]), 
	.B1(out_sel[9]), 
	.B2(I9[25]), 
	.Z(O4[25])); 
	AO_CELL inst_5_25 ( 
	.A1(out_sel[10]), 
	.A2(I10[25]), 
	.B1(out_sel[11]), 
	.B2(I11[25]), 
	.Z(O5[25])); 
	AO_CELL inst_6_25 ( 
	.A1(out_sel[12]), 
	.A2(I12[25]), 
	.B1(out_sel[13]), 
	.B2(I13[25]), 
	.Z(O6[25])); 
	AO_CELL inst_7_25 ( 
	.A1(out_sel[14]), 
	.A2(I14[25]), 
	.B1(out_sel[15]), 
	.B2(I15[25]), 
	.Z(O7[25])); 
	AO_CELL inst_8_25 ( 
	.A1(out_sel[16]), 
	.A2(I16[25]), 
	.B1(out_sel[17]), 
	.B2(I17[25]), 
	.Z(O8[25])); 
	AO_CELL inst_0_26 ( 
	.A1(out_sel[0]), 
	.A2(I0[26]), 
	.B1(out_sel[1]), 
	.B2(I1[26]), 
	.Z(O0[26])); 
	AO_CELL inst_1_26 ( 
	.A1(out_sel[2]), 
	.A2(I2[26]), 
	.B1(out_sel[3]), 
	.B2(I3[26]), 
	.Z(O1[26])); 
	AO_CELL inst_2_26 ( 
	.A1(out_sel[4]), 
	.A2(I4[26]), 
	.B1(out_sel[5]), 
	.B2(I5[26]), 
	.Z(O2[26])); 
	AO_CELL inst_3_26 ( 
	.A1(out_sel[6]), 
	.A2(I6[26]), 
	.B1(out_sel[7]), 
	.B2(I7[26]), 
	.Z(O3[26])); 
	AO_CELL inst_4_26 ( 
	.A1(out_sel[8]), 
	.A2(I8[26]), 
	.B1(out_sel[9]), 
	.B2(I9[26]), 
	.Z(O4[26])); 
	AO_CELL inst_5_26 ( 
	.A1(out_sel[10]), 
	.A2(I10[26]), 
	.B1(out_sel[11]), 
	.B2(I11[26]), 
	.Z(O5[26])); 
	AO_CELL inst_6_26 ( 
	.A1(out_sel[12]), 
	.A2(I12[26]), 
	.B1(out_sel[13]), 
	.B2(I13[26]), 
	.Z(O6[26])); 
	AO_CELL inst_7_26 ( 
	.A1(out_sel[14]), 
	.A2(I14[26]), 
	.B1(out_sel[15]), 
	.B2(I15[26]), 
	.Z(O7[26])); 
	AO_CELL inst_8_26 ( 
	.A1(out_sel[16]), 
	.A2(I16[26]), 
	.B1(out_sel[17]), 
	.B2(I17[26]), 
	.Z(O8[26])); 
	AO_CELL inst_0_27 ( 
	.A1(out_sel[0]), 
	.A2(I0[27]), 
	.B1(out_sel[1]), 
	.B2(I1[27]), 
	.Z(O0[27])); 
	AO_CELL inst_1_27 ( 
	.A1(out_sel[2]), 
	.A2(I2[27]), 
	.B1(out_sel[3]), 
	.B2(I3[27]), 
	.Z(O1[27])); 
	AO_CELL inst_2_27 ( 
	.A1(out_sel[4]), 
	.A2(I4[27]), 
	.B1(out_sel[5]), 
	.B2(I5[27]), 
	.Z(O2[27])); 
	AO_CELL inst_3_27 ( 
	.A1(out_sel[6]), 
	.A2(I6[27]), 
	.B1(out_sel[7]), 
	.B2(I7[27]), 
	.Z(O3[27])); 
	AO_CELL inst_4_27 ( 
	.A1(out_sel[8]), 
	.A2(I8[27]), 
	.B1(out_sel[9]), 
	.B2(I9[27]), 
	.Z(O4[27])); 
	AO_CELL inst_5_27 ( 
	.A1(out_sel[10]), 
	.A2(I10[27]), 
	.B1(out_sel[11]), 
	.B2(I11[27]), 
	.Z(O5[27])); 
	AO_CELL inst_6_27 ( 
	.A1(out_sel[12]), 
	.A2(I12[27]), 
	.B1(out_sel[13]), 
	.B2(I13[27]), 
	.Z(O6[27])); 
	AO_CELL inst_7_27 ( 
	.A1(out_sel[14]), 
	.A2(I14[27]), 
	.B1(out_sel[15]), 
	.B2(I15[27]), 
	.Z(O7[27])); 
	AO_CELL inst_8_27 ( 
	.A1(out_sel[16]), 
	.A2(I16[27]), 
	.B1(out_sel[17]), 
	.B2(I17[27]), 
	.Z(O8[27])); 
	AO_CELL inst_0_28 ( 
	.A1(out_sel[0]), 
	.A2(I0[28]), 
	.B1(out_sel[1]), 
	.B2(I1[28]), 
	.Z(O0[28])); 
	AO_CELL inst_1_28 ( 
	.A1(out_sel[2]), 
	.A2(I2[28]), 
	.B1(out_sel[3]), 
	.B2(I3[28]), 
	.Z(O1[28])); 
	AO_CELL inst_2_28 ( 
	.A1(out_sel[4]), 
	.A2(I4[28]), 
	.B1(out_sel[5]), 
	.B2(I5[28]), 
	.Z(O2[28])); 
	AO_CELL inst_3_28 ( 
	.A1(out_sel[6]), 
	.A2(I6[28]), 
	.B1(out_sel[7]), 
	.B2(I7[28]), 
	.Z(O3[28])); 
	AO_CELL inst_4_28 ( 
	.A1(out_sel[8]), 
	.A2(I8[28]), 
	.B1(out_sel[9]), 
	.B2(I9[28]), 
	.Z(O4[28])); 
	AO_CELL inst_5_28 ( 
	.A1(out_sel[10]), 
	.A2(I10[28]), 
	.B1(out_sel[11]), 
	.B2(I11[28]), 
	.Z(O5[28])); 
	AO_CELL inst_6_28 ( 
	.A1(out_sel[12]), 
	.A2(I12[28]), 
	.B1(out_sel[13]), 
	.B2(I13[28]), 
	.Z(O6[28])); 
	AO_CELL inst_7_28 ( 
	.A1(out_sel[14]), 
	.A2(I14[28]), 
	.B1(out_sel[15]), 
	.B2(I15[28]), 
	.Z(O7[28])); 
	AO_CELL inst_8_28 ( 
	.A1(out_sel[16]), 
	.A2(I16[28]), 
	.B1(out_sel[17]), 
	.B2(I17[28]), 
	.Z(O8[28])); 
	AO_CELL inst_0_29 ( 
	.A1(out_sel[0]), 
	.A2(I0[29]), 
	.B1(out_sel[1]), 
	.B2(I1[29]), 
	.Z(O0[29])); 
	AO_CELL inst_1_29 ( 
	.A1(out_sel[2]), 
	.A2(I2[29]), 
	.B1(out_sel[3]), 
	.B2(I3[29]), 
	.Z(O1[29])); 
	AO_CELL inst_2_29 ( 
	.A1(out_sel[4]), 
	.A2(I4[29]), 
	.B1(out_sel[5]), 
	.B2(I5[29]), 
	.Z(O2[29])); 
	AO_CELL inst_3_29 ( 
	.A1(out_sel[6]), 
	.A2(I6[29]), 
	.B1(out_sel[7]), 
	.B2(I7[29]), 
	.Z(O3[29])); 
	AO_CELL inst_4_29 ( 
	.A1(out_sel[8]), 
	.A2(I8[29]), 
	.B1(out_sel[9]), 
	.B2(I9[29]), 
	.Z(O4[29])); 
	AO_CELL inst_5_29 ( 
	.A1(out_sel[10]), 
	.A2(I10[29]), 
	.B1(out_sel[11]), 
	.B2(I11[29]), 
	.Z(O5[29])); 
	AO_CELL inst_6_29 ( 
	.A1(out_sel[12]), 
	.A2(I12[29]), 
	.B1(out_sel[13]), 
	.B2(I13[29]), 
	.Z(O6[29])); 
	AO_CELL inst_7_29 ( 
	.A1(out_sel[14]), 
	.A2(I14[29]), 
	.B1(out_sel[15]), 
	.B2(I15[29]), 
	.Z(O7[29])); 
	AO_CELL inst_8_29 ( 
	.A1(out_sel[16]), 
	.A2(I16[29]), 
	.B1(out_sel[17]), 
	.B2(I17[29]), 
	.Z(O8[29])); 
	AO_CELL inst_0_30 ( 
	.A1(out_sel[0]), 
	.A2(I0[30]), 
	.B1(out_sel[1]), 
	.B2(I1[30]), 
	.Z(O0[30])); 
	AO_CELL inst_1_30 ( 
	.A1(out_sel[2]), 
	.A2(I2[30]), 
	.B1(out_sel[3]), 
	.B2(I3[30]), 
	.Z(O1[30])); 
	AO_CELL inst_2_30 ( 
	.A1(out_sel[4]), 
	.A2(I4[30]), 
	.B1(out_sel[5]), 
	.B2(I5[30]), 
	.Z(O2[30])); 
	AO_CELL inst_3_30 ( 
	.A1(out_sel[6]), 
	.A2(I6[30]), 
	.B1(out_sel[7]), 
	.B2(I7[30]), 
	.Z(O3[30])); 
	AO_CELL inst_4_30 ( 
	.A1(out_sel[8]), 
	.A2(I8[30]), 
	.B1(out_sel[9]), 
	.B2(I9[30]), 
	.Z(O4[30])); 
	AO_CELL inst_5_30 ( 
	.A1(out_sel[10]), 
	.A2(I10[30]), 
	.B1(out_sel[11]), 
	.B2(I11[30]), 
	.Z(O5[30])); 
	AO_CELL inst_6_30 ( 
	.A1(out_sel[12]), 
	.A2(I12[30]), 
	.B1(out_sel[13]), 
	.B2(I13[30]), 
	.Z(O6[30])); 
	AO_CELL inst_7_30 ( 
	.A1(out_sel[14]), 
	.A2(I14[30]), 
	.B1(out_sel[15]), 
	.B2(I15[30]), 
	.Z(O7[30])); 
	AO_CELL inst_8_30 ( 
	.A1(out_sel[16]), 
	.A2(I16[30]), 
	.B1(out_sel[17]), 
	.B2(I17[30]), 
	.Z(O8[30])); 
	AO_CELL inst_0_31 ( 
	.A1(out_sel[0]), 
	.A2(I0[31]), 
	.B1(out_sel[1]), 
	.B2(I1[31]), 
	.Z(O0[31])); 
	AO_CELL inst_1_31 ( 
	.A1(out_sel[2]), 
	.A2(I2[31]), 
	.B1(out_sel[3]), 
	.B2(I3[31]), 
	.Z(O1[31])); 
	AO_CELL inst_2_31 ( 
	.A1(out_sel[4]), 
	.A2(I4[31]), 
	.B1(out_sel[5]), 
	.B2(I5[31]), 
	.Z(O2[31])); 
	AO_CELL inst_3_31 ( 
	.A1(out_sel[6]), 
	.A2(I6[31]), 
	.B1(out_sel[7]), 
	.B2(I7[31]), 
	.Z(O3[31])); 
	AO_CELL inst_4_31 ( 
	.A1(out_sel[8]), 
	.A2(I8[31]), 
	.B1(out_sel[9]), 
	.B2(I9[31]), 
	.Z(O4[31])); 
	AO_CELL inst_5_31 ( 
	.A1(out_sel[10]), 
	.A2(I10[31]), 
	.B1(out_sel[11]), 
	.B2(I11[31]), 
	.Z(O5[31])); 
	AO_CELL inst_6_31 ( 
	.A1(out_sel[12]), 
	.A2(I12[31]), 
	.B1(out_sel[13]), 
	.B2(I13[31]), 
	.Z(O6[31])); 
	AO_CELL inst_7_31 ( 
	.A1(out_sel[14]), 
	.A2(I14[31]), 
	.B1(out_sel[15]), 
	.B2(I15[31]), 
	.Z(O7[31])); 
	AO_CELL inst_8_31 ( 
	.A1(out_sel[16]), 
	.A2(I16[31]), 
	.B1(out_sel[17]), 
	.B2(I17[31]), 
	.Z(O8[31])); 
endmodule 

module mux_aoi_16_32 ( 
	input logic  [31 : 0] I[15:0], 
	input logic  [3 : 0] S ,
	output logic  [15 : 0] out_sel,
	output logic [31 : 0] O); 
	logic  [31 : 0] O_int0;
	logic  [31 : 0] O_int1;
	logic  [31 : 0] O_int2;
	logic  [31 : 0] O_int3;
	logic  [31 : 0] O_int4;
	logic  [31 : 0] O_int5;
	logic  [31 : 0] O_int6;
	logic  [31 : 0] O_int7;

precoder_32_16 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_32_16 u_mux_logic ( 
	.I0 (I[0]),
	.I1 (I[1]),
	.I2 (I[2]),
	.I3 (I[3]),
	.I4 (I[4]),
	.I5 (I[5]),
	.I6 (I[6]),
	.I7 (I[7]),
	.I8 (I[8]),
	.I9 (I[9]),
	.I10 (I[10]),
	.I11 (I[11]),
	.I12 (I[12]),
	.I13 (I[13]),
	.I14 (I[14]),
	.I15 (I[15]),
	.out_sel(out_sel), 
	.O0(O_int0), 
	.O1(O_int1), 
	.O2(O_int2), 
	.O3(O_int3), 
	.O4(O_int4), 
	.O5(O_int5), 
	.O6(O_int6), 
	.O7(O_int7)); 
	assign O = (  	O_int0 | 	O_int1 | 	O_int2 | 	O_int3 | 	O_int4 | 	O_int5 | 	O_int6 | 	O_int7 	); 

endmodule 

module precoder_32_16 (
	input logic  [3 : 0] S ,
	output logic  [15 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		4'd0    :   out_sel = 16'b0000000000000001;
		4'd1    :   out_sel = 16'b0000000000000010;
		4'd2    :   out_sel = 16'b0000000000000100;
		4'd3    :   out_sel = 16'b0000000000001000;
		4'd4    :   out_sel = 16'b0000000000010000;
		4'd5    :   out_sel = 16'b0000000000100000;
		4'd6    :   out_sel = 16'b0000000001000000;
		4'd7    :   out_sel = 16'b0000000010000000;
		4'd8    :   out_sel = 16'b0000000100000000;
		4'd9    :   out_sel = 16'b0000001000000000;
		4'd10    :   out_sel = 16'b0000010000000000;
		4'd11    :   out_sel = 16'b0000100000000000;
		4'd12    :   out_sel = 16'b0001000000000000;
		4'd13    :   out_sel = 16'b0010000000000000;
		4'd14    :   out_sel = 16'b0100000000000000;
		4'd15    :   out_sel = 16'b1000000000000000;
		default :   out_sel = 16'b0;
	endcase 
end 

endmodule 

module mux_logic_32_16 ( 
	input logic  [15 : 0] out_sel,
	input logic  [31 : 0] I0, 
	input logic  [31 : 0] I1, 
	input logic  [31 : 0] I2, 
	input logic  [31 : 0] I3, 
	input logic  [31 : 0] I4, 
	input logic  [31 : 0] I5, 
	input logic  [31 : 0] I6, 
	input logic  [31 : 0] I7, 
	input logic  [31 : 0] I8, 
	input logic  [31 : 0] I9, 
	input logic  [31 : 0] I10, 
	input logic  [31 : 0] I11, 
	input logic  [31 : 0] I12, 
	input logic  [31 : 0] I13, 
	input logic  [31 : 0] I14, 
	input logic  [31 : 0] I15, 
	output logic  [31 : 0] O0, 
	output logic  [31 : 0] O1, 
	output logic  [31 : 0] O2, 
	output logic  [31 : 0] O3, 
	output logic  [31 : 0] O4, 
	output logic  [31 : 0] O5, 
	output logic  [31 : 0] O6, 
	output logic  [31 : 0] O7); 
	AO_CELL inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	AO_CELL inst_1_0 ( 
	.A1(out_sel[2]), 
	.A2(I2[0]), 
	.B1(out_sel[3]), 
	.B2(I3[0]), 
	.Z(O1[0])); 
	AO_CELL inst_2_0 ( 
	.A1(out_sel[4]), 
	.A2(I4[0]), 
	.B1(out_sel[5]), 
	.B2(I5[0]), 
	.Z(O2[0])); 
	AO_CELL inst_3_0 ( 
	.A1(out_sel[6]), 
	.A2(I6[0]), 
	.B1(out_sel[7]), 
	.B2(I7[0]), 
	.Z(O3[0])); 
	AO_CELL inst_4_0 ( 
	.A1(out_sel[8]), 
	.A2(I8[0]), 
	.B1(out_sel[9]), 
	.B2(I9[0]), 
	.Z(O4[0])); 
	AO_CELL inst_5_0 ( 
	.A1(out_sel[10]), 
	.A2(I10[0]), 
	.B1(out_sel[11]), 
	.B2(I11[0]), 
	.Z(O5[0])); 
	AO_CELL inst_6_0 ( 
	.A1(out_sel[12]), 
	.A2(I12[0]), 
	.B1(out_sel[13]), 
	.B2(I13[0]), 
	.Z(O6[0])); 
	AO_CELL inst_7_0 ( 
	.A1(out_sel[14]), 
	.A2(I14[0]), 
	.B1(out_sel[15]), 
	.B2(I15[0]), 
	.Z(O7[0])); 
	AO_CELL inst_0_1 ( 
	.A1(out_sel[0]), 
	.A2(I0[1]), 
	.B1(out_sel[1]), 
	.B2(I1[1]), 
	.Z(O0[1])); 
	AO_CELL inst_1_1 ( 
	.A1(out_sel[2]), 
	.A2(I2[1]), 
	.B1(out_sel[3]), 
	.B2(I3[1]), 
	.Z(O1[1])); 
	AO_CELL inst_2_1 ( 
	.A1(out_sel[4]), 
	.A2(I4[1]), 
	.B1(out_sel[5]), 
	.B2(I5[1]), 
	.Z(O2[1])); 
	AO_CELL inst_3_1 ( 
	.A1(out_sel[6]), 
	.A2(I6[1]), 
	.B1(out_sel[7]), 
	.B2(I7[1]), 
	.Z(O3[1])); 
	AO_CELL inst_4_1 ( 
	.A1(out_sel[8]), 
	.A2(I8[1]), 
	.B1(out_sel[9]), 
	.B2(I9[1]), 
	.Z(O4[1])); 
	AO_CELL inst_5_1 ( 
	.A1(out_sel[10]), 
	.A2(I10[1]), 
	.B1(out_sel[11]), 
	.B2(I11[1]), 
	.Z(O5[1])); 
	AO_CELL inst_6_1 ( 
	.A1(out_sel[12]), 
	.A2(I12[1]), 
	.B1(out_sel[13]), 
	.B2(I13[1]), 
	.Z(O6[1])); 
	AO_CELL inst_7_1 ( 
	.A1(out_sel[14]), 
	.A2(I14[1]), 
	.B1(out_sel[15]), 
	.B2(I15[1]), 
	.Z(O7[1])); 
	AO_CELL inst_0_2 ( 
	.A1(out_sel[0]), 
	.A2(I0[2]), 
	.B1(out_sel[1]), 
	.B2(I1[2]), 
	.Z(O0[2])); 
	AO_CELL inst_1_2 ( 
	.A1(out_sel[2]), 
	.A2(I2[2]), 
	.B1(out_sel[3]), 
	.B2(I3[2]), 
	.Z(O1[2])); 
	AO_CELL inst_2_2 ( 
	.A1(out_sel[4]), 
	.A2(I4[2]), 
	.B1(out_sel[5]), 
	.B2(I5[2]), 
	.Z(O2[2])); 
	AO_CELL inst_3_2 ( 
	.A1(out_sel[6]), 
	.A2(I6[2]), 
	.B1(out_sel[7]), 
	.B2(I7[2]), 
	.Z(O3[2])); 
	AO_CELL inst_4_2 ( 
	.A1(out_sel[8]), 
	.A2(I8[2]), 
	.B1(out_sel[9]), 
	.B2(I9[2]), 
	.Z(O4[2])); 
	AO_CELL inst_5_2 ( 
	.A1(out_sel[10]), 
	.A2(I10[2]), 
	.B1(out_sel[11]), 
	.B2(I11[2]), 
	.Z(O5[2])); 
	AO_CELL inst_6_2 ( 
	.A1(out_sel[12]), 
	.A2(I12[2]), 
	.B1(out_sel[13]), 
	.B2(I13[2]), 
	.Z(O6[2])); 
	AO_CELL inst_7_2 ( 
	.A1(out_sel[14]), 
	.A2(I14[2]), 
	.B1(out_sel[15]), 
	.B2(I15[2]), 
	.Z(O7[2])); 
	AO_CELL inst_0_3 ( 
	.A1(out_sel[0]), 
	.A2(I0[3]), 
	.B1(out_sel[1]), 
	.B2(I1[3]), 
	.Z(O0[3])); 
	AO_CELL inst_1_3 ( 
	.A1(out_sel[2]), 
	.A2(I2[3]), 
	.B1(out_sel[3]), 
	.B2(I3[3]), 
	.Z(O1[3])); 
	AO_CELL inst_2_3 ( 
	.A1(out_sel[4]), 
	.A2(I4[3]), 
	.B1(out_sel[5]), 
	.B2(I5[3]), 
	.Z(O2[3])); 
	AO_CELL inst_3_3 ( 
	.A1(out_sel[6]), 
	.A2(I6[3]), 
	.B1(out_sel[7]), 
	.B2(I7[3]), 
	.Z(O3[3])); 
	AO_CELL inst_4_3 ( 
	.A1(out_sel[8]), 
	.A2(I8[3]), 
	.B1(out_sel[9]), 
	.B2(I9[3]), 
	.Z(O4[3])); 
	AO_CELL inst_5_3 ( 
	.A1(out_sel[10]), 
	.A2(I10[3]), 
	.B1(out_sel[11]), 
	.B2(I11[3]), 
	.Z(O5[3])); 
	AO_CELL inst_6_3 ( 
	.A1(out_sel[12]), 
	.A2(I12[3]), 
	.B1(out_sel[13]), 
	.B2(I13[3]), 
	.Z(O6[3])); 
	AO_CELL inst_7_3 ( 
	.A1(out_sel[14]), 
	.A2(I14[3]), 
	.B1(out_sel[15]), 
	.B2(I15[3]), 
	.Z(O7[3])); 
	AO_CELL inst_0_4 ( 
	.A1(out_sel[0]), 
	.A2(I0[4]), 
	.B1(out_sel[1]), 
	.B2(I1[4]), 
	.Z(O0[4])); 
	AO_CELL inst_1_4 ( 
	.A1(out_sel[2]), 
	.A2(I2[4]), 
	.B1(out_sel[3]), 
	.B2(I3[4]), 
	.Z(O1[4])); 
	AO_CELL inst_2_4 ( 
	.A1(out_sel[4]), 
	.A2(I4[4]), 
	.B1(out_sel[5]), 
	.B2(I5[4]), 
	.Z(O2[4])); 
	AO_CELL inst_3_4 ( 
	.A1(out_sel[6]), 
	.A2(I6[4]), 
	.B1(out_sel[7]), 
	.B2(I7[4]), 
	.Z(O3[4])); 
	AO_CELL inst_4_4 ( 
	.A1(out_sel[8]), 
	.A2(I8[4]), 
	.B1(out_sel[9]), 
	.B2(I9[4]), 
	.Z(O4[4])); 
	AO_CELL inst_5_4 ( 
	.A1(out_sel[10]), 
	.A2(I10[4]), 
	.B1(out_sel[11]), 
	.B2(I11[4]), 
	.Z(O5[4])); 
	AO_CELL inst_6_4 ( 
	.A1(out_sel[12]), 
	.A2(I12[4]), 
	.B1(out_sel[13]), 
	.B2(I13[4]), 
	.Z(O6[4])); 
	AO_CELL inst_7_4 ( 
	.A1(out_sel[14]), 
	.A2(I14[4]), 
	.B1(out_sel[15]), 
	.B2(I15[4]), 
	.Z(O7[4])); 
	AO_CELL inst_0_5 ( 
	.A1(out_sel[0]), 
	.A2(I0[5]), 
	.B1(out_sel[1]), 
	.B2(I1[5]), 
	.Z(O0[5])); 
	AO_CELL inst_1_5 ( 
	.A1(out_sel[2]), 
	.A2(I2[5]), 
	.B1(out_sel[3]), 
	.B2(I3[5]), 
	.Z(O1[5])); 
	AO_CELL inst_2_5 ( 
	.A1(out_sel[4]), 
	.A2(I4[5]), 
	.B1(out_sel[5]), 
	.B2(I5[5]), 
	.Z(O2[5])); 
	AO_CELL inst_3_5 ( 
	.A1(out_sel[6]), 
	.A2(I6[5]), 
	.B1(out_sel[7]), 
	.B2(I7[5]), 
	.Z(O3[5])); 
	AO_CELL inst_4_5 ( 
	.A1(out_sel[8]), 
	.A2(I8[5]), 
	.B1(out_sel[9]), 
	.B2(I9[5]), 
	.Z(O4[5])); 
	AO_CELL inst_5_5 ( 
	.A1(out_sel[10]), 
	.A2(I10[5]), 
	.B1(out_sel[11]), 
	.B2(I11[5]), 
	.Z(O5[5])); 
	AO_CELL inst_6_5 ( 
	.A1(out_sel[12]), 
	.A2(I12[5]), 
	.B1(out_sel[13]), 
	.B2(I13[5]), 
	.Z(O6[5])); 
	AO_CELL inst_7_5 ( 
	.A1(out_sel[14]), 
	.A2(I14[5]), 
	.B1(out_sel[15]), 
	.B2(I15[5]), 
	.Z(O7[5])); 
	AO_CELL inst_0_6 ( 
	.A1(out_sel[0]), 
	.A2(I0[6]), 
	.B1(out_sel[1]), 
	.B2(I1[6]), 
	.Z(O0[6])); 
	AO_CELL inst_1_6 ( 
	.A1(out_sel[2]), 
	.A2(I2[6]), 
	.B1(out_sel[3]), 
	.B2(I3[6]), 
	.Z(O1[6])); 
	AO_CELL inst_2_6 ( 
	.A1(out_sel[4]), 
	.A2(I4[6]), 
	.B1(out_sel[5]), 
	.B2(I5[6]), 
	.Z(O2[6])); 
	AO_CELL inst_3_6 ( 
	.A1(out_sel[6]), 
	.A2(I6[6]), 
	.B1(out_sel[7]), 
	.B2(I7[6]), 
	.Z(O3[6])); 
	AO_CELL inst_4_6 ( 
	.A1(out_sel[8]), 
	.A2(I8[6]), 
	.B1(out_sel[9]), 
	.B2(I9[6]), 
	.Z(O4[6])); 
	AO_CELL inst_5_6 ( 
	.A1(out_sel[10]), 
	.A2(I10[6]), 
	.B1(out_sel[11]), 
	.B2(I11[6]), 
	.Z(O5[6])); 
	AO_CELL inst_6_6 ( 
	.A1(out_sel[12]), 
	.A2(I12[6]), 
	.B1(out_sel[13]), 
	.B2(I13[6]), 
	.Z(O6[6])); 
	AO_CELL inst_7_6 ( 
	.A1(out_sel[14]), 
	.A2(I14[6]), 
	.B1(out_sel[15]), 
	.B2(I15[6]), 
	.Z(O7[6])); 
	AO_CELL inst_0_7 ( 
	.A1(out_sel[0]), 
	.A2(I0[7]), 
	.B1(out_sel[1]), 
	.B2(I1[7]), 
	.Z(O0[7])); 
	AO_CELL inst_1_7 ( 
	.A1(out_sel[2]), 
	.A2(I2[7]), 
	.B1(out_sel[3]), 
	.B2(I3[7]), 
	.Z(O1[7])); 
	AO_CELL inst_2_7 ( 
	.A1(out_sel[4]), 
	.A2(I4[7]), 
	.B1(out_sel[5]), 
	.B2(I5[7]), 
	.Z(O2[7])); 
	AO_CELL inst_3_7 ( 
	.A1(out_sel[6]), 
	.A2(I6[7]), 
	.B1(out_sel[7]), 
	.B2(I7[7]), 
	.Z(O3[7])); 
	AO_CELL inst_4_7 ( 
	.A1(out_sel[8]), 
	.A2(I8[7]), 
	.B1(out_sel[9]), 
	.B2(I9[7]), 
	.Z(O4[7])); 
	AO_CELL inst_5_7 ( 
	.A1(out_sel[10]), 
	.A2(I10[7]), 
	.B1(out_sel[11]), 
	.B2(I11[7]), 
	.Z(O5[7])); 
	AO_CELL inst_6_7 ( 
	.A1(out_sel[12]), 
	.A2(I12[7]), 
	.B1(out_sel[13]), 
	.B2(I13[7]), 
	.Z(O6[7])); 
	AO_CELL inst_7_7 ( 
	.A1(out_sel[14]), 
	.A2(I14[7]), 
	.B1(out_sel[15]), 
	.B2(I15[7]), 
	.Z(O7[7])); 
	AO_CELL inst_0_8 ( 
	.A1(out_sel[0]), 
	.A2(I0[8]), 
	.B1(out_sel[1]), 
	.B2(I1[8]), 
	.Z(O0[8])); 
	AO_CELL inst_1_8 ( 
	.A1(out_sel[2]), 
	.A2(I2[8]), 
	.B1(out_sel[3]), 
	.B2(I3[8]), 
	.Z(O1[8])); 
	AO_CELL inst_2_8 ( 
	.A1(out_sel[4]), 
	.A2(I4[8]), 
	.B1(out_sel[5]), 
	.B2(I5[8]), 
	.Z(O2[8])); 
	AO_CELL inst_3_8 ( 
	.A1(out_sel[6]), 
	.A2(I6[8]), 
	.B1(out_sel[7]), 
	.B2(I7[8]), 
	.Z(O3[8])); 
	AO_CELL inst_4_8 ( 
	.A1(out_sel[8]), 
	.A2(I8[8]), 
	.B1(out_sel[9]), 
	.B2(I9[8]), 
	.Z(O4[8])); 
	AO_CELL inst_5_8 ( 
	.A1(out_sel[10]), 
	.A2(I10[8]), 
	.B1(out_sel[11]), 
	.B2(I11[8]), 
	.Z(O5[8])); 
	AO_CELL inst_6_8 ( 
	.A1(out_sel[12]), 
	.A2(I12[8]), 
	.B1(out_sel[13]), 
	.B2(I13[8]), 
	.Z(O6[8])); 
	AO_CELL inst_7_8 ( 
	.A1(out_sel[14]), 
	.A2(I14[8]), 
	.B1(out_sel[15]), 
	.B2(I15[8]), 
	.Z(O7[8])); 
	AO_CELL inst_0_9 ( 
	.A1(out_sel[0]), 
	.A2(I0[9]), 
	.B1(out_sel[1]), 
	.B2(I1[9]), 
	.Z(O0[9])); 
	AO_CELL inst_1_9 ( 
	.A1(out_sel[2]), 
	.A2(I2[9]), 
	.B1(out_sel[3]), 
	.B2(I3[9]), 
	.Z(O1[9])); 
	AO_CELL inst_2_9 ( 
	.A1(out_sel[4]), 
	.A2(I4[9]), 
	.B1(out_sel[5]), 
	.B2(I5[9]), 
	.Z(O2[9])); 
	AO_CELL inst_3_9 ( 
	.A1(out_sel[6]), 
	.A2(I6[9]), 
	.B1(out_sel[7]), 
	.B2(I7[9]), 
	.Z(O3[9])); 
	AO_CELL inst_4_9 ( 
	.A1(out_sel[8]), 
	.A2(I8[9]), 
	.B1(out_sel[9]), 
	.B2(I9[9]), 
	.Z(O4[9])); 
	AO_CELL inst_5_9 ( 
	.A1(out_sel[10]), 
	.A2(I10[9]), 
	.B1(out_sel[11]), 
	.B2(I11[9]), 
	.Z(O5[9])); 
	AO_CELL inst_6_9 ( 
	.A1(out_sel[12]), 
	.A2(I12[9]), 
	.B1(out_sel[13]), 
	.B2(I13[9]), 
	.Z(O6[9])); 
	AO_CELL inst_7_9 ( 
	.A1(out_sel[14]), 
	.A2(I14[9]), 
	.B1(out_sel[15]), 
	.B2(I15[9]), 
	.Z(O7[9])); 
	AO_CELL inst_0_10 ( 
	.A1(out_sel[0]), 
	.A2(I0[10]), 
	.B1(out_sel[1]), 
	.B2(I1[10]), 
	.Z(O0[10])); 
	AO_CELL inst_1_10 ( 
	.A1(out_sel[2]), 
	.A2(I2[10]), 
	.B1(out_sel[3]), 
	.B2(I3[10]), 
	.Z(O1[10])); 
	AO_CELL inst_2_10 ( 
	.A1(out_sel[4]), 
	.A2(I4[10]), 
	.B1(out_sel[5]), 
	.B2(I5[10]), 
	.Z(O2[10])); 
	AO_CELL inst_3_10 ( 
	.A1(out_sel[6]), 
	.A2(I6[10]), 
	.B1(out_sel[7]), 
	.B2(I7[10]), 
	.Z(O3[10])); 
	AO_CELL inst_4_10 ( 
	.A1(out_sel[8]), 
	.A2(I8[10]), 
	.B1(out_sel[9]), 
	.B2(I9[10]), 
	.Z(O4[10])); 
	AO_CELL inst_5_10 ( 
	.A1(out_sel[10]), 
	.A2(I10[10]), 
	.B1(out_sel[11]), 
	.B2(I11[10]), 
	.Z(O5[10])); 
	AO_CELL inst_6_10 ( 
	.A1(out_sel[12]), 
	.A2(I12[10]), 
	.B1(out_sel[13]), 
	.B2(I13[10]), 
	.Z(O6[10])); 
	AO_CELL inst_7_10 ( 
	.A1(out_sel[14]), 
	.A2(I14[10]), 
	.B1(out_sel[15]), 
	.B2(I15[10]), 
	.Z(O7[10])); 
	AO_CELL inst_0_11 ( 
	.A1(out_sel[0]), 
	.A2(I0[11]), 
	.B1(out_sel[1]), 
	.B2(I1[11]), 
	.Z(O0[11])); 
	AO_CELL inst_1_11 ( 
	.A1(out_sel[2]), 
	.A2(I2[11]), 
	.B1(out_sel[3]), 
	.B2(I3[11]), 
	.Z(O1[11])); 
	AO_CELL inst_2_11 ( 
	.A1(out_sel[4]), 
	.A2(I4[11]), 
	.B1(out_sel[5]), 
	.B2(I5[11]), 
	.Z(O2[11])); 
	AO_CELL inst_3_11 ( 
	.A1(out_sel[6]), 
	.A2(I6[11]), 
	.B1(out_sel[7]), 
	.B2(I7[11]), 
	.Z(O3[11])); 
	AO_CELL inst_4_11 ( 
	.A1(out_sel[8]), 
	.A2(I8[11]), 
	.B1(out_sel[9]), 
	.B2(I9[11]), 
	.Z(O4[11])); 
	AO_CELL inst_5_11 ( 
	.A1(out_sel[10]), 
	.A2(I10[11]), 
	.B1(out_sel[11]), 
	.B2(I11[11]), 
	.Z(O5[11])); 
	AO_CELL inst_6_11 ( 
	.A1(out_sel[12]), 
	.A2(I12[11]), 
	.B1(out_sel[13]), 
	.B2(I13[11]), 
	.Z(O6[11])); 
	AO_CELL inst_7_11 ( 
	.A1(out_sel[14]), 
	.A2(I14[11]), 
	.B1(out_sel[15]), 
	.B2(I15[11]), 
	.Z(O7[11])); 
	AO_CELL inst_0_12 ( 
	.A1(out_sel[0]), 
	.A2(I0[12]), 
	.B1(out_sel[1]), 
	.B2(I1[12]), 
	.Z(O0[12])); 
	AO_CELL inst_1_12 ( 
	.A1(out_sel[2]), 
	.A2(I2[12]), 
	.B1(out_sel[3]), 
	.B2(I3[12]), 
	.Z(O1[12])); 
	AO_CELL inst_2_12 ( 
	.A1(out_sel[4]), 
	.A2(I4[12]), 
	.B1(out_sel[5]), 
	.B2(I5[12]), 
	.Z(O2[12])); 
	AO_CELL inst_3_12 ( 
	.A1(out_sel[6]), 
	.A2(I6[12]), 
	.B1(out_sel[7]), 
	.B2(I7[12]), 
	.Z(O3[12])); 
	AO_CELL inst_4_12 ( 
	.A1(out_sel[8]), 
	.A2(I8[12]), 
	.B1(out_sel[9]), 
	.B2(I9[12]), 
	.Z(O4[12])); 
	AO_CELL inst_5_12 ( 
	.A1(out_sel[10]), 
	.A2(I10[12]), 
	.B1(out_sel[11]), 
	.B2(I11[12]), 
	.Z(O5[12])); 
	AO_CELL inst_6_12 ( 
	.A1(out_sel[12]), 
	.A2(I12[12]), 
	.B1(out_sel[13]), 
	.B2(I13[12]), 
	.Z(O6[12])); 
	AO_CELL inst_7_12 ( 
	.A1(out_sel[14]), 
	.A2(I14[12]), 
	.B1(out_sel[15]), 
	.B2(I15[12]), 
	.Z(O7[12])); 
	AO_CELL inst_0_13 ( 
	.A1(out_sel[0]), 
	.A2(I0[13]), 
	.B1(out_sel[1]), 
	.B2(I1[13]), 
	.Z(O0[13])); 
	AO_CELL inst_1_13 ( 
	.A1(out_sel[2]), 
	.A2(I2[13]), 
	.B1(out_sel[3]), 
	.B2(I3[13]), 
	.Z(O1[13])); 
	AO_CELL inst_2_13 ( 
	.A1(out_sel[4]), 
	.A2(I4[13]), 
	.B1(out_sel[5]), 
	.B2(I5[13]), 
	.Z(O2[13])); 
	AO_CELL inst_3_13 ( 
	.A1(out_sel[6]), 
	.A2(I6[13]), 
	.B1(out_sel[7]), 
	.B2(I7[13]), 
	.Z(O3[13])); 
	AO_CELL inst_4_13 ( 
	.A1(out_sel[8]), 
	.A2(I8[13]), 
	.B1(out_sel[9]), 
	.B2(I9[13]), 
	.Z(O4[13])); 
	AO_CELL inst_5_13 ( 
	.A1(out_sel[10]), 
	.A2(I10[13]), 
	.B1(out_sel[11]), 
	.B2(I11[13]), 
	.Z(O5[13])); 
	AO_CELL inst_6_13 ( 
	.A1(out_sel[12]), 
	.A2(I12[13]), 
	.B1(out_sel[13]), 
	.B2(I13[13]), 
	.Z(O6[13])); 
	AO_CELL inst_7_13 ( 
	.A1(out_sel[14]), 
	.A2(I14[13]), 
	.B1(out_sel[15]), 
	.B2(I15[13]), 
	.Z(O7[13])); 
	AO_CELL inst_0_14 ( 
	.A1(out_sel[0]), 
	.A2(I0[14]), 
	.B1(out_sel[1]), 
	.B2(I1[14]), 
	.Z(O0[14])); 
	AO_CELL inst_1_14 ( 
	.A1(out_sel[2]), 
	.A2(I2[14]), 
	.B1(out_sel[3]), 
	.B2(I3[14]), 
	.Z(O1[14])); 
	AO_CELL inst_2_14 ( 
	.A1(out_sel[4]), 
	.A2(I4[14]), 
	.B1(out_sel[5]), 
	.B2(I5[14]), 
	.Z(O2[14])); 
	AO_CELL inst_3_14 ( 
	.A1(out_sel[6]), 
	.A2(I6[14]), 
	.B1(out_sel[7]), 
	.B2(I7[14]), 
	.Z(O3[14])); 
	AO_CELL inst_4_14 ( 
	.A1(out_sel[8]), 
	.A2(I8[14]), 
	.B1(out_sel[9]), 
	.B2(I9[14]), 
	.Z(O4[14])); 
	AO_CELL inst_5_14 ( 
	.A1(out_sel[10]), 
	.A2(I10[14]), 
	.B1(out_sel[11]), 
	.B2(I11[14]), 
	.Z(O5[14])); 
	AO_CELL inst_6_14 ( 
	.A1(out_sel[12]), 
	.A2(I12[14]), 
	.B1(out_sel[13]), 
	.B2(I13[14]), 
	.Z(O6[14])); 
	AO_CELL inst_7_14 ( 
	.A1(out_sel[14]), 
	.A2(I14[14]), 
	.B1(out_sel[15]), 
	.B2(I15[14]), 
	.Z(O7[14])); 
	AO_CELL inst_0_15 ( 
	.A1(out_sel[0]), 
	.A2(I0[15]), 
	.B1(out_sel[1]), 
	.B2(I1[15]), 
	.Z(O0[15])); 
	AO_CELL inst_1_15 ( 
	.A1(out_sel[2]), 
	.A2(I2[15]), 
	.B1(out_sel[3]), 
	.B2(I3[15]), 
	.Z(O1[15])); 
	AO_CELL inst_2_15 ( 
	.A1(out_sel[4]), 
	.A2(I4[15]), 
	.B1(out_sel[5]), 
	.B2(I5[15]), 
	.Z(O2[15])); 
	AO_CELL inst_3_15 ( 
	.A1(out_sel[6]), 
	.A2(I6[15]), 
	.B1(out_sel[7]), 
	.B2(I7[15]), 
	.Z(O3[15])); 
	AO_CELL inst_4_15 ( 
	.A1(out_sel[8]), 
	.A2(I8[15]), 
	.B1(out_sel[9]), 
	.B2(I9[15]), 
	.Z(O4[15])); 
	AO_CELL inst_5_15 ( 
	.A1(out_sel[10]), 
	.A2(I10[15]), 
	.B1(out_sel[11]), 
	.B2(I11[15]), 
	.Z(O5[15])); 
	AO_CELL inst_6_15 ( 
	.A1(out_sel[12]), 
	.A2(I12[15]), 
	.B1(out_sel[13]), 
	.B2(I13[15]), 
	.Z(O6[15])); 
	AO_CELL inst_7_15 ( 
	.A1(out_sel[14]), 
	.A2(I14[15]), 
	.B1(out_sel[15]), 
	.B2(I15[15]), 
	.Z(O7[15])); 
	AO_CELL inst_0_16 ( 
	.A1(out_sel[0]), 
	.A2(I0[16]), 
	.B1(out_sel[1]), 
	.B2(I1[16]), 
	.Z(O0[16])); 
	AO_CELL inst_1_16 ( 
	.A1(out_sel[2]), 
	.A2(I2[16]), 
	.B1(out_sel[3]), 
	.B2(I3[16]), 
	.Z(O1[16])); 
	AO_CELL inst_2_16 ( 
	.A1(out_sel[4]), 
	.A2(I4[16]), 
	.B1(out_sel[5]), 
	.B2(I5[16]), 
	.Z(O2[16])); 
	AO_CELL inst_3_16 ( 
	.A1(out_sel[6]), 
	.A2(I6[16]), 
	.B1(out_sel[7]), 
	.B2(I7[16]), 
	.Z(O3[16])); 
	AO_CELL inst_4_16 ( 
	.A1(out_sel[8]), 
	.A2(I8[16]), 
	.B1(out_sel[9]), 
	.B2(I9[16]), 
	.Z(O4[16])); 
	AO_CELL inst_5_16 ( 
	.A1(out_sel[10]), 
	.A2(I10[16]), 
	.B1(out_sel[11]), 
	.B2(I11[16]), 
	.Z(O5[16])); 
	AO_CELL inst_6_16 ( 
	.A1(out_sel[12]), 
	.A2(I12[16]), 
	.B1(out_sel[13]), 
	.B2(I13[16]), 
	.Z(O6[16])); 
	AO_CELL inst_7_16 ( 
	.A1(out_sel[14]), 
	.A2(I14[16]), 
	.B1(out_sel[15]), 
	.B2(I15[16]), 
	.Z(O7[16])); 
	AO_CELL inst_0_17 ( 
	.A1(out_sel[0]), 
	.A2(I0[17]), 
	.B1(out_sel[1]), 
	.B2(I1[17]), 
	.Z(O0[17])); 
	AO_CELL inst_1_17 ( 
	.A1(out_sel[2]), 
	.A2(I2[17]), 
	.B1(out_sel[3]), 
	.B2(I3[17]), 
	.Z(O1[17])); 
	AO_CELL inst_2_17 ( 
	.A1(out_sel[4]), 
	.A2(I4[17]), 
	.B1(out_sel[5]), 
	.B2(I5[17]), 
	.Z(O2[17])); 
	AO_CELL inst_3_17 ( 
	.A1(out_sel[6]), 
	.A2(I6[17]), 
	.B1(out_sel[7]), 
	.B2(I7[17]), 
	.Z(O3[17])); 
	AO_CELL inst_4_17 ( 
	.A1(out_sel[8]), 
	.A2(I8[17]), 
	.B1(out_sel[9]), 
	.B2(I9[17]), 
	.Z(O4[17])); 
	AO_CELL inst_5_17 ( 
	.A1(out_sel[10]), 
	.A2(I10[17]), 
	.B1(out_sel[11]), 
	.B2(I11[17]), 
	.Z(O5[17])); 
	AO_CELL inst_6_17 ( 
	.A1(out_sel[12]), 
	.A2(I12[17]), 
	.B1(out_sel[13]), 
	.B2(I13[17]), 
	.Z(O6[17])); 
	AO_CELL inst_7_17 ( 
	.A1(out_sel[14]), 
	.A2(I14[17]), 
	.B1(out_sel[15]), 
	.B2(I15[17]), 
	.Z(O7[17])); 
	AO_CELL inst_0_18 ( 
	.A1(out_sel[0]), 
	.A2(I0[18]), 
	.B1(out_sel[1]), 
	.B2(I1[18]), 
	.Z(O0[18])); 
	AO_CELL inst_1_18 ( 
	.A1(out_sel[2]), 
	.A2(I2[18]), 
	.B1(out_sel[3]), 
	.B2(I3[18]), 
	.Z(O1[18])); 
	AO_CELL inst_2_18 ( 
	.A1(out_sel[4]), 
	.A2(I4[18]), 
	.B1(out_sel[5]), 
	.B2(I5[18]), 
	.Z(O2[18])); 
	AO_CELL inst_3_18 ( 
	.A1(out_sel[6]), 
	.A2(I6[18]), 
	.B1(out_sel[7]), 
	.B2(I7[18]), 
	.Z(O3[18])); 
	AO_CELL inst_4_18 ( 
	.A1(out_sel[8]), 
	.A2(I8[18]), 
	.B1(out_sel[9]), 
	.B2(I9[18]), 
	.Z(O4[18])); 
	AO_CELL inst_5_18 ( 
	.A1(out_sel[10]), 
	.A2(I10[18]), 
	.B1(out_sel[11]), 
	.B2(I11[18]), 
	.Z(O5[18])); 
	AO_CELL inst_6_18 ( 
	.A1(out_sel[12]), 
	.A2(I12[18]), 
	.B1(out_sel[13]), 
	.B2(I13[18]), 
	.Z(O6[18])); 
	AO_CELL inst_7_18 ( 
	.A1(out_sel[14]), 
	.A2(I14[18]), 
	.B1(out_sel[15]), 
	.B2(I15[18]), 
	.Z(O7[18])); 
	AO_CELL inst_0_19 ( 
	.A1(out_sel[0]), 
	.A2(I0[19]), 
	.B1(out_sel[1]), 
	.B2(I1[19]), 
	.Z(O0[19])); 
	AO_CELL inst_1_19 ( 
	.A1(out_sel[2]), 
	.A2(I2[19]), 
	.B1(out_sel[3]), 
	.B2(I3[19]), 
	.Z(O1[19])); 
	AO_CELL inst_2_19 ( 
	.A1(out_sel[4]), 
	.A2(I4[19]), 
	.B1(out_sel[5]), 
	.B2(I5[19]), 
	.Z(O2[19])); 
	AO_CELL inst_3_19 ( 
	.A1(out_sel[6]), 
	.A2(I6[19]), 
	.B1(out_sel[7]), 
	.B2(I7[19]), 
	.Z(O3[19])); 
	AO_CELL inst_4_19 ( 
	.A1(out_sel[8]), 
	.A2(I8[19]), 
	.B1(out_sel[9]), 
	.B2(I9[19]), 
	.Z(O4[19])); 
	AO_CELL inst_5_19 ( 
	.A1(out_sel[10]), 
	.A2(I10[19]), 
	.B1(out_sel[11]), 
	.B2(I11[19]), 
	.Z(O5[19])); 
	AO_CELL inst_6_19 ( 
	.A1(out_sel[12]), 
	.A2(I12[19]), 
	.B1(out_sel[13]), 
	.B2(I13[19]), 
	.Z(O6[19])); 
	AO_CELL inst_7_19 ( 
	.A1(out_sel[14]), 
	.A2(I14[19]), 
	.B1(out_sel[15]), 
	.B2(I15[19]), 
	.Z(O7[19])); 
	AO_CELL inst_0_20 ( 
	.A1(out_sel[0]), 
	.A2(I0[20]), 
	.B1(out_sel[1]), 
	.B2(I1[20]), 
	.Z(O0[20])); 
	AO_CELL inst_1_20 ( 
	.A1(out_sel[2]), 
	.A2(I2[20]), 
	.B1(out_sel[3]), 
	.B2(I3[20]), 
	.Z(O1[20])); 
	AO_CELL inst_2_20 ( 
	.A1(out_sel[4]), 
	.A2(I4[20]), 
	.B1(out_sel[5]), 
	.B2(I5[20]), 
	.Z(O2[20])); 
	AO_CELL inst_3_20 ( 
	.A1(out_sel[6]), 
	.A2(I6[20]), 
	.B1(out_sel[7]), 
	.B2(I7[20]), 
	.Z(O3[20])); 
	AO_CELL inst_4_20 ( 
	.A1(out_sel[8]), 
	.A2(I8[20]), 
	.B1(out_sel[9]), 
	.B2(I9[20]), 
	.Z(O4[20])); 
	AO_CELL inst_5_20 ( 
	.A1(out_sel[10]), 
	.A2(I10[20]), 
	.B1(out_sel[11]), 
	.B2(I11[20]), 
	.Z(O5[20])); 
	AO_CELL inst_6_20 ( 
	.A1(out_sel[12]), 
	.A2(I12[20]), 
	.B1(out_sel[13]), 
	.B2(I13[20]), 
	.Z(O6[20])); 
	AO_CELL inst_7_20 ( 
	.A1(out_sel[14]), 
	.A2(I14[20]), 
	.B1(out_sel[15]), 
	.B2(I15[20]), 
	.Z(O7[20])); 
	AO_CELL inst_0_21 ( 
	.A1(out_sel[0]), 
	.A2(I0[21]), 
	.B1(out_sel[1]), 
	.B2(I1[21]), 
	.Z(O0[21])); 
	AO_CELL inst_1_21 ( 
	.A1(out_sel[2]), 
	.A2(I2[21]), 
	.B1(out_sel[3]), 
	.B2(I3[21]), 
	.Z(O1[21])); 
	AO_CELL inst_2_21 ( 
	.A1(out_sel[4]), 
	.A2(I4[21]), 
	.B1(out_sel[5]), 
	.B2(I5[21]), 
	.Z(O2[21])); 
	AO_CELL inst_3_21 ( 
	.A1(out_sel[6]), 
	.A2(I6[21]), 
	.B1(out_sel[7]), 
	.B2(I7[21]), 
	.Z(O3[21])); 
	AO_CELL inst_4_21 ( 
	.A1(out_sel[8]), 
	.A2(I8[21]), 
	.B1(out_sel[9]), 
	.B2(I9[21]), 
	.Z(O4[21])); 
	AO_CELL inst_5_21 ( 
	.A1(out_sel[10]), 
	.A2(I10[21]), 
	.B1(out_sel[11]), 
	.B2(I11[21]), 
	.Z(O5[21])); 
	AO_CELL inst_6_21 ( 
	.A1(out_sel[12]), 
	.A2(I12[21]), 
	.B1(out_sel[13]), 
	.B2(I13[21]), 
	.Z(O6[21])); 
	AO_CELL inst_7_21 ( 
	.A1(out_sel[14]), 
	.A2(I14[21]), 
	.B1(out_sel[15]), 
	.B2(I15[21]), 
	.Z(O7[21])); 
	AO_CELL inst_0_22 ( 
	.A1(out_sel[0]), 
	.A2(I0[22]), 
	.B1(out_sel[1]), 
	.B2(I1[22]), 
	.Z(O0[22])); 
	AO_CELL inst_1_22 ( 
	.A1(out_sel[2]), 
	.A2(I2[22]), 
	.B1(out_sel[3]), 
	.B2(I3[22]), 
	.Z(O1[22])); 
	AO_CELL inst_2_22 ( 
	.A1(out_sel[4]), 
	.A2(I4[22]), 
	.B1(out_sel[5]), 
	.B2(I5[22]), 
	.Z(O2[22])); 
	AO_CELL inst_3_22 ( 
	.A1(out_sel[6]), 
	.A2(I6[22]), 
	.B1(out_sel[7]), 
	.B2(I7[22]), 
	.Z(O3[22])); 
	AO_CELL inst_4_22 ( 
	.A1(out_sel[8]), 
	.A2(I8[22]), 
	.B1(out_sel[9]), 
	.B2(I9[22]), 
	.Z(O4[22])); 
	AO_CELL inst_5_22 ( 
	.A1(out_sel[10]), 
	.A2(I10[22]), 
	.B1(out_sel[11]), 
	.B2(I11[22]), 
	.Z(O5[22])); 
	AO_CELL inst_6_22 ( 
	.A1(out_sel[12]), 
	.A2(I12[22]), 
	.B1(out_sel[13]), 
	.B2(I13[22]), 
	.Z(O6[22])); 
	AO_CELL inst_7_22 ( 
	.A1(out_sel[14]), 
	.A2(I14[22]), 
	.B1(out_sel[15]), 
	.B2(I15[22]), 
	.Z(O7[22])); 
	AO_CELL inst_0_23 ( 
	.A1(out_sel[0]), 
	.A2(I0[23]), 
	.B1(out_sel[1]), 
	.B2(I1[23]), 
	.Z(O0[23])); 
	AO_CELL inst_1_23 ( 
	.A1(out_sel[2]), 
	.A2(I2[23]), 
	.B1(out_sel[3]), 
	.B2(I3[23]), 
	.Z(O1[23])); 
	AO_CELL inst_2_23 ( 
	.A1(out_sel[4]), 
	.A2(I4[23]), 
	.B1(out_sel[5]), 
	.B2(I5[23]), 
	.Z(O2[23])); 
	AO_CELL inst_3_23 ( 
	.A1(out_sel[6]), 
	.A2(I6[23]), 
	.B1(out_sel[7]), 
	.B2(I7[23]), 
	.Z(O3[23])); 
	AO_CELL inst_4_23 ( 
	.A1(out_sel[8]), 
	.A2(I8[23]), 
	.B1(out_sel[9]), 
	.B2(I9[23]), 
	.Z(O4[23])); 
	AO_CELL inst_5_23 ( 
	.A1(out_sel[10]), 
	.A2(I10[23]), 
	.B1(out_sel[11]), 
	.B2(I11[23]), 
	.Z(O5[23])); 
	AO_CELL inst_6_23 ( 
	.A1(out_sel[12]), 
	.A2(I12[23]), 
	.B1(out_sel[13]), 
	.B2(I13[23]), 
	.Z(O6[23])); 
	AO_CELL inst_7_23 ( 
	.A1(out_sel[14]), 
	.A2(I14[23]), 
	.B1(out_sel[15]), 
	.B2(I15[23]), 
	.Z(O7[23])); 
	AO_CELL inst_0_24 ( 
	.A1(out_sel[0]), 
	.A2(I0[24]), 
	.B1(out_sel[1]), 
	.B2(I1[24]), 
	.Z(O0[24])); 
	AO_CELL inst_1_24 ( 
	.A1(out_sel[2]), 
	.A2(I2[24]), 
	.B1(out_sel[3]), 
	.B2(I3[24]), 
	.Z(O1[24])); 
	AO_CELL inst_2_24 ( 
	.A1(out_sel[4]), 
	.A2(I4[24]), 
	.B1(out_sel[5]), 
	.B2(I5[24]), 
	.Z(O2[24])); 
	AO_CELL inst_3_24 ( 
	.A1(out_sel[6]), 
	.A2(I6[24]), 
	.B1(out_sel[7]), 
	.B2(I7[24]), 
	.Z(O3[24])); 
	AO_CELL inst_4_24 ( 
	.A1(out_sel[8]), 
	.A2(I8[24]), 
	.B1(out_sel[9]), 
	.B2(I9[24]), 
	.Z(O4[24])); 
	AO_CELL inst_5_24 ( 
	.A1(out_sel[10]), 
	.A2(I10[24]), 
	.B1(out_sel[11]), 
	.B2(I11[24]), 
	.Z(O5[24])); 
	AO_CELL inst_6_24 ( 
	.A1(out_sel[12]), 
	.A2(I12[24]), 
	.B1(out_sel[13]), 
	.B2(I13[24]), 
	.Z(O6[24])); 
	AO_CELL inst_7_24 ( 
	.A1(out_sel[14]), 
	.A2(I14[24]), 
	.B1(out_sel[15]), 
	.B2(I15[24]), 
	.Z(O7[24])); 
	AO_CELL inst_0_25 ( 
	.A1(out_sel[0]), 
	.A2(I0[25]), 
	.B1(out_sel[1]), 
	.B2(I1[25]), 
	.Z(O0[25])); 
	AO_CELL inst_1_25 ( 
	.A1(out_sel[2]), 
	.A2(I2[25]), 
	.B1(out_sel[3]), 
	.B2(I3[25]), 
	.Z(O1[25])); 
	AO_CELL inst_2_25 ( 
	.A1(out_sel[4]), 
	.A2(I4[25]), 
	.B1(out_sel[5]), 
	.B2(I5[25]), 
	.Z(O2[25])); 
	AO_CELL inst_3_25 ( 
	.A1(out_sel[6]), 
	.A2(I6[25]), 
	.B1(out_sel[7]), 
	.B2(I7[25]), 
	.Z(O3[25])); 
	AO_CELL inst_4_25 ( 
	.A1(out_sel[8]), 
	.A2(I8[25]), 
	.B1(out_sel[9]), 
	.B2(I9[25]), 
	.Z(O4[25])); 
	AO_CELL inst_5_25 ( 
	.A1(out_sel[10]), 
	.A2(I10[25]), 
	.B1(out_sel[11]), 
	.B2(I11[25]), 
	.Z(O5[25])); 
	AO_CELL inst_6_25 ( 
	.A1(out_sel[12]), 
	.A2(I12[25]), 
	.B1(out_sel[13]), 
	.B2(I13[25]), 
	.Z(O6[25])); 
	AO_CELL inst_7_25 ( 
	.A1(out_sel[14]), 
	.A2(I14[25]), 
	.B1(out_sel[15]), 
	.B2(I15[25]), 
	.Z(O7[25])); 
	AO_CELL inst_0_26 ( 
	.A1(out_sel[0]), 
	.A2(I0[26]), 
	.B1(out_sel[1]), 
	.B2(I1[26]), 
	.Z(O0[26])); 
	AO_CELL inst_1_26 ( 
	.A1(out_sel[2]), 
	.A2(I2[26]), 
	.B1(out_sel[3]), 
	.B2(I3[26]), 
	.Z(O1[26])); 
	AO_CELL inst_2_26 ( 
	.A1(out_sel[4]), 
	.A2(I4[26]), 
	.B1(out_sel[5]), 
	.B2(I5[26]), 
	.Z(O2[26])); 
	AO_CELL inst_3_26 ( 
	.A1(out_sel[6]), 
	.A2(I6[26]), 
	.B1(out_sel[7]), 
	.B2(I7[26]), 
	.Z(O3[26])); 
	AO_CELL inst_4_26 ( 
	.A1(out_sel[8]), 
	.A2(I8[26]), 
	.B1(out_sel[9]), 
	.B2(I9[26]), 
	.Z(O4[26])); 
	AO_CELL inst_5_26 ( 
	.A1(out_sel[10]), 
	.A2(I10[26]), 
	.B1(out_sel[11]), 
	.B2(I11[26]), 
	.Z(O5[26])); 
	AO_CELL inst_6_26 ( 
	.A1(out_sel[12]), 
	.A2(I12[26]), 
	.B1(out_sel[13]), 
	.B2(I13[26]), 
	.Z(O6[26])); 
	AO_CELL inst_7_26 ( 
	.A1(out_sel[14]), 
	.A2(I14[26]), 
	.B1(out_sel[15]), 
	.B2(I15[26]), 
	.Z(O7[26])); 
	AO_CELL inst_0_27 ( 
	.A1(out_sel[0]), 
	.A2(I0[27]), 
	.B1(out_sel[1]), 
	.B2(I1[27]), 
	.Z(O0[27])); 
	AO_CELL inst_1_27 ( 
	.A1(out_sel[2]), 
	.A2(I2[27]), 
	.B1(out_sel[3]), 
	.B2(I3[27]), 
	.Z(O1[27])); 
	AO_CELL inst_2_27 ( 
	.A1(out_sel[4]), 
	.A2(I4[27]), 
	.B1(out_sel[5]), 
	.B2(I5[27]), 
	.Z(O2[27])); 
	AO_CELL inst_3_27 ( 
	.A1(out_sel[6]), 
	.A2(I6[27]), 
	.B1(out_sel[7]), 
	.B2(I7[27]), 
	.Z(O3[27])); 
	AO_CELL inst_4_27 ( 
	.A1(out_sel[8]), 
	.A2(I8[27]), 
	.B1(out_sel[9]), 
	.B2(I9[27]), 
	.Z(O4[27])); 
	AO_CELL inst_5_27 ( 
	.A1(out_sel[10]), 
	.A2(I10[27]), 
	.B1(out_sel[11]), 
	.B2(I11[27]), 
	.Z(O5[27])); 
	AO_CELL inst_6_27 ( 
	.A1(out_sel[12]), 
	.A2(I12[27]), 
	.B1(out_sel[13]), 
	.B2(I13[27]), 
	.Z(O6[27])); 
	AO_CELL inst_7_27 ( 
	.A1(out_sel[14]), 
	.A2(I14[27]), 
	.B1(out_sel[15]), 
	.B2(I15[27]), 
	.Z(O7[27])); 
	AO_CELL inst_0_28 ( 
	.A1(out_sel[0]), 
	.A2(I0[28]), 
	.B1(out_sel[1]), 
	.B2(I1[28]), 
	.Z(O0[28])); 
	AO_CELL inst_1_28 ( 
	.A1(out_sel[2]), 
	.A2(I2[28]), 
	.B1(out_sel[3]), 
	.B2(I3[28]), 
	.Z(O1[28])); 
	AO_CELL inst_2_28 ( 
	.A1(out_sel[4]), 
	.A2(I4[28]), 
	.B1(out_sel[5]), 
	.B2(I5[28]), 
	.Z(O2[28])); 
	AO_CELL inst_3_28 ( 
	.A1(out_sel[6]), 
	.A2(I6[28]), 
	.B1(out_sel[7]), 
	.B2(I7[28]), 
	.Z(O3[28])); 
	AO_CELL inst_4_28 ( 
	.A1(out_sel[8]), 
	.A2(I8[28]), 
	.B1(out_sel[9]), 
	.B2(I9[28]), 
	.Z(O4[28])); 
	AO_CELL inst_5_28 ( 
	.A1(out_sel[10]), 
	.A2(I10[28]), 
	.B1(out_sel[11]), 
	.B2(I11[28]), 
	.Z(O5[28])); 
	AO_CELL inst_6_28 ( 
	.A1(out_sel[12]), 
	.A2(I12[28]), 
	.B1(out_sel[13]), 
	.B2(I13[28]), 
	.Z(O6[28])); 
	AO_CELL inst_7_28 ( 
	.A1(out_sel[14]), 
	.A2(I14[28]), 
	.B1(out_sel[15]), 
	.B2(I15[28]), 
	.Z(O7[28])); 
	AO_CELL inst_0_29 ( 
	.A1(out_sel[0]), 
	.A2(I0[29]), 
	.B1(out_sel[1]), 
	.B2(I1[29]), 
	.Z(O0[29])); 
	AO_CELL inst_1_29 ( 
	.A1(out_sel[2]), 
	.A2(I2[29]), 
	.B1(out_sel[3]), 
	.B2(I3[29]), 
	.Z(O1[29])); 
	AO_CELL inst_2_29 ( 
	.A1(out_sel[4]), 
	.A2(I4[29]), 
	.B1(out_sel[5]), 
	.B2(I5[29]), 
	.Z(O2[29])); 
	AO_CELL inst_3_29 ( 
	.A1(out_sel[6]), 
	.A2(I6[29]), 
	.B1(out_sel[7]), 
	.B2(I7[29]), 
	.Z(O3[29])); 
	AO_CELL inst_4_29 ( 
	.A1(out_sel[8]), 
	.A2(I8[29]), 
	.B1(out_sel[9]), 
	.B2(I9[29]), 
	.Z(O4[29])); 
	AO_CELL inst_5_29 ( 
	.A1(out_sel[10]), 
	.A2(I10[29]), 
	.B1(out_sel[11]), 
	.B2(I11[29]), 
	.Z(O5[29])); 
	AO_CELL inst_6_29 ( 
	.A1(out_sel[12]), 
	.A2(I12[29]), 
	.B1(out_sel[13]), 
	.B2(I13[29]), 
	.Z(O6[29])); 
	AO_CELL inst_7_29 ( 
	.A1(out_sel[14]), 
	.A2(I14[29]), 
	.B1(out_sel[15]), 
	.B2(I15[29]), 
	.Z(O7[29])); 
	AO_CELL inst_0_30 ( 
	.A1(out_sel[0]), 
	.A2(I0[30]), 
	.B1(out_sel[1]), 
	.B2(I1[30]), 
	.Z(O0[30])); 
	AO_CELL inst_1_30 ( 
	.A1(out_sel[2]), 
	.A2(I2[30]), 
	.B1(out_sel[3]), 
	.B2(I3[30]), 
	.Z(O1[30])); 
	AO_CELL inst_2_30 ( 
	.A1(out_sel[4]), 
	.A2(I4[30]), 
	.B1(out_sel[5]), 
	.B2(I5[30]), 
	.Z(O2[30])); 
	AO_CELL inst_3_30 ( 
	.A1(out_sel[6]), 
	.A2(I6[30]), 
	.B1(out_sel[7]), 
	.B2(I7[30]), 
	.Z(O3[30])); 
	AO_CELL inst_4_30 ( 
	.A1(out_sel[8]), 
	.A2(I8[30]), 
	.B1(out_sel[9]), 
	.B2(I9[30]), 
	.Z(O4[30])); 
	AO_CELL inst_5_30 ( 
	.A1(out_sel[10]), 
	.A2(I10[30]), 
	.B1(out_sel[11]), 
	.B2(I11[30]), 
	.Z(O5[30])); 
	AO_CELL inst_6_30 ( 
	.A1(out_sel[12]), 
	.A2(I12[30]), 
	.B1(out_sel[13]), 
	.B2(I13[30]), 
	.Z(O6[30])); 
	AO_CELL inst_7_30 ( 
	.A1(out_sel[14]), 
	.A2(I14[30]), 
	.B1(out_sel[15]), 
	.B2(I15[30]), 
	.Z(O7[30])); 
	AO_CELL inst_0_31 ( 
	.A1(out_sel[0]), 
	.A2(I0[31]), 
	.B1(out_sel[1]), 
	.B2(I1[31]), 
	.Z(O0[31])); 
	AO_CELL inst_1_31 ( 
	.A1(out_sel[2]), 
	.A2(I2[31]), 
	.B1(out_sel[3]), 
	.B2(I3[31]), 
	.Z(O1[31])); 
	AO_CELL inst_2_31 ( 
	.A1(out_sel[4]), 
	.A2(I4[31]), 
	.B1(out_sel[5]), 
	.B2(I5[31]), 
	.Z(O2[31])); 
	AO_CELL inst_3_31 ( 
	.A1(out_sel[6]), 
	.A2(I6[31]), 
	.B1(out_sel[7]), 
	.B2(I7[31]), 
	.Z(O3[31])); 
	AO_CELL inst_4_31 ( 
	.A1(out_sel[8]), 
	.A2(I8[31]), 
	.B1(out_sel[9]), 
	.B2(I9[31]), 
	.Z(O4[31])); 
	AO_CELL inst_5_31 ( 
	.A1(out_sel[10]), 
	.A2(I10[31]), 
	.B1(out_sel[11]), 
	.B2(I11[31]), 
	.Z(O5[31])); 
	AO_CELL inst_6_31 ( 
	.A1(out_sel[12]), 
	.A2(I12[31]), 
	.B1(out_sel[13]), 
	.B2(I13[31]), 
	.Z(O6[31])); 
	AO_CELL inst_7_31 ( 
	.A1(out_sel[14]), 
	.A2(I14[31]), 
	.B1(out_sel[15]), 
	.B2(I15[31]), 
	.Z(O7[31])); 
endmodule 

module mux_aoi_13_32 ( 
	input logic  [31 : 0] I[12:0], 
	input logic  [3 : 0] S ,
	output logic  [15 : 0] out_sel,
	output logic [31 : 0] O); 
	logic  [31 : 0] O_int0;
	logic  [31 : 0] O_int1;
	logic  [31 : 0] O_int2;
	logic  [31 : 0] O_int3;
	logic  [31 : 0] O_int4;
	logic  [31 : 0] O_int5;
	logic  [31 : 0] O_int6;

precoder_32_13 u_precoder ( 
	.S(S), 
	.out_sel(out_sel)); 

mux_logic_32_13 u_mux_logic ( 
	.I0 (I[0]),
	.I1 (I[1]),
	.I2 (I[2]),
	.I3 (I[3]),
	.I4 (I[4]),
	.I5 (I[5]),
	.I6 (I[6]),
	.I7 (I[7]),
	.I8 (I[8]),
	.I9 (I[9]),
	.I10 (I[10]),
	.I11 (I[11]),
	.I12 (I[12]),
	.out_sel(out_sel), 
	.O0(O_int0), 
	.O1(O_int1), 
	.O2(O_int2), 
	.O3(O_int3), 
	.O4(O_int4), 
	.O5(O_int5), 
	.O6(O_int6)); 
	assign O = (  	O_int0 | 	O_int1 | 	O_int2 | 	O_int3 | 	O_int4 | 	O_int5 | 	O_int6 	); 

endmodule 

module precoder_32_13 (
	input logic  [3 : 0] S ,
	output logic  [15 : 0] out_sel );

always_comb begin: mux_sel
	case (S) 
		4'd0    :   out_sel = 16'b0000000000000001;
		4'd1    :   out_sel = 16'b0000000000000010;
		4'd2    :   out_sel = 16'b0000000000000100;
		4'd3    :   out_sel = 16'b0000000000001000;
		4'd4    :   out_sel = 16'b0000000000010000;
		4'd5    :   out_sel = 16'b0000000000100000;
		4'd6    :   out_sel = 16'b0000000001000000;
		4'd7    :   out_sel = 16'b0000000010000000;
		4'd8    :   out_sel = 16'b0000000100000000;
		4'd9    :   out_sel = 16'b0000001000000000;
		4'd10    :   out_sel = 16'b0000010000000000;
		4'd11    :   out_sel = 16'b0000100000000000;
		4'd12    :   out_sel = 16'b0001000000000000;
		default :   out_sel = 16'b0;
	endcase 
end 

endmodule 

module mux_logic_32_13 ( 
	input logic  [15 : 0] out_sel,
	input logic  [31 : 0] I0, 
	input logic  [31 : 0] I1, 
	input logic  [31 : 0] I2, 
	input logic  [31 : 0] I3, 
	input logic  [31 : 0] I4, 
	input logic  [31 : 0] I5, 
	input logic  [31 : 0] I6, 
	input logic  [31 : 0] I7, 
	input logic  [31 : 0] I8, 
	input logic  [31 : 0] I9, 
	input logic  [31 : 0] I10, 
	input logic  [31 : 0] I11, 
	input logic  [31 : 0] I12, 
	output logic  [31 : 0] O0, 
	output logic  [31 : 0] O1, 
	output logic  [31 : 0] O2, 
	output logic  [31 : 0] O3, 
	output logic  [31 : 0] O4, 
	output logic  [31 : 0] O5, 
	output logic  [31 : 0] O6); 
	AO_CELL inst_0_0 ( 
	.A1(out_sel[0]), 
	.A2(I0[0]), 
	.B1(out_sel[1]), 
	.B2(I1[0]), 
	.Z(O0[0])); 
	AO_CELL inst_1_0 ( 
	.A1(out_sel[2]), 
	.A2(I2[0]), 
	.B1(out_sel[3]), 
	.B2(I3[0]), 
	.Z(O1[0])); 
	AO_CELL inst_2_0 ( 
	.A1(out_sel[4]), 
	.A2(I4[0]), 
	.B1(out_sel[5]), 
	.B2(I5[0]), 
	.Z(O2[0])); 
	AO_CELL inst_3_0 ( 
	.A1(out_sel[6]), 
	.A2(I6[0]), 
	.B1(out_sel[7]), 
	.B2(I7[0]), 
	.Z(O3[0])); 
	AO_CELL inst_4_0 ( 
	.A1(out_sel[8]), 
	.A2(I8[0]), 
	.B1(out_sel[9]), 
	.B2(I9[0]), 
	.Z(O4[0])); 
	AO_CELL inst_5_0 ( 
	.A1(out_sel[10]), 
	.A2(I10[0]), 
	.B1(out_sel[11]), 
	.B2(I11[0]), 
	.Z(O5[0])); 
	AN_CELL inst_and_0 ( 
	.A1(out_sel[12]), 
	.A2(I12[0]), 
	.Z(O6[0])); 
	AO_CELL inst_0_1 ( 
	.A1(out_sel[0]), 
	.A2(I0[1]), 
	.B1(out_sel[1]), 
	.B2(I1[1]), 
	.Z(O0[1])); 
	AO_CELL inst_1_1 ( 
	.A1(out_sel[2]), 
	.A2(I2[1]), 
	.B1(out_sel[3]), 
	.B2(I3[1]), 
	.Z(O1[1])); 
	AO_CELL inst_2_1 ( 
	.A1(out_sel[4]), 
	.A2(I4[1]), 
	.B1(out_sel[5]), 
	.B2(I5[1]), 
	.Z(O2[1])); 
	AO_CELL inst_3_1 ( 
	.A1(out_sel[6]), 
	.A2(I6[1]), 
	.B1(out_sel[7]), 
	.B2(I7[1]), 
	.Z(O3[1])); 
	AO_CELL inst_4_1 ( 
	.A1(out_sel[8]), 
	.A2(I8[1]), 
	.B1(out_sel[9]), 
	.B2(I9[1]), 
	.Z(O4[1])); 
	AO_CELL inst_5_1 ( 
	.A1(out_sel[10]), 
	.A2(I10[1]), 
	.B1(out_sel[11]), 
	.B2(I11[1]), 
	.Z(O5[1])); 
	AN_CELL inst_and_1 ( 
	.A1(out_sel[12]), 
	.A2(I12[1]), 
	.Z(O6[1])); 
	AO_CELL inst_0_2 ( 
	.A1(out_sel[0]), 
	.A2(I0[2]), 
	.B1(out_sel[1]), 
	.B2(I1[2]), 
	.Z(O0[2])); 
	AO_CELL inst_1_2 ( 
	.A1(out_sel[2]), 
	.A2(I2[2]), 
	.B1(out_sel[3]), 
	.B2(I3[2]), 
	.Z(O1[2])); 
	AO_CELL inst_2_2 ( 
	.A1(out_sel[4]), 
	.A2(I4[2]), 
	.B1(out_sel[5]), 
	.B2(I5[2]), 
	.Z(O2[2])); 
	AO_CELL inst_3_2 ( 
	.A1(out_sel[6]), 
	.A2(I6[2]), 
	.B1(out_sel[7]), 
	.B2(I7[2]), 
	.Z(O3[2])); 
	AO_CELL inst_4_2 ( 
	.A1(out_sel[8]), 
	.A2(I8[2]), 
	.B1(out_sel[9]), 
	.B2(I9[2]), 
	.Z(O4[2])); 
	AO_CELL inst_5_2 ( 
	.A1(out_sel[10]), 
	.A2(I10[2]), 
	.B1(out_sel[11]), 
	.B2(I11[2]), 
	.Z(O5[2])); 
	AN_CELL inst_and_2 ( 
	.A1(out_sel[12]), 
	.A2(I12[2]), 
	.Z(O6[2])); 
	AO_CELL inst_0_3 ( 
	.A1(out_sel[0]), 
	.A2(I0[3]), 
	.B1(out_sel[1]), 
	.B2(I1[3]), 
	.Z(O0[3])); 
	AO_CELL inst_1_3 ( 
	.A1(out_sel[2]), 
	.A2(I2[3]), 
	.B1(out_sel[3]), 
	.B2(I3[3]), 
	.Z(O1[3])); 
	AO_CELL inst_2_3 ( 
	.A1(out_sel[4]), 
	.A2(I4[3]), 
	.B1(out_sel[5]), 
	.B2(I5[3]), 
	.Z(O2[3])); 
	AO_CELL inst_3_3 ( 
	.A1(out_sel[6]), 
	.A2(I6[3]), 
	.B1(out_sel[7]), 
	.B2(I7[3]), 
	.Z(O3[3])); 
	AO_CELL inst_4_3 ( 
	.A1(out_sel[8]), 
	.A2(I8[3]), 
	.B1(out_sel[9]), 
	.B2(I9[3]), 
	.Z(O4[3])); 
	AO_CELL inst_5_3 ( 
	.A1(out_sel[10]), 
	.A2(I10[3]), 
	.B1(out_sel[11]), 
	.B2(I11[3]), 
	.Z(O5[3])); 
	AN_CELL inst_and_3 ( 
	.A1(out_sel[12]), 
	.A2(I12[3]), 
	.Z(O6[3])); 
	AO_CELL inst_0_4 ( 
	.A1(out_sel[0]), 
	.A2(I0[4]), 
	.B1(out_sel[1]), 
	.B2(I1[4]), 
	.Z(O0[4])); 
	AO_CELL inst_1_4 ( 
	.A1(out_sel[2]), 
	.A2(I2[4]), 
	.B1(out_sel[3]), 
	.B2(I3[4]), 
	.Z(O1[4])); 
	AO_CELL inst_2_4 ( 
	.A1(out_sel[4]), 
	.A2(I4[4]), 
	.B1(out_sel[5]), 
	.B2(I5[4]), 
	.Z(O2[4])); 
	AO_CELL inst_3_4 ( 
	.A1(out_sel[6]), 
	.A2(I6[4]), 
	.B1(out_sel[7]), 
	.B2(I7[4]), 
	.Z(O3[4])); 
	AO_CELL inst_4_4 ( 
	.A1(out_sel[8]), 
	.A2(I8[4]), 
	.B1(out_sel[9]), 
	.B2(I9[4]), 
	.Z(O4[4])); 
	AO_CELL inst_5_4 ( 
	.A1(out_sel[10]), 
	.A2(I10[4]), 
	.B1(out_sel[11]), 
	.B2(I11[4]), 
	.Z(O5[4])); 
	AN_CELL inst_and_4 ( 
	.A1(out_sel[12]), 
	.A2(I12[4]), 
	.Z(O6[4])); 
	AO_CELL inst_0_5 ( 
	.A1(out_sel[0]), 
	.A2(I0[5]), 
	.B1(out_sel[1]), 
	.B2(I1[5]), 
	.Z(O0[5])); 
	AO_CELL inst_1_5 ( 
	.A1(out_sel[2]), 
	.A2(I2[5]), 
	.B1(out_sel[3]), 
	.B2(I3[5]), 
	.Z(O1[5])); 
	AO_CELL inst_2_5 ( 
	.A1(out_sel[4]), 
	.A2(I4[5]), 
	.B1(out_sel[5]), 
	.B2(I5[5]), 
	.Z(O2[5])); 
	AO_CELL inst_3_5 ( 
	.A1(out_sel[6]), 
	.A2(I6[5]), 
	.B1(out_sel[7]), 
	.B2(I7[5]), 
	.Z(O3[5])); 
	AO_CELL inst_4_5 ( 
	.A1(out_sel[8]), 
	.A2(I8[5]), 
	.B1(out_sel[9]), 
	.B2(I9[5]), 
	.Z(O4[5])); 
	AO_CELL inst_5_5 ( 
	.A1(out_sel[10]), 
	.A2(I10[5]), 
	.B1(out_sel[11]), 
	.B2(I11[5]), 
	.Z(O5[5])); 
	AN_CELL inst_and_5 ( 
	.A1(out_sel[12]), 
	.A2(I12[5]), 
	.Z(O6[5])); 
	AO_CELL inst_0_6 ( 
	.A1(out_sel[0]), 
	.A2(I0[6]), 
	.B1(out_sel[1]), 
	.B2(I1[6]), 
	.Z(O0[6])); 
	AO_CELL inst_1_6 ( 
	.A1(out_sel[2]), 
	.A2(I2[6]), 
	.B1(out_sel[3]), 
	.B2(I3[6]), 
	.Z(O1[6])); 
	AO_CELL inst_2_6 ( 
	.A1(out_sel[4]), 
	.A2(I4[6]), 
	.B1(out_sel[5]), 
	.B2(I5[6]), 
	.Z(O2[6])); 
	AO_CELL inst_3_6 ( 
	.A1(out_sel[6]), 
	.A2(I6[6]), 
	.B1(out_sel[7]), 
	.B2(I7[6]), 
	.Z(O3[6])); 
	AO_CELL inst_4_6 ( 
	.A1(out_sel[8]), 
	.A2(I8[6]), 
	.B1(out_sel[9]), 
	.B2(I9[6]), 
	.Z(O4[6])); 
	AO_CELL inst_5_6 ( 
	.A1(out_sel[10]), 
	.A2(I10[6]), 
	.B1(out_sel[11]), 
	.B2(I11[6]), 
	.Z(O5[6])); 
	AN_CELL inst_and_6 ( 
	.A1(out_sel[12]), 
	.A2(I12[6]), 
	.Z(O6[6])); 
	AO_CELL inst_0_7 ( 
	.A1(out_sel[0]), 
	.A2(I0[7]), 
	.B1(out_sel[1]), 
	.B2(I1[7]), 
	.Z(O0[7])); 
	AO_CELL inst_1_7 ( 
	.A1(out_sel[2]), 
	.A2(I2[7]), 
	.B1(out_sel[3]), 
	.B2(I3[7]), 
	.Z(O1[7])); 
	AO_CELL inst_2_7 ( 
	.A1(out_sel[4]), 
	.A2(I4[7]), 
	.B1(out_sel[5]), 
	.B2(I5[7]), 
	.Z(O2[7])); 
	AO_CELL inst_3_7 ( 
	.A1(out_sel[6]), 
	.A2(I6[7]), 
	.B1(out_sel[7]), 
	.B2(I7[7]), 
	.Z(O3[7])); 
	AO_CELL inst_4_7 ( 
	.A1(out_sel[8]), 
	.A2(I8[7]), 
	.B1(out_sel[9]), 
	.B2(I9[7]), 
	.Z(O4[7])); 
	AO_CELL inst_5_7 ( 
	.A1(out_sel[10]), 
	.A2(I10[7]), 
	.B1(out_sel[11]), 
	.B2(I11[7]), 
	.Z(O5[7])); 
	AN_CELL inst_and_7 ( 
	.A1(out_sel[12]), 
	.A2(I12[7]), 
	.Z(O6[7])); 
	AO_CELL inst_0_8 ( 
	.A1(out_sel[0]), 
	.A2(I0[8]), 
	.B1(out_sel[1]), 
	.B2(I1[8]), 
	.Z(O0[8])); 
	AO_CELL inst_1_8 ( 
	.A1(out_sel[2]), 
	.A2(I2[8]), 
	.B1(out_sel[3]), 
	.B2(I3[8]), 
	.Z(O1[8])); 
	AO_CELL inst_2_8 ( 
	.A1(out_sel[4]), 
	.A2(I4[8]), 
	.B1(out_sel[5]), 
	.B2(I5[8]), 
	.Z(O2[8])); 
	AO_CELL inst_3_8 ( 
	.A1(out_sel[6]), 
	.A2(I6[8]), 
	.B1(out_sel[7]), 
	.B2(I7[8]), 
	.Z(O3[8])); 
	AO_CELL inst_4_8 ( 
	.A1(out_sel[8]), 
	.A2(I8[8]), 
	.B1(out_sel[9]), 
	.B2(I9[8]), 
	.Z(O4[8])); 
	AO_CELL inst_5_8 ( 
	.A1(out_sel[10]), 
	.A2(I10[8]), 
	.B1(out_sel[11]), 
	.B2(I11[8]), 
	.Z(O5[8])); 
	AN_CELL inst_and_8 ( 
	.A1(out_sel[12]), 
	.A2(I12[8]), 
	.Z(O6[8])); 
	AO_CELL inst_0_9 ( 
	.A1(out_sel[0]), 
	.A2(I0[9]), 
	.B1(out_sel[1]), 
	.B2(I1[9]), 
	.Z(O0[9])); 
	AO_CELL inst_1_9 ( 
	.A1(out_sel[2]), 
	.A2(I2[9]), 
	.B1(out_sel[3]), 
	.B2(I3[9]), 
	.Z(O1[9])); 
	AO_CELL inst_2_9 ( 
	.A1(out_sel[4]), 
	.A2(I4[9]), 
	.B1(out_sel[5]), 
	.B2(I5[9]), 
	.Z(O2[9])); 
	AO_CELL inst_3_9 ( 
	.A1(out_sel[6]), 
	.A2(I6[9]), 
	.B1(out_sel[7]), 
	.B2(I7[9]), 
	.Z(O3[9])); 
	AO_CELL inst_4_9 ( 
	.A1(out_sel[8]), 
	.A2(I8[9]), 
	.B1(out_sel[9]), 
	.B2(I9[9]), 
	.Z(O4[9])); 
	AO_CELL inst_5_9 ( 
	.A1(out_sel[10]), 
	.A2(I10[9]), 
	.B1(out_sel[11]), 
	.B2(I11[9]), 
	.Z(O5[9])); 
	AN_CELL inst_and_9 ( 
	.A1(out_sel[12]), 
	.A2(I12[9]), 
	.Z(O6[9])); 
	AO_CELL inst_0_10 ( 
	.A1(out_sel[0]), 
	.A2(I0[10]), 
	.B1(out_sel[1]), 
	.B2(I1[10]), 
	.Z(O0[10])); 
	AO_CELL inst_1_10 ( 
	.A1(out_sel[2]), 
	.A2(I2[10]), 
	.B1(out_sel[3]), 
	.B2(I3[10]), 
	.Z(O1[10])); 
	AO_CELL inst_2_10 ( 
	.A1(out_sel[4]), 
	.A2(I4[10]), 
	.B1(out_sel[5]), 
	.B2(I5[10]), 
	.Z(O2[10])); 
	AO_CELL inst_3_10 ( 
	.A1(out_sel[6]), 
	.A2(I6[10]), 
	.B1(out_sel[7]), 
	.B2(I7[10]), 
	.Z(O3[10])); 
	AO_CELL inst_4_10 ( 
	.A1(out_sel[8]), 
	.A2(I8[10]), 
	.B1(out_sel[9]), 
	.B2(I9[10]), 
	.Z(O4[10])); 
	AO_CELL inst_5_10 ( 
	.A1(out_sel[10]), 
	.A2(I10[10]), 
	.B1(out_sel[11]), 
	.B2(I11[10]), 
	.Z(O5[10])); 
	AN_CELL inst_and_10 ( 
	.A1(out_sel[12]), 
	.A2(I12[10]), 
	.Z(O6[10])); 
	AO_CELL inst_0_11 ( 
	.A1(out_sel[0]), 
	.A2(I0[11]), 
	.B1(out_sel[1]), 
	.B2(I1[11]), 
	.Z(O0[11])); 
	AO_CELL inst_1_11 ( 
	.A1(out_sel[2]), 
	.A2(I2[11]), 
	.B1(out_sel[3]), 
	.B2(I3[11]), 
	.Z(O1[11])); 
	AO_CELL inst_2_11 ( 
	.A1(out_sel[4]), 
	.A2(I4[11]), 
	.B1(out_sel[5]), 
	.B2(I5[11]), 
	.Z(O2[11])); 
	AO_CELL inst_3_11 ( 
	.A1(out_sel[6]), 
	.A2(I6[11]), 
	.B1(out_sel[7]), 
	.B2(I7[11]), 
	.Z(O3[11])); 
	AO_CELL inst_4_11 ( 
	.A1(out_sel[8]), 
	.A2(I8[11]), 
	.B1(out_sel[9]), 
	.B2(I9[11]), 
	.Z(O4[11])); 
	AO_CELL inst_5_11 ( 
	.A1(out_sel[10]), 
	.A2(I10[11]), 
	.B1(out_sel[11]), 
	.B2(I11[11]), 
	.Z(O5[11])); 
	AN_CELL inst_and_11 ( 
	.A1(out_sel[12]), 
	.A2(I12[11]), 
	.Z(O6[11])); 
	AO_CELL inst_0_12 ( 
	.A1(out_sel[0]), 
	.A2(I0[12]), 
	.B1(out_sel[1]), 
	.B2(I1[12]), 
	.Z(O0[12])); 
	AO_CELL inst_1_12 ( 
	.A1(out_sel[2]), 
	.A2(I2[12]), 
	.B1(out_sel[3]), 
	.B2(I3[12]), 
	.Z(O1[12])); 
	AO_CELL inst_2_12 ( 
	.A1(out_sel[4]), 
	.A2(I4[12]), 
	.B1(out_sel[5]), 
	.B2(I5[12]), 
	.Z(O2[12])); 
	AO_CELL inst_3_12 ( 
	.A1(out_sel[6]), 
	.A2(I6[12]), 
	.B1(out_sel[7]), 
	.B2(I7[12]), 
	.Z(O3[12])); 
	AO_CELL inst_4_12 ( 
	.A1(out_sel[8]), 
	.A2(I8[12]), 
	.B1(out_sel[9]), 
	.B2(I9[12]), 
	.Z(O4[12])); 
	AO_CELL inst_5_12 ( 
	.A1(out_sel[10]), 
	.A2(I10[12]), 
	.B1(out_sel[11]), 
	.B2(I11[12]), 
	.Z(O5[12])); 
	AN_CELL inst_and_12 ( 
	.A1(out_sel[12]), 
	.A2(I12[12]), 
	.Z(O6[12])); 
	AO_CELL inst_0_13 ( 
	.A1(out_sel[0]), 
	.A2(I0[13]), 
	.B1(out_sel[1]), 
	.B2(I1[13]), 
	.Z(O0[13])); 
	AO_CELL inst_1_13 ( 
	.A1(out_sel[2]), 
	.A2(I2[13]), 
	.B1(out_sel[3]), 
	.B2(I3[13]), 
	.Z(O1[13])); 
	AO_CELL inst_2_13 ( 
	.A1(out_sel[4]), 
	.A2(I4[13]), 
	.B1(out_sel[5]), 
	.B2(I5[13]), 
	.Z(O2[13])); 
	AO_CELL inst_3_13 ( 
	.A1(out_sel[6]), 
	.A2(I6[13]), 
	.B1(out_sel[7]), 
	.B2(I7[13]), 
	.Z(O3[13])); 
	AO_CELL inst_4_13 ( 
	.A1(out_sel[8]), 
	.A2(I8[13]), 
	.B1(out_sel[9]), 
	.B2(I9[13]), 
	.Z(O4[13])); 
	AO_CELL inst_5_13 ( 
	.A1(out_sel[10]), 
	.A2(I10[13]), 
	.B1(out_sel[11]), 
	.B2(I11[13]), 
	.Z(O5[13])); 
	AN_CELL inst_and_13 ( 
	.A1(out_sel[12]), 
	.A2(I12[13]), 
	.Z(O6[13])); 
	AO_CELL inst_0_14 ( 
	.A1(out_sel[0]), 
	.A2(I0[14]), 
	.B1(out_sel[1]), 
	.B2(I1[14]), 
	.Z(O0[14])); 
	AO_CELL inst_1_14 ( 
	.A1(out_sel[2]), 
	.A2(I2[14]), 
	.B1(out_sel[3]), 
	.B2(I3[14]), 
	.Z(O1[14])); 
	AO_CELL inst_2_14 ( 
	.A1(out_sel[4]), 
	.A2(I4[14]), 
	.B1(out_sel[5]), 
	.B2(I5[14]), 
	.Z(O2[14])); 
	AO_CELL inst_3_14 ( 
	.A1(out_sel[6]), 
	.A2(I6[14]), 
	.B1(out_sel[7]), 
	.B2(I7[14]), 
	.Z(O3[14])); 
	AO_CELL inst_4_14 ( 
	.A1(out_sel[8]), 
	.A2(I8[14]), 
	.B1(out_sel[9]), 
	.B2(I9[14]), 
	.Z(O4[14])); 
	AO_CELL inst_5_14 ( 
	.A1(out_sel[10]), 
	.A2(I10[14]), 
	.B1(out_sel[11]), 
	.B2(I11[14]), 
	.Z(O5[14])); 
	AN_CELL inst_and_14 ( 
	.A1(out_sel[12]), 
	.A2(I12[14]), 
	.Z(O6[14])); 
	AO_CELL inst_0_15 ( 
	.A1(out_sel[0]), 
	.A2(I0[15]), 
	.B1(out_sel[1]), 
	.B2(I1[15]), 
	.Z(O0[15])); 
	AO_CELL inst_1_15 ( 
	.A1(out_sel[2]), 
	.A2(I2[15]), 
	.B1(out_sel[3]), 
	.B2(I3[15]), 
	.Z(O1[15])); 
	AO_CELL inst_2_15 ( 
	.A1(out_sel[4]), 
	.A2(I4[15]), 
	.B1(out_sel[5]), 
	.B2(I5[15]), 
	.Z(O2[15])); 
	AO_CELL inst_3_15 ( 
	.A1(out_sel[6]), 
	.A2(I6[15]), 
	.B1(out_sel[7]), 
	.B2(I7[15]), 
	.Z(O3[15])); 
	AO_CELL inst_4_15 ( 
	.A1(out_sel[8]), 
	.A2(I8[15]), 
	.B1(out_sel[9]), 
	.B2(I9[15]), 
	.Z(O4[15])); 
	AO_CELL inst_5_15 ( 
	.A1(out_sel[10]), 
	.A2(I10[15]), 
	.B1(out_sel[11]), 
	.B2(I11[15]), 
	.Z(O5[15])); 
	AN_CELL inst_and_15 ( 
	.A1(out_sel[12]), 
	.A2(I12[15]), 
	.Z(O6[15])); 
	AO_CELL inst_0_16 ( 
	.A1(out_sel[0]), 
	.A2(I0[16]), 
	.B1(out_sel[1]), 
	.B2(I1[16]), 
	.Z(O0[16])); 
	AO_CELL inst_1_16 ( 
	.A1(out_sel[2]), 
	.A2(I2[16]), 
	.B1(out_sel[3]), 
	.B2(I3[16]), 
	.Z(O1[16])); 
	AO_CELL inst_2_16 ( 
	.A1(out_sel[4]), 
	.A2(I4[16]), 
	.B1(out_sel[5]), 
	.B2(I5[16]), 
	.Z(O2[16])); 
	AO_CELL inst_3_16 ( 
	.A1(out_sel[6]), 
	.A2(I6[16]), 
	.B1(out_sel[7]), 
	.B2(I7[16]), 
	.Z(O3[16])); 
	AO_CELL inst_4_16 ( 
	.A1(out_sel[8]), 
	.A2(I8[16]), 
	.B1(out_sel[9]), 
	.B2(I9[16]), 
	.Z(O4[16])); 
	AO_CELL inst_5_16 ( 
	.A1(out_sel[10]), 
	.A2(I10[16]), 
	.B1(out_sel[11]), 
	.B2(I11[16]), 
	.Z(O5[16])); 
	AN_CELL inst_and_16 ( 
	.A1(out_sel[12]), 
	.A2(I12[16]), 
	.Z(O6[16])); 
	AO_CELL inst_0_17 ( 
	.A1(out_sel[0]), 
	.A2(I0[17]), 
	.B1(out_sel[1]), 
	.B2(I1[17]), 
	.Z(O0[17])); 
	AO_CELL inst_1_17 ( 
	.A1(out_sel[2]), 
	.A2(I2[17]), 
	.B1(out_sel[3]), 
	.B2(I3[17]), 
	.Z(O1[17])); 
	AO_CELL inst_2_17 ( 
	.A1(out_sel[4]), 
	.A2(I4[17]), 
	.B1(out_sel[5]), 
	.B2(I5[17]), 
	.Z(O2[17])); 
	AO_CELL inst_3_17 ( 
	.A1(out_sel[6]), 
	.A2(I6[17]), 
	.B1(out_sel[7]), 
	.B2(I7[17]), 
	.Z(O3[17])); 
	AO_CELL inst_4_17 ( 
	.A1(out_sel[8]), 
	.A2(I8[17]), 
	.B1(out_sel[9]), 
	.B2(I9[17]), 
	.Z(O4[17])); 
	AO_CELL inst_5_17 ( 
	.A1(out_sel[10]), 
	.A2(I10[17]), 
	.B1(out_sel[11]), 
	.B2(I11[17]), 
	.Z(O5[17])); 
	AN_CELL inst_and_17 ( 
	.A1(out_sel[12]), 
	.A2(I12[17]), 
	.Z(O6[17])); 
	AO_CELL inst_0_18 ( 
	.A1(out_sel[0]), 
	.A2(I0[18]), 
	.B1(out_sel[1]), 
	.B2(I1[18]), 
	.Z(O0[18])); 
	AO_CELL inst_1_18 ( 
	.A1(out_sel[2]), 
	.A2(I2[18]), 
	.B1(out_sel[3]), 
	.B2(I3[18]), 
	.Z(O1[18])); 
	AO_CELL inst_2_18 ( 
	.A1(out_sel[4]), 
	.A2(I4[18]), 
	.B1(out_sel[5]), 
	.B2(I5[18]), 
	.Z(O2[18])); 
	AO_CELL inst_3_18 ( 
	.A1(out_sel[6]), 
	.A2(I6[18]), 
	.B1(out_sel[7]), 
	.B2(I7[18]), 
	.Z(O3[18])); 
	AO_CELL inst_4_18 ( 
	.A1(out_sel[8]), 
	.A2(I8[18]), 
	.B1(out_sel[9]), 
	.B2(I9[18]), 
	.Z(O4[18])); 
	AO_CELL inst_5_18 ( 
	.A1(out_sel[10]), 
	.A2(I10[18]), 
	.B1(out_sel[11]), 
	.B2(I11[18]), 
	.Z(O5[18])); 
	AN_CELL inst_and_18 ( 
	.A1(out_sel[12]), 
	.A2(I12[18]), 
	.Z(O6[18])); 
	AO_CELL inst_0_19 ( 
	.A1(out_sel[0]), 
	.A2(I0[19]), 
	.B1(out_sel[1]), 
	.B2(I1[19]), 
	.Z(O0[19])); 
	AO_CELL inst_1_19 ( 
	.A1(out_sel[2]), 
	.A2(I2[19]), 
	.B1(out_sel[3]), 
	.B2(I3[19]), 
	.Z(O1[19])); 
	AO_CELL inst_2_19 ( 
	.A1(out_sel[4]), 
	.A2(I4[19]), 
	.B1(out_sel[5]), 
	.B2(I5[19]), 
	.Z(O2[19])); 
	AO_CELL inst_3_19 ( 
	.A1(out_sel[6]), 
	.A2(I6[19]), 
	.B1(out_sel[7]), 
	.B2(I7[19]), 
	.Z(O3[19])); 
	AO_CELL inst_4_19 ( 
	.A1(out_sel[8]), 
	.A2(I8[19]), 
	.B1(out_sel[9]), 
	.B2(I9[19]), 
	.Z(O4[19])); 
	AO_CELL inst_5_19 ( 
	.A1(out_sel[10]), 
	.A2(I10[19]), 
	.B1(out_sel[11]), 
	.B2(I11[19]), 
	.Z(O5[19])); 
	AN_CELL inst_and_19 ( 
	.A1(out_sel[12]), 
	.A2(I12[19]), 
	.Z(O6[19])); 
	AO_CELL inst_0_20 ( 
	.A1(out_sel[0]), 
	.A2(I0[20]), 
	.B1(out_sel[1]), 
	.B2(I1[20]), 
	.Z(O0[20])); 
	AO_CELL inst_1_20 ( 
	.A1(out_sel[2]), 
	.A2(I2[20]), 
	.B1(out_sel[3]), 
	.B2(I3[20]), 
	.Z(O1[20])); 
	AO_CELL inst_2_20 ( 
	.A1(out_sel[4]), 
	.A2(I4[20]), 
	.B1(out_sel[5]), 
	.B2(I5[20]), 
	.Z(O2[20])); 
	AO_CELL inst_3_20 ( 
	.A1(out_sel[6]), 
	.A2(I6[20]), 
	.B1(out_sel[7]), 
	.B2(I7[20]), 
	.Z(O3[20])); 
	AO_CELL inst_4_20 ( 
	.A1(out_sel[8]), 
	.A2(I8[20]), 
	.B1(out_sel[9]), 
	.B2(I9[20]), 
	.Z(O4[20])); 
	AO_CELL inst_5_20 ( 
	.A1(out_sel[10]), 
	.A2(I10[20]), 
	.B1(out_sel[11]), 
	.B2(I11[20]), 
	.Z(O5[20])); 
	AN_CELL inst_and_20 ( 
	.A1(out_sel[12]), 
	.A2(I12[20]), 
	.Z(O6[20])); 
	AO_CELL inst_0_21 ( 
	.A1(out_sel[0]), 
	.A2(I0[21]), 
	.B1(out_sel[1]), 
	.B2(I1[21]), 
	.Z(O0[21])); 
	AO_CELL inst_1_21 ( 
	.A1(out_sel[2]), 
	.A2(I2[21]), 
	.B1(out_sel[3]), 
	.B2(I3[21]), 
	.Z(O1[21])); 
	AO_CELL inst_2_21 ( 
	.A1(out_sel[4]), 
	.A2(I4[21]), 
	.B1(out_sel[5]), 
	.B2(I5[21]), 
	.Z(O2[21])); 
	AO_CELL inst_3_21 ( 
	.A1(out_sel[6]), 
	.A2(I6[21]), 
	.B1(out_sel[7]), 
	.B2(I7[21]), 
	.Z(O3[21])); 
	AO_CELL inst_4_21 ( 
	.A1(out_sel[8]), 
	.A2(I8[21]), 
	.B1(out_sel[9]), 
	.B2(I9[21]), 
	.Z(O4[21])); 
	AO_CELL inst_5_21 ( 
	.A1(out_sel[10]), 
	.A2(I10[21]), 
	.B1(out_sel[11]), 
	.B2(I11[21]), 
	.Z(O5[21])); 
	AN_CELL inst_and_21 ( 
	.A1(out_sel[12]), 
	.A2(I12[21]), 
	.Z(O6[21])); 
	AO_CELL inst_0_22 ( 
	.A1(out_sel[0]), 
	.A2(I0[22]), 
	.B1(out_sel[1]), 
	.B2(I1[22]), 
	.Z(O0[22])); 
	AO_CELL inst_1_22 ( 
	.A1(out_sel[2]), 
	.A2(I2[22]), 
	.B1(out_sel[3]), 
	.B2(I3[22]), 
	.Z(O1[22])); 
	AO_CELL inst_2_22 ( 
	.A1(out_sel[4]), 
	.A2(I4[22]), 
	.B1(out_sel[5]), 
	.B2(I5[22]), 
	.Z(O2[22])); 
	AO_CELL inst_3_22 ( 
	.A1(out_sel[6]), 
	.A2(I6[22]), 
	.B1(out_sel[7]), 
	.B2(I7[22]), 
	.Z(O3[22])); 
	AO_CELL inst_4_22 ( 
	.A1(out_sel[8]), 
	.A2(I8[22]), 
	.B1(out_sel[9]), 
	.B2(I9[22]), 
	.Z(O4[22])); 
	AO_CELL inst_5_22 ( 
	.A1(out_sel[10]), 
	.A2(I10[22]), 
	.B1(out_sel[11]), 
	.B2(I11[22]), 
	.Z(O5[22])); 
	AN_CELL inst_and_22 ( 
	.A1(out_sel[12]), 
	.A2(I12[22]), 
	.Z(O6[22])); 
	AO_CELL inst_0_23 ( 
	.A1(out_sel[0]), 
	.A2(I0[23]), 
	.B1(out_sel[1]), 
	.B2(I1[23]), 
	.Z(O0[23])); 
	AO_CELL inst_1_23 ( 
	.A1(out_sel[2]), 
	.A2(I2[23]), 
	.B1(out_sel[3]), 
	.B2(I3[23]), 
	.Z(O1[23])); 
	AO_CELL inst_2_23 ( 
	.A1(out_sel[4]), 
	.A2(I4[23]), 
	.B1(out_sel[5]), 
	.B2(I5[23]), 
	.Z(O2[23])); 
	AO_CELL inst_3_23 ( 
	.A1(out_sel[6]), 
	.A2(I6[23]), 
	.B1(out_sel[7]), 
	.B2(I7[23]), 
	.Z(O3[23])); 
	AO_CELL inst_4_23 ( 
	.A1(out_sel[8]), 
	.A2(I8[23]), 
	.B1(out_sel[9]), 
	.B2(I9[23]), 
	.Z(O4[23])); 
	AO_CELL inst_5_23 ( 
	.A1(out_sel[10]), 
	.A2(I10[23]), 
	.B1(out_sel[11]), 
	.B2(I11[23]), 
	.Z(O5[23])); 
	AN_CELL inst_and_23 ( 
	.A1(out_sel[12]), 
	.A2(I12[23]), 
	.Z(O6[23])); 
	AO_CELL inst_0_24 ( 
	.A1(out_sel[0]), 
	.A2(I0[24]), 
	.B1(out_sel[1]), 
	.B2(I1[24]), 
	.Z(O0[24])); 
	AO_CELL inst_1_24 ( 
	.A1(out_sel[2]), 
	.A2(I2[24]), 
	.B1(out_sel[3]), 
	.B2(I3[24]), 
	.Z(O1[24])); 
	AO_CELL inst_2_24 ( 
	.A1(out_sel[4]), 
	.A2(I4[24]), 
	.B1(out_sel[5]), 
	.B2(I5[24]), 
	.Z(O2[24])); 
	AO_CELL inst_3_24 ( 
	.A1(out_sel[6]), 
	.A2(I6[24]), 
	.B1(out_sel[7]), 
	.B2(I7[24]), 
	.Z(O3[24])); 
	AO_CELL inst_4_24 ( 
	.A1(out_sel[8]), 
	.A2(I8[24]), 
	.B1(out_sel[9]), 
	.B2(I9[24]), 
	.Z(O4[24])); 
	AO_CELL inst_5_24 ( 
	.A1(out_sel[10]), 
	.A2(I10[24]), 
	.B1(out_sel[11]), 
	.B2(I11[24]), 
	.Z(O5[24])); 
	AN_CELL inst_and_24 ( 
	.A1(out_sel[12]), 
	.A2(I12[24]), 
	.Z(O6[24])); 
	AO_CELL inst_0_25 ( 
	.A1(out_sel[0]), 
	.A2(I0[25]), 
	.B1(out_sel[1]), 
	.B2(I1[25]), 
	.Z(O0[25])); 
	AO_CELL inst_1_25 ( 
	.A1(out_sel[2]), 
	.A2(I2[25]), 
	.B1(out_sel[3]), 
	.B2(I3[25]), 
	.Z(O1[25])); 
	AO_CELL inst_2_25 ( 
	.A1(out_sel[4]), 
	.A2(I4[25]), 
	.B1(out_sel[5]), 
	.B2(I5[25]), 
	.Z(O2[25])); 
	AO_CELL inst_3_25 ( 
	.A1(out_sel[6]), 
	.A2(I6[25]), 
	.B1(out_sel[7]), 
	.B2(I7[25]), 
	.Z(O3[25])); 
	AO_CELL inst_4_25 ( 
	.A1(out_sel[8]), 
	.A2(I8[25]), 
	.B1(out_sel[9]), 
	.B2(I9[25]), 
	.Z(O4[25])); 
	AO_CELL inst_5_25 ( 
	.A1(out_sel[10]), 
	.A2(I10[25]), 
	.B1(out_sel[11]), 
	.B2(I11[25]), 
	.Z(O5[25])); 
	AN_CELL inst_and_25 ( 
	.A1(out_sel[12]), 
	.A2(I12[25]), 
	.Z(O6[25])); 
	AO_CELL inst_0_26 ( 
	.A1(out_sel[0]), 
	.A2(I0[26]), 
	.B1(out_sel[1]), 
	.B2(I1[26]), 
	.Z(O0[26])); 
	AO_CELL inst_1_26 ( 
	.A1(out_sel[2]), 
	.A2(I2[26]), 
	.B1(out_sel[3]), 
	.B2(I3[26]), 
	.Z(O1[26])); 
	AO_CELL inst_2_26 ( 
	.A1(out_sel[4]), 
	.A2(I4[26]), 
	.B1(out_sel[5]), 
	.B2(I5[26]), 
	.Z(O2[26])); 
	AO_CELL inst_3_26 ( 
	.A1(out_sel[6]), 
	.A2(I6[26]), 
	.B1(out_sel[7]), 
	.B2(I7[26]), 
	.Z(O3[26])); 
	AO_CELL inst_4_26 ( 
	.A1(out_sel[8]), 
	.A2(I8[26]), 
	.B1(out_sel[9]), 
	.B2(I9[26]), 
	.Z(O4[26])); 
	AO_CELL inst_5_26 ( 
	.A1(out_sel[10]), 
	.A2(I10[26]), 
	.B1(out_sel[11]), 
	.B2(I11[26]), 
	.Z(O5[26])); 
	AN_CELL inst_and_26 ( 
	.A1(out_sel[12]), 
	.A2(I12[26]), 
	.Z(O6[26])); 
	AO_CELL inst_0_27 ( 
	.A1(out_sel[0]), 
	.A2(I0[27]), 
	.B1(out_sel[1]), 
	.B2(I1[27]), 
	.Z(O0[27])); 
	AO_CELL inst_1_27 ( 
	.A1(out_sel[2]), 
	.A2(I2[27]), 
	.B1(out_sel[3]), 
	.B2(I3[27]), 
	.Z(O1[27])); 
	AO_CELL inst_2_27 ( 
	.A1(out_sel[4]), 
	.A2(I4[27]), 
	.B1(out_sel[5]), 
	.B2(I5[27]), 
	.Z(O2[27])); 
	AO_CELL inst_3_27 ( 
	.A1(out_sel[6]), 
	.A2(I6[27]), 
	.B1(out_sel[7]), 
	.B2(I7[27]), 
	.Z(O3[27])); 
	AO_CELL inst_4_27 ( 
	.A1(out_sel[8]), 
	.A2(I8[27]), 
	.B1(out_sel[9]), 
	.B2(I9[27]), 
	.Z(O4[27])); 
	AO_CELL inst_5_27 ( 
	.A1(out_sel[10]), 
	.A2(I10[27]), 
	.B1(out_sel[11]), 
	.B2(I11[27]), 
	.Z(O5[27])); 
	AN_CELL inst_and_27 ( 
	.A1(out_sel[12]), 
	.A2(I12[27]), 
	.Z(O6[27])); 
	AO_CELL inst_0_28 ( 
	.A1(out_sel[0]), 
	.A2(I0[28]), 
	.B1(out_sel[1]), 
	.B2(I1[28]), 
	.Z(O0[28])); 
	AO_CELL inst_1_28 ( 
	.A1(out_sel[2]), 
	.A2(I2[28]), 
	.B1(out_sel[3]), 
	.B2(I3[28]), 
	.Z(O1[28])); 
	AO_CELL inst_2_28 ( 
	.A1(out_sel[4]), 
	.A2(I4[28]), 
	.B1(out_sel[5]), 
	.B2(I5[28]), 
	.Z(O2[28])); 
	AO_CELL inst_3_28 ( 
	.A1(out_sel[6]), 
	.A2(I6[28]), 
	.B1(out_sel[7]), 
	.B2(I7[28]), 
	.Z(O3[28])); 
	AO_CELL inst_4_28 ( 
	.A1(out_sel[8]), 
	.A2(I8[28]), 
	.B1(out_sel[9]), 
	.B2(I9[28]), 
	.Z(O4[28])); 
	AO_CELL inst_5_28 ( 
	.A1(out_sel[10]), 
	.A2(I10[28]), 
	.B1(out_sel[11]), 
	.B2(I11[28]), 
	.Z(O5[28])); 
	AN_CELL inst_and_28 ( 
	.A1(out_sel[12]), 
	.A2(I12[28]), 
	.Z(O6[28])); 
	AO_CELL inst_0_29 ( 
	.A1(out_sel[0]), 
	.A2(I0[29]), 
	.B1(out_sel[1]), 
	.B2(I1[29]), 
	.Z(O0[29])); 
	AO_CELL inst_1_29 ( 
	.A1(out_sel[2]), 
	.A2(I2[29]), 
	.B1(out_sel[3]), 
	.B2(I3[29]), 
	.Z(O1[29])); 
	AO_CELL inst_2_29 ( 
	.A1(out_sel[4]), 
	.A2(I4[29]), 
	.B1(out_sel[5]), 
	.B2(I5[29]), 
	.Z(O2[29])); 
	AO_CELL inst_3_29 ( 
	.A1(out_sel[6]), 
	.A2(I6[29]), 
	.B1(out_sel[7]), 
	.B2(I7[29]), 
	.Z(O3[29])); 
	AO_CELL inst_4_29 ( 
	.A1(out_sel[8]), 
	.A2(I8[29]), 
	.B1(out_sel[9]), 
	.B2(I9[29]), 
	.Z(O4[29])); 
	AO_CELL inst_5_29 ( 
	.A1(out_sel[10]), 
	.A2(I10[29]), 
	.B1(out_sel[11]), 
	.B2(I11[29]), 
	.Z(O5[29])); 
	AN_CELL inst_and_29 ( 
	.A1(out_sel[12]), 
	.A2(I12[29]), 
	.Z(O6[29])); 
	AO_CELL inst_0_30 ( 
	.A1(out_sel[0]), 
	.A2(I0[30]), 
	.B1(out_sel[1]), 
	.B2(I1[30]), 
	.Z(O0[30])); 
	AO_CELL inst_1_30 ( 
	.A1(out_sel[2]), 
	.A2(I2[30]), 
	.B1(out_sel[3]), 
	.B2(I3[30]), 
	.Z(O1[30])); 
	AO_CELL inst_2_30 ( 
	.A1(out_sel[4]), 
	.A2(I4[30]), 
	.B1(out_sel[5]), 
	.B2(I5[30]), 
	.Z(O2[30])); 
	AO_CELL inst_3_30 ( 
	.A1(out_sel[6]), 
	.A2(I6[30]), 
	.B1(out_sel[7]), 
	.B2(I7[30]), 
	.Z(O3[30])); 
	AO_CELL inst_4_30 ( 
	.A1(out_sel[8]), 
	.A2(I8[30]), 
	.B1(out_sel[9]), 
	.B2(I9[30]), 
	.Z(O4[30])); 
	AO_CELL inst_5_30 ( 
	.A1(out_sel[10]), 
	.A2(I10[30]), 
	.B1(out_sel[11]), 
	.B2(I11[30]), 
	.Z(O5[30])); 
	AN_CELL inst_and_30 ( 
	.A1(out_sel[12]), 
	.A2(I12[30]), 
	.Z(O6[30])); 
	AO_CELL inst_0_31 ( 
	.A1(out_sel[0]), 
	.A2(I0[31]), 
	.B1(out_sel[1]), 
	.B2(I1[31]), 
	.Z(O0[31])); 
	AO_CELL inst_1_31 ( 
	.A1(out_sel[2]), 
	.A2(I2[31]), 
	.B1(out_sel[3]), 
	.B2(I3[31]), 
	.Z(O1[31])); 
	AO_CELL inst_2_31 ( 
	.A1(out_sel[4]), 
	.A2(I4[31]), 
	.B1(out_sel[5]), 
	.B2(I5[31]), 
	.Z(O2[31])); 
	AO_CELL inst_3_31 ( 
	.A1(out_sel[6]), 
	.A2(I6[31]), 
	.B1(out_sel[7]), 
	.B2(I7[31]), 
	.Z(O3[31])); 
	AO_CELL inst_4_31 ( 
	.A1(out_sel[8]), 
	.A2(I8[31]), 
	.B1(out_sel[9]), 
	.B2(I9[31]), 
	.Z(O4[31])); 
	AO_CELL inst_5_31 ( 
	.A1(out_sel[10]), 
	.A2(I10[31]), 
	.B1(out_sel[11]), 
	.B2(I11[31]), 
	.Z(O5[31])); 
	AN_CELL inst_and_31 ( 
	.A1(out_sel[12]), 
	.A2(I12[31]), 
	.Z(O6[31])); 
endmodule 

module mantle_wire__typeBitIn32 (
    output [31:0] in,
    input [31:0] out
);
assign in = out;
endmodule

module mantle_wire__typeBitIn17 (
    output [16:0] in,
    input [16:0] out
);
assign in = out;
endmodule

module mantle_wire__typeBit8 (
    input [7:0] in,
    output [7:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit4 (
    input [3:0] in,
    output [3:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit32 (
    input [31:0] in,
    output [31:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit17 (
    input [16:0] in,
    output [16:0] out
);
assign out = in;
endmodule

module regCE_arst #(
    parameter width = 1,
    parameter init = 1
) (
    input [width-1:0] in,
    input ce,
    output [width-1:0] out,
    input clk,
    input arst
);
  reg [width-1:0] value;
  always @(posedge clk, posedge arst) begin
    if (arst) begin
      value <= init;
    end
    else if (ce) begin
      value <= in;
    end
  end
  assign out = value;
endmodule

module io_core (
  input logic clk,
  input logic clk_en,
  input logic f2io_1,
  input logic [16:0] f2io_17,
  input logic f2io_17_valid,
  input logic f2io_1_valid,
  input logic flush,
  input logic glb2io_1,
  input logic [16:0] glb2io_17,
  input logic glb2io_17_valid,
  input logic glb2io_1_valid,
  input logic io2f_17_ready,
  input logic io2f_1_ready,
  input logic io2glb_17_ready,
  input logic io2glb_1_ready,
  input logic rst_n,
  input logic tile_en,
  output logic f2io_17_ready,
  output logic f2io_1_ready,
  output logic glb2io_17_ready,
  output logic glb2io_1_ready,
  output logic io2f_1,
  output logic [16:0] io2f_17,
  output logic io2f_17_valid,
  output logic io2f_1_valid,
  output logic io2glb_1,
  output logic [16:0] io2glb_17,
  output logic io2glb_17_valid,
  output logic io2glb_1_valid
);

logic [0:0][16:0] f2io_2_io2glb_17_data_out;
logic f2io_2_io2glb_17_empty;
logic f2io_2_io2glb_17_full;
logic [0:0] f2io_2_io2glb_1_data_out;
logic f2io_2_io2glb_1_empty;
logic f2io_2_io2glb_1_full;
logic gclk;
logic glb2io_2_io2f_17_empty;
logic glb2io_2_io2f_17_full;
logic glb2io_2_io2f_1_empty;
logic glb2io_2_io2f_1_full;
assign gclk = clk & tile_en;
assign io2glb_1 = f2io_2_io2glb_1_data_out;
assign f2io_1_ready = ~f2io_2_io2glb_1_full;
assign io2glb_1_valid = ~f2io_2_io2glb_1_empty;
assign glb2io_1_ready = ~glb2io_2_io2f_1_full;
assign io2f_1_valid = ~glb2io_2_io2f_1_empty;
assign io2glb_17 = f2io_2_io2glb_17_data_out[0][16:0];
assign f2io_17_ready = ~f2io_2_io2glb_17_full;
assign io2glb_17_valid = ~f2io_2_io2glb_17_empty;
assign glb2io_17_ready = ~glb2io_2_io2f_17_full;
assign io2f_17_valid = ~glb2io_2_io2f_17_empty;
reg_fifo_depth_2_w_1_afd_1_iocore_nof f2io_2_io2glb_1 (
  .clk(clk),
  .clk_en(clk_en),
  .data_in(f2io_1),
  .flush(flush),
  .pop(io2glb_1_ready),
  .push(f2io_1_valid),
  .rst_n(rst_n),
  .data_out(f2io_2_io2glb_1_data_out),
  .empty(f2io_2_io2glb_1_empty),
  .full(f2io_2_io2glb_1_full)
);

reg_fifo_depth_2_w_1_afd_1_iocore_nof glb2io_2_io2f_1 (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(glb2io_1),
  .flush(flush),
  .pop(io2f_1_ready),
  .push(glb2io_1_valid),
  .rst_n(rst_n),
  .data_out(io2f_1),
  .empty(glb2io_2_io2f_1_empty),
  .full(glb2io_2_io2f_1_full)
);

reg_fifo_depth_2_w_17_afd_1_iocore_nof f2io_2_io2glb_17 (
  .clk(clk),
  .clk_en(clk_en),
  .data_in(f2io_17),
  .flush(flush),
  .pop(io2glb_17_ready),
  .push(f2io_17_valid),
  .rst_n(rst_n),
  .data_out(f2io_2_io2glb_17_data_out),
  .empty(f2io_2_io2glb_17_empty),
  .full(f2io_2_io2glb_17_full)
);

reg_fifo_depth_2_w_17_afd_1_iocore_nof glb2io_2_io2f_17 (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(glb2io_17),
  .flush(flush),
  .pop(io2f_17_ready),
  .push(glb2io_17_valid),
  .rst_n(rst_n),
  .data_out(io2f_17),
  .empty(glb2io_2_io2f_17_empty),
  .full(glb2io_2_io2f_17_full)
);

endmodule   // io_core

module io_core_W (
  input logic clk,
  input logic clk_en,
  input logic f2io_1,
  input logic [16:0] f2io_17,
  input logic f2io_17_valid,
  input logic f2io_1_valid,
  input logic flush,
  input logic glb2io_1,
  input logic [16:0] glb2io_17,
  input logic glb2io_17_valid,
  input logic glb2io_1_valid,
  input logic io2f_17_ready,
  input logic io2f_1_ready,
  input logic io2glb_17_ready,
  input logic io2glb_1_ready,
  input logic rst_n,
  input logic tile_en,
  output logic f2io_17_ready,
  output logic f2io_1_ready,
  output logic glb2io_17_ready,
  output logic glb2io_1_ready,
  output logic io2f_1,
  output logic [16:0] io2f_17,
  output logic io2f_17_valid,
  output logic io2f_1_valid,
  output logic io2glb_1,
  output logic [16:0] io2glb_17,
  output logic io2glb_17_valid,
  output logic io2glb_1_valid
);

io_core io_core (
  .clk(clk),
  .clk_en(clk_en),
  .f2io_1(f2io_1),
  .f2io_17(f2io_17),
  .f2io_17_valid(f2io_17_valid),
  .f2io_1_valid(f2io_1_valid),
  .flush(flush),
  .glb2io_1(glb2io_1),
  .glb2io_17(glb2io_17),
  .glb2io_17_valid(glb2io_17_valid),
  .glb2io_1_valid(glb2io_1_valid),
  .io2f_17_ready(io2f_17_ready),
  .io2f_1_ready(io2f_1_ready),
  .io2glb_17_ready(io2glb_17_ready),
  .io2glb_1_ready(io2glb_1_ready),
  .rst_n(rst_n),
  .tile_en(tile_en),
  .f2io_17_ready(f2io_17_ready),
  .f2io_1_ready(f2io_1_ready),
  .glb2io_17_ready(glb2io_17_ready),
  .glb2io_1_ready(glb2io_1_ready),
  .io2f_1(io2f_1),
  .io2f_17(io2f_17),
  .io2f_17_valid(io2f_17_valid),
  .io2f_1_valid(io2f_1_valid),
  .io2glb_1(io2glb_1),
  .io2glb_17(io2glb_17),
  .io2glb_17_valid(io2glb_17_valid),
  .io2glb_1_valid(io2glb_1_valid)
);

endmodule   // io_core_W

module reg_fifo_depth_2_w_17_afd_1_iocore_nof (
  input logic clk,
  input logic clk_en,
  input logic [0:0] [16:0] data_in,
  input logic flush,
  input logic pop,
  input logic push,
  input logic rst_n,
  output logic almost_full,
  output logic [0:0] [16:0] data_out,
  output logic empty,
  output logic full,
  output logic valid
);

logic [1:0] num_items;
logic passthru;
logic rd_ptr;
logic read;
logic [1:0][0:0][16:0] reg_array;
logic wr_ptr;
logic write;
assign full = num_items == 2'h2;
assign almost_full = num_items >= 2'h1;
assign empty = num_items == 2'h0;
assign read = pop & (~passthru) & (~empty);
assign passthru = 1'h0;
assign write = push & (~passthru) & (~full);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_items <= 2'h0;
  end
  else if (flush) begin
    num_items <= 2'h0;
  end
  else if (clk_en) begin
    if (write & (~read)) begin
      num_items <= num_items + 2'h1;
    end
    else if ((~write) & read) begin
      num_items <= num_items - 2'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    reg_array <= 34'h0;
  end
  else if (flush) begin
    reg_array <= 34'h0;
  end
  else if (clk_en) begin
    if (write) begin
      reg_array[wr_ptr] <= data_in;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    wr_ptr <= 1'h0;
  end
  else if (flush) begin
    wr_ptr <= 1'h0;
  end
  else if (clk_en) begin
    if (write) begin
      if (wr_ptr == 1'h1) begin
        wr_ptr <= 1'h0;
      end
      else wr_ptr <= wr_ptr + 1'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    rd_ptr <= 1'h0;
  end
  else if (flush) begin
    rd_ptr <= 1'h0;
  end
  else if (clk_en) begin
    if (read) begin
      rd_ptr <= rd_ptr + 1'h1;
    end
  end
end
always_comb begin
  if (passthru) begin
    data_out = data_in;
  end
  else data_out = reg_array[rd_ptr];
end
always_comb begin
  valid = (~empty) | passthru;
end
endmodule   // reg_fifo_depth_2_w_17_afd_1_iocore_nof

module reg_fifo_depth_2_w_1_afd_1_iocore_nof (
  input logic clk,
  input logic clk_en,
  input logic [0:0] data_in,
  input logic flush,
  input logic pop,
  input logic push,
  input logic rst_n,
  output logic almost_full,
  output logic [0:0] data_out,
  output logic empty,
  output logic full,
  output logic valid
);

logic [1:0] num_items;
logic passthru;
logic rd_ptr;
logic read;
logic [1:0][0:0] reg_array;
logic wr_ptr;
logic write;
assign full = num_items == 2'h2;
assign almost_full = num_items >= 2'h1;
assign empty = num_items == 2'h0;
assign read = pop & (~passthru) & (~empty);
assign passthru = 1'h0;
assign write = push & (~passthru) & (~full);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_items <= 2'h0;
  end
  else if (flush) begin
    num_items <= 2'h0;
  end
  else if (clk_en) begin
    if (write & (~read)) begin
      num_items <= num_items + 2'h1;
    end
    else if ((~write) & read) begin
      num_items <= num_items - 2'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    reg_array <= 2'h0;
  end
  else if (flush) begin
    reg_array <= 2'h0;
  end
  else if (clk_en) begin
    if (write) begin
      reg_array[wr_ptr] <= data_in;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    wr_ptr <= 1'h0;
  end
  else if (flush) begin
    wr_ptr <= 1'h0;
  end
  else if (clk_en) begin
    if (write) begin
      if (wr_ptr == 1'h1) begin
        wr_ptr <= 1'h0;
      end
      else wr_ptr <= wr_ptr + 1'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    rd_ptr <= 1'h0;
  end
  else if (flush) begin
    rd_ptr <= 1'h0;
  end
  else if (clk_en) begin
    if (read) begin
      rd_ptr <= rd_ptr + 1'h1;
    end
  end
end
always_comb begin
  if (passthru) begin
    data_out = data_in;
  end
  else data_out = reg_array[rd_ptr];
end
always_comb begin
  valid = (~empty) | passthru;
end
endmodule   // reg_fifo_depth_2_w_1_afd_1_iocore_nof


typedef struct packed {
    logic [1:0] west;
    logic [1:0] east;
    logic [1:0] south;
} pcfg_broadcast_mux_t;

typedef struct packed {
    logic rd_en;
    logic [18:0] rd_addr;
} rdrq_packet_t;

typedef struct packed {
    logic wr_en;
    logic [7:0] wr_strb;
    logic [16:0] wr_addr;
    logic [63:0] wr_data;
} wr_bank_packet_t;

typedef struct packed {
    logic mode;
    logic [15:0] relocation_value;
    logic relocation_is_msb;
} pcfg_dma_ctrl_t;

typedef struct packed {
    logic wr_en;
    logic [7:0] wr_strb;
    logic [18:0] wr_addr;
    logic [63:0] wr_data;
} wr_packet_t;

typedef struct packed {
    logic [1:0] mode;
    logic [1:0] valid_mode;
    logic [1:0] data_mux;
    logic num_repeat;
} store_dma_ctrl_t;

typedef struct packed {
    logic tile_connected;
    logic [5:0] latency;
} cfg_pcfg_network_t;

typedef struct packed {
    logic tile_connected;
    logic [5:0] latency;
} cfg_data_network_t;

typedef struct packed {
    logic rd_en;
    logic wr_en;
    logic [31:0] addr;
    logic [31:0] data;
} cgra_cfg_t;

typedef struct packed {
    logic [63:0] rd_data;
    logic rd_data_valid;
} rdrs_packet_t;

typedef struct packed {
wr_packet_t wr;
rdrq_packet_t rdrq;
rdrs_packet_t rdrs;
} packet_t;

typedef struct packed {
    logic [1:0] mode;
    logic [1:0] valid_mode;
    logic flush_mode;
    logic [1:0] data_mux;
    logic num_repeat;
} load_dma_ctrl_t;

typedef struct packed {
    logic [18:0] start_addr;
    logic [15:0] cycle_start_addr;
    logic [3:0] dim;
    logic [31:0] range_0;
    logic [19:0] stride_0;
    logic [15:0] cycle_stride_0;
    logic [31:0] range_1;
    logic [19:0] stride_1;
    logic [15:0] cycle_stride_1;
    logic [31:0] range_2;
    logic [19:0] stride_2;
    logic [15:0] cycle_stride_2;
    logic [31:0] range_3;
    logic [19:0] stride_3;
    logic [15:0] cycle_stride_3;
    logic [31:0] range_4;
    logic [19:0] stride_4;
    logic [15:0] cycle_stride_4;
    logic [31:0] range_5;
    logic [19:0] stride_5;
    logic [15:0] cycle_stride_5;
    logic [31:0] range_6;
    logic [19:0] stride_6;
    logic [15:0] cycle_stride_6;
    logic [31:0] range_7;
    logic [19:0] stride_7;
    logic [15:0] cycle_stride_7;
} load_dma_header_t;

typedef struct packed {
    logic [18:0] start_addr;
    logic [15:0] num_cfg;
} pcfg_dma_header_t;

typedef struct packed {
rdrq_packet_t rdrq;
rdrs_packet_t rdrs;
} rd_packet_t;

typedef struct packed {
    logic rd_en;
    logic [16:0] rd_addr;
} rdrq_bank_packet_t;

typedef struct packed {
    logic [18:0] start_addr;
    logic [15:0] cycle_start_addr;
    logic [3:0] dim;
    logic [31:0] range_0;
    logic [19:0] stride_0;
    logic [15:0] cycle_stride_0;
    logic [31:0] range_1;
    logic [19:0] stride_1;
    logic [15:0] cycle_stride_1;
    logic [31:0] range_2;
    logic [19:0] stride_2;
    logic [15:0] cycle_stride_2;
    logic [31:0] range_3;
    logic [19:0] stride_3;
    logic [15:0] cycle_stride_3;
    logic [31:0] range_4;
    logic [19:0] stride_4;
    logic [15:0] cycle_stride_4;
    logic [31:0] range_5;
    logic [19:0] stride_5;
    logic [15:0] cycle_stride_5;
    logic [31:0] range_6;
    logic [19:0] stride_6;
    logic [15:0] cycle_stride_6;
} store_dma_header_t;

interface glb_tile_ifc_A_12_D_32;
  logic [11:0] rd_addr;
  logic rd_clk_en;
  logic [31:0] rd_data;
  logic rd_data_valid;
  logic rd_en;
  logic [11:0] wr_addr;
  logic wr_clk_en;
  logic [31:0] wr_data;
  logic wr_en;
  modport master(input rd_data, input rd_data_valid, output rd_addr, output rd_clk_en, output rd_en, output wr_addr, output wr_clk_en, output wr_data, output wr_en);
  modport slave(input rd_addr, input rd_clk_en, input rd_en, input wr_addr, input wr_clk_en, input wr_data, input wr_en, output rd_data, output rd_data_valid);
endinterface

interface glb_tile_ifc_A_19_D_32;
  logic [18:0] rd_addr;
  logic rd_clk_en;
  logic [31:0] rd_data;
  logic rd_data_valid;
  logic rd_en;
  logic [18:0] wr_addr;
  logic wr_clk_en;
  logic [31:0] wr_data;
  logic wr_en;
  modport master(input rd_data, input rd_data_valid, output rd_addr, output rd_clk_en, output rd_en, output wr_addr, output wr_clk_en, output wr_data, output wr_en);
  modport slave(input rd_addr, input rd_clk_en, input rd_en, input wr_addr, input wr_clk_en, input wr_data, input wr_en, output rd_data, output rd_data_valid);
endinterface

interface glb_tile_ifc_A_19_D_64;
  logic [18:0] rd_addr;
  logic rd_clk_en;
  logic [63:0] rd_data;
  logic rd_data_valid;
  logic rd_en;
  logic [18:0] wr_addr;
  logic wr_clk_en;
  logic [63:0] wr_data;
  logic wr_en;
  logic [7:0] wr_strb;
  modport master(input rd_data, input rd_data_valid, output rd_addr, output rd_clk_en, output rd_en, output wr_addr, output wr_clk_en, output wr_data, output wr_en, output wr_strb);
  modport slave(input rd_addr, input rd_clk_en, input rd_en, input wr_addr, input wr_clk_en, input wr_data, input wr_en, input wr_strb, output rd_data, output rd_data_valid);
endinterface

module IN12LP_S1DB_W04096B064M08S2_HB (
  input logic [11:0] A,
  input logic [63:0] BW,
  input logic CEN,
  input logic CLK,
  input logic [63:0] D,
  input logic MA_SAWL0,
  input logic MA_SAWL1,
  input logic MA_STABAS0,
  input logic MA_STABAS1,
  input logic MA_VD0,
  input logic MA_VD1,
  input logic MA_WL0,
  input logic MA_WL1,
  input logic MA_WRAS0,
  input logic MA_WRAS1,
  input logic MA_WRT,
  input logic RDWEN,
  input logic T_LOGIC,
  input logic T_Q_RST,
  output logic [63:0] Q
);

logic [63:0] data_array [4095:0];

always_ff @(posedge CLK) begin
  if (CEN == 1'h0) begin
    Q <= data_array[A];
    if (RDWEN == 1'h0) begin
      for (int unsigned i = 0; i < 64; i += 1) begin
          if (BW[6'(i)]) begin
            data_array[A][6'(i)] <= D[6'(i)];
          end
        end
    end
  end
end
endmodule   // IN12LP_S1DB_W04096B064M08S2_HB

module SC7P5T_CKGPRELATNX1_SSC14R (
  input logic CLK,
  input logic E,
  input logic TE,
  output logic Z
);

logic enable_latch;
always_latch begin
  if (~CLK) begin
    enable_latch = E;
  end
end
assign Z = CLK & enable_latch;
endmodule   // SC7P5T_CKGPRELATNX1_SSC14R

module clk_gate (
  input logic clk,
  input logic enable,
  output logic gclk
);

SC7P5T_CKGPRELATNX1_SSC14R CG_CELL (
  .CLK(clk),
  .E(enable),
  .TE(1'h0),
  .Z(gclk)
);

endmodule   // clk_gate

module glb_addr_gen_7 #(
  parameter addr_width = 32'h10,
  parameter loop_level = 32'h7
)
(
  input logic clk,
  input logic clk_en,
  input logic [2:0] mux_sel,
  input logic reset,
  input logic restart,
  input logic [addr_width-1:0] start_addr,
  input logic step,
  input logic [loop_level-1:0] [addr_width-1:0] strides,
  output logic [addr_width-1:0] addr_out
);

logic [addr_width-1:0] current_addr;
assign addr_out = start_addr + current_addr;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    current_addr <= 16'h0;
  end
  else if (clk_en) begin
    if (restart) begin
      current_addr <= 16'h0;
    end
    else if (step) begin
      current_addr <= current_addr + strides[mux_sel];
    end
  end
end
endmodule   // glb_addr_gen_7

module glb_addr_gen_8 #(
  parameter addr_width = 32'h10,
  parameter loop_level = 32'h8
)
(
  input logic clk,
  input logic clk_en,
  input logic [2:0] mux_sel,
  input logic reset,
  input logic restart,
  input logic [addr_width-1:0] start_addr,
  input logic step,
  input logic [loop_level-1:0] [addr_width-1:0] strides,
  output logic [addr_width-1:0] addr_out
);

logic [addr_width-1:0] current_addr;
assign addr_out = start_addr + current_addr;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    current_addr <= 16'h0;
  end
  else if (clk_en) begin
    if (restart) begin
      current_addr <= 16'h0;
    end
    else if (step) begin
      current_addr <= current_addr + strides[mux_sel];
    end
  end
end
endmodule   // glb_addr_gen_8

module glb_bank (
  input logic clk,
  input rdrq_bank_packet_t rdrq_packet,
  input logic reset,
  input wr_bank_packet_t wr_packet,
  output rdrs_packet_t rdrs_packet
);

logic [16:0] mem_addr;
logic [63:0] mem_data_in;
logic [63:0] mem_data_in_bit_sel;
logic [63:0] mem_data_out;
logic mem_rd_en;
logic mem_wr_en;
logic [63:0] packet_rd_data_r;
logic packet_rd_en_d;
logic [63:0] wr_data_bit_sel;
assign wr_data_bit_sel[0] = wr_packet.wr_strb[0];
assign wr_data_bit_sel[1] = wr_packet.wr_strb[0];
assign wr_data_bit_sel[2] = wr_packet.wr_strb[0];
assign wr_data_bit_sel[3] = wr_packet.wr_strb[0];
assign wr_data_bit_sel[4] = wr_packet.wr_strb[0];
assign wr_data_bit_sel[5] = wr_packet.wr_strb[0];
assign wr_data_bit_sel[6] = wr_packet.wr_strb[0];
assign wr_data_bit_sel[7] = wr_packet.wr_strb[0];
assign wr_data_bit_sel[8] = wr_packet.wr_strb[1];
assign wr_data_bit_sel[9] = wr_packet.wr_strb[1];
assign wr_data_bit_sel[10] = wr_packet.wr_strb[1];
assign wr_data_bit_sel[11] = wr_packet.wr_strb[1];
assign wr_data_bit_sel[12] = wr_packet.wr_strb[1];
assign wr_data_bit_sel[13] = wr_packet.wr_strb[1];
assign wr_data_bit_sel[14] = wr_packet.wr_strb[1];
assign wr_data_bit_sel[15] = wr_packet.wr_strb[1];
assign wr_data_bit_sel[16] = wr_packet.wr_strb[2];
assign wr_data_bit_sel[17] = wr_packet.wr_strb[2];
assign wr_data_bit_sel[18] = wr_packet.wr_strb[2];
assign wr_data_bit_sel[19] = wr_packet.wr_strb[2];
assign wr_data_bit_sel[20] = wr_packet.wr_strb[2];
assign wr_data_bit_sel[21] = wr_packet.wr_strb[2];
assign wr_data_bit_sel[22] = wr_packet.wr_strb[2];
assign wr_data_bit_sel[23] = wr_packet.wr_strb[2];
assign wr_data_bit_sel[24] = wr_packet.wr_strb[3];
assign wr_data_bit_sel[25] = wr_packet.wr_strb[3];
assign wr_data_bit_sel[26] = wr_packet.wr_strb[3];
assign wr_data_bit_sel[27] = wr_packet.wr_strb[3];
assign wr_data_bit_sel[28] = wr_packet.wr_strb[3];
assign wr_data_bit_sel[29] = wr_packet.wr_strb[3];
assign wr_data_bit_sel[30] = wr_packet.wr_strb[3];
assign wr_data_bit_sel[31] = wr_packet.wr_strb[3];
assign wr_data_bit_sel[32] = wr_packet.wr_strb[4];
assign wr_data_bit_sel[33] = wr_packet.wr_strb[4];
assign wr_data_bit_sel[34] = wr_packet.wr_strb[4];
assign wr_data_bit_sel[35] = wr_packet.wr_strb[4];
assign wr_data_bit_sel[36] = wr_packet.wr_strb[4];
assign wr_data_bit_sel[37] = wr_packet.wr_strb[4];
assign wr_data_bit_sel[38] = wr_packet.wr_strb[4];
assign wr_data_bit_sel[39] = wr_packet.wr_strb[4];
assign wr_data_bit_sel[40] = wr_packet.wr_strb[5];
assign wr_data_bit_sel[41] = wr_packet.wr_strb[5];
assign wr_data_bit_sel[42] = wr_packet.wr_strb[5];
assign wr_data_bit_sel[43] = wr_packet.wr_strb[5];
assign wr_data_bit_sel[44] = wr_packet.wr_strb[5];
assign wr_data_bit_sel[45] = wr_packet.wr_strb[5];
assign wr_data_bit_sel[46] = wr_packet.wr_strb[5];
assign wr_data_bit_sel[47] = wr_packet.wr_strb[5];
assign wr_data_bit_sel[48] = wr_packet.wr_strb[6];
assign wr_data_bit_sel[49] = wr_packet.wr_strb[6];
assign wr_data_bit_sel[50] = wr_packet.wr_strb[6];
assign wr_data_bit_sel[51] = wr_packet.wr_strb[6];
assign wr_data_bit_sel[52] = wr_packet.wr_strb[6];
assign wr_data_bit_sel[53] = wr_packet.wr_strb[6];
assign wr_data_bit_sel[54] = wr_packet.wr_strb[6];
assign wr_data_bit_sel[55] = wr_packet.wr_strb[6];
assign wr_data_bit_sel[56] = wr_packet.wr_strb[7];
assign wr_data_bit_sel[57] = wr_packet.wr_strb[7];
assign wr_data_bit_sel[58] = wr_packet.wr_strb[7];
assign wr_data_bit_sel[59] = wr_packet.wr_strb[7];
assign wr_data_bit_sel[60] = wr_packet.wr_strb[7];
assign wr_data_bit_sel[61] = wr_packet.wr_strb[7];
assign wr_data_bit_sel[62] = wr_packet.wr_strb[7];
assign wr_data_bit_sel[63] = wr_packet.wr_strb[7];
always_comb begin
  if (wr_packet.wr_en) begin
    mem_wr_en = 1'h1;
    mem_rd_en = 1'h0;
    mem_addr = wr_packet.wr_addr;
    mem_data_in = wr_packet.wr_data;
    mem_data_in_bit_sel = wr_data_bit_sel;
  end
  else if (rdrq_packet.rd_en) begin
    mem_wr_en = 1'h0;
    mem_rd_en = 1'h1;
    mem_addr = rdrq_packet.rd_addr;
    mem_data_in = 64'h0;
    mem_data_in_bit_sel = 64'h0;
  end
  else begin
    mem_wr_en = 1'h0;
    mem_rd_en = 1'h0;
    mem_addr = 17'h0;
    mem_data_in = 64'h0;
    mem_data_in_bit_sel = 64'h0;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    packet_rd_data_r <= 64'h0;
  end
  else packet_rd_data_r <= rdrs_packet.rd_data;
end
always_comb begin
  if (packet_rd_en_d) begin
    rdrs_packet.rd_data = mem_data_out;
  end
  else rdrs_packet.rd_data = packet_rd_data_r;
  rdrs_packet.rd_data_valid = packet_rd_en_d;
end
glb_bank_memory glb_bank_memory (
  .addr(mem_addr),
  .clk(clk),
  .data_in(mem_data_in),
  .data_in_bit_sel(mem_data_in_bit_sel),
  .ren(mem_rd_en),
  .reset(reset),
  .wen(mem_wr_en),
  .data_out(mem_data_out)
);

pipeline_w_1_d_1 packet_rdrq_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(rdrq_packet.rd_en),
  .reset(reset),
  .out_(packet_rd_en_d)
);

endmodule   // glb_bank

module glb_bank_memory (
  input logic [16:0] addr,
  input logic clk,
  input logic [63:0] data_in,
  input logic [63:0] data_in_bit_sel,
  input logic ren,
  input logic reset,
  input logic wen,
  output logic [63:0] data_out
);

logic glb_bank_sram_gen_CEB;
logic glb_bank_sram_gen_WEB;
logic [13:0] sram_addr;
logic [13:0] sram_addr_d;
logic sram_cen;
logic sram_cen_d;
logic [63:0] sram_data_in;
logic [63:0] sram_data_in_bit_sel;
logic [63:0] sram_data_in_bit_sel_d;
logic [63:0] sram_data_in_d;
logic [63:0] sram_data_out;
logic [143:0] sram_signals_pipeline_in_;
logic [143:0] sram_signals_pipeline_out_;
logic sram_wen;
logic sram_wen_d;
assign sram_signals_pipeline_in_ = {sram_wen, sram_cen, sram_addr, sram_data_in, sram_data_in_bit_sel};
assign {sram_wen_d, sram_cen_d, sram_addr_d, sram_data_in_d, sram_data_in_bit_sel_d} = sram_signals_pipeline_out_;
assign glb_bank_sram_gen_CEB = ~sram_cen_d;
assign glb_bank_sram_gen_WEB = ~sram_wen_d;
always_comb begin
  sram_wen = wen;
  sram_cen = wen | ren;
  sram_addr = addr[16:3];
  sram_data_in = data_in;
  sram_data_in_bit_sel = data_in_bit_sel;
  data_out = sram_data_out;
end
pipeline_w_144_d_0 sram_signals_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(sram_signals_pipeline_in_),
  .reset(reset),
  .out_(sram_signals_pipeline_out_)
);

glb_bank_sram_gen_14 glb_bank_sram_gen (
  .A(sram_addr_d),
  .BW(sram_data_in_bit_sel_d),
  .CEB(glb_bank_sram_gen_CEB),
  .CLK(clk),
  .D(sram_data_in_d),
  .RESET(reset),
  .WEB(glb_bank_sram_gen_WEB),
  .Q(sram_data_out)
);

endmodule   // glb_bank_memory

module glb_bank_mux (
  input logic cfg_pcfg_tile_connected_next,
  input logic cfg_pcfg_tile_connected_prev,
  input logic cfg_tile_connected_next,
  input logic cfg_tile_connected_prev,
  input logic clk,
  input logic glb_tile_id,
  input rdrq_packet_t rdrq_packet_dma2bank,
  input rdrq_packet_t rdrq_packet_pcfgdma2bank,
  input rdrq_packet_t rdrq_packet_pcfgring2bank,
  input rdrq_packet_t rdrq_packet_procsw2bank,
  input rdrq_packet_t rdrq_packet_ring2bank,
  input rdrs_packet_t [1:0] rdrs_packet_bankarr2sw,
  input logic reset,
  input wr_packet_t wr_packet_dma2bank,
  input wr_packet_t wr_packet_procsw2bank,
  input wr_packet_t wr_packet_ring2bank,
  output rdrq_bank_packet_t [1:0] rdrq_packet_sw2bankarr,
  output rdrs_packet_t rdrs_packet_bank2dma,
  output rdrs_packet_t rdrs_packet_bank2pcfgdma,
  output rdrs_packet_t rdrs_packet_bank2pcfgring,
  output rdrs_packet_t rdrs_packet_bank2procsw,
  output rdrs_packet_t rdrs_packet_bank2ring,
  output wr_bank_packet_t [1:0] wr_packet_sw2bankarr
);

typedef enum logic[1:0] {
  none = 2'h0,
  proc = 2'h1,
  strm = 2'h2,
  pcfg = 2'h3
} rd_type_e;
rd_type_e rd_type_0;
rd_type_e rd_type_1;
rd_type_e rd_type_d_0;
rd_type_e rd_type_d_1;
logic [3:0] rd_type_pipeline_1_in_;
logic [3:0] rd_type_pipeline_1_out_;
rdrq_bank_packet_t [1:0] rdrq_packet_sw2bankarr_w;
logic [17:0] rdrq_sw2bank_pipeline_0_out_;
logic [17:0] rdrq_sw2bank_pipeline_1_out_;
logic [64:0] rdrs_bank2sw_pipeline_0_out_;
logic [64:0] rdrs_bank2sw_pipeline_1_out_;
rdrs_packet_t [1:0] rdrs_packet_bankarr2sw_d;
wr_bank_packet_t [1:0] wr_packet_sw2bankarr_w;
logic [89:0] wr_sw2bank_pipeline_0_out_;
logic [89:0] wr_sw2bank_pipeline_1_out_;
assign wr_packet_sw2bankarr[0] = wr_sw2bank_pipeline_0_out_;
assign wr_packet_sw2bankarr[1] = wr_sw2bank_pipeline_1_out_;
assign rdrq_packet_sw2bankarr[0] = rdrq_sw2bank_pipeline_0_out_;
assign rdrq_packet_sw2bankarr[1] = rdrq_sw2bank_pipeline_1_out_;
assign rd_type_pipeline_1_in_ = {rd_type_0, rd_type_1};
assign {rd_type_d_0, rd_type_d_1} = rd_type_pipeline_1_out_;
assign rdrs_packet_bankarr2sw_d[0] = rdrs_bank2sw_pipeline_0_out_;
assign rdrs_packet_bankarr2sw_d[1] = rdrs_bank2sw_pipeline_1_out_;
always_comb begin
  if ((wr_packet_procsw2bank.wr_en == 1'h1) & (wr_packet_procsw2bank.wr_addr[18] == glb_tile_id) & (wr_packet_procsw2bank.wr_addr[17] == 1'h0)) begin
    wr_packet_sw2bankarr_w[0].wr_en = wr_packet_procsw2bank.wr_en;
    wr_packet_sw2bankarr_w[0].wr_addr = wr_packet_procsw2bank.wr_addr[16:0];
    wr_packet_sw2bankarr_w[0].wr_strb = wr_packet_procsw2bank.wr_strb;
    wr_packet_sw2bankarr_w[0].wr_data = wr_packet_procsw2bank.wr_data;
  end
  else if ((wr_packet_dma2bank.wr_en == 1'h1) & (~cfg_tile_connected_prev) & (~cfg_tile_connected_next) & (wr_packet_dma2bank.wr_addr[18] == glb_tile_id) & (wr_packet_dma2bank.wr_addr[17] == 1'h0)) begin
    wr_packet_sw2bankarr_w[0].wr_en = wr_packet_dma2bank.wr_en;
    wr_packet_sw2bankarr_w[0].wr_addr = wr_packet_dma2bank.wr_addr[16:0];
    wr_packet_sw2bankarr_w[0].wr_strb = wr_packet_dma2bank.wr_strb;
    wr_packet_sw2bankarr_w[0].wr_data = wr_packet_dma2bank.wr_data;
  end
  else if ((wr_packet_ring2bank.wr_en == 1'h1) & (wr_packet_ring2bank.wr_addr[18] == glb_tile_id) & (wr_packet_ring2bank.wr_addr[17] == 1'h0)) begin
    wr_packet_sw2bankarr_w[0].wr_en = wr_packet_ring2bank.wr_en;
    wr_packet_sw2bankarr_w[0].wr_addr = wr_packet_ring2bank.wr_addr[16:0];
    wr_packet_sw2bankarr_w[0].wr_strb = wr_packet_ring2bank.wr_strb;
    wr_packet_sw2bankarr_w[0].wr_data = wr_packet_ring2bank.wr_data;
  end
  else wr_packet_sw2bankarr_w[0] = 90'h0;
end
always_comb begin
  if ((wr_packet_procsw2bank.wr_en == 1'h1) & (wr_packet_procsw2bank.wr_addr[18] == glb_tile_id) & (wr_packet_procsw2bank.wr_addr[17] == 1'h1)) begin
    wr_packet_sw2bankarr_w[1].wr_en = wr_packet_procsw2bank.wr_en;
    wr_packet_sw2bankarr_w[1].wr_addr = wr_packet_procsw2bank.wr_addr[16:0];
    wr_packet_sw2bankarr_w[1].wr_strb = wr_packet_procsw2bank.wr_strb;
    wr_packet_sw2bankarr_w[1].wr_data = wr_packet_procsw2bank.wr_data;
  end
  else if ((wr_packet_dma2bank.wr_en == 1'h1) & (~cfg_tile_connected_prev) & (~cfg_tile_connected_next) & (wr_packet_dma2bank.wr_addr[18] == glb_tile_id) & (wr_packet_dma2bank.wr_addr[17] == 1'h1)) begin
    wr_packet_sw2bankarr_w[1].wr_en = wr_packet_dma2bank.wr_en;
    wr_packet_sw2bankarr_w[1].wr_addr = wr_packet_dma2bank.wr_addr[16:0];
    wr_packet_sw2bankarr_w[1].wr_strb = wr_packet_dma2bank.wr_strb;
    wr_packet_sw2bankarr_w[1].wr_data = wr_packet_dma2bank.wr_data;
  end
  else if ((wr_packet_ring2bank.wr_en == 1'h1) & (wr_packet_ring2bank.wr_addr[18] == glb_tile_id) & (wr_packet_ring2bank.wr_addr[17] == 1'h1)) begin
    wr_packet_sw2bankarr_w[1].wr_en = wr_packet_ring2bank.wr_en;
    wr_packet_sw2bankarr_w[1].wr_addr = wr_packet_ring2bank.wr_addr[16:0];
    wr_packet_sw2bankarr_w[1].wr_strb = wr_packet_ring2bank.wr_strb;
    wr_packet_sw2bankarr_w[1].wr_data = wr_packet_ring2bank.wr_data;
  end
  else wr_packet_sw2bankarr_w[1] = 90'h0;
end
always_comb begin
  if ((rdrq_packet_procsw2bank.rd_en == 1'h1) & (rdrq_packet_procsw2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_procsw2bank.rd_addr[17] == 1'h0)) begin
    rdrq_packet_sw2bankarr_w[0].rd_en = rdrq_packet_procsw2bank.rd_en;
    rdrq_packet_sw2bankarr_w[0].rd_addr = rdrq_packet_procsw2bank.rd_addr[16:0];
    rd_type_0 = proc;
  end
  else if ((rdrq_packet_pcfgdma2bank.rd_en == 1'h1) & (~cfg_pcfg_tile_connected_prev) & (~cfg_pcfg_tile_connected_next) & (rdrq_packet_pcfgdma2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_pcfgdma2bank.rd_addr[17] == 1'h0)) begin
    rdrq_packet_sw2bankarr_w[0].rd_en = rdrq_packet_pcfgdma2bank.rd_en;
    rdrq_packet_sw2bankarr_w[0].rd_addr = rdrq_packet_pcfgdma2bank.rd_addr[16:0];
    rd_type_0 = pcfg;
  end
  else if ((rdrq_packet_pcfgring2bank.rd_en == 1'h1) & (rdrq_packet_pcfgring2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_pcfgring2bank.rd_addr[17] == 1'h0)) begin
    rdrq_packet_sw2bankarr_w[0].rd_en = rdrq_packet_pcfgring2bank.rd_en;
    rdrq_packet_sw2bankarr_w[0].rd_addr = rdrq_packet_pcfgring2bank.rd_addr[16:0];
    rd_type_0 = pcfg;
  end
  else if ((rdrq_packet_dma2bank.rd_en == 1'h1) & (~cfg_tile_connected_prev) & (~cfg_tile_connected_next) & (rdrq_packet_dma2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_dma2bank.rd_addr[17] == 1'h0)) begin
    rdrq_packet_sw2bankarr_w[0].rd_en = rdrq_packet_dma2bank.rd_en;
    rdrq_packet_sw2bankarr_w[0].rd_addr = rdrq_packet_dma2bank.rd_addr[16:0];
    rd_type_0 = strm;
  end
  else if ((rdrq_packet_ring2bank.rd_en == 1'h1) & (rdrq_packet_ring2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_ring2bank.rd_addr[17] == 1'h0)) begin
    rdrq_packet_sw2bankarr_w[0].rd_en = rdrq_packet_ring2bank.rd_en;
    rdrq_packet_sw2bankarr_w[0].rd_addr = rdrq_packet_ring2bank.rd_addr[16:0];
    rd_type_0 = strm;
  end
  else begin
    rdrq_packet_sw2bankarr_w[0] = 18'h0;
    rd_type_0 = none;
  end
end
always_comb begin
  if ((rdrq_packet_procsw2bank.rd_en == 1'h1) & (rdrq_packet_procsw2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_procsw2bank.rd_addr[17] == 1'h1)) begin
    rdrq_packet_sw2bankarr_w[1].rd_en = rdrq_packet_procsw2bank.rd_en;
    rdrq_packet_sw2bankarr_w[1].rd_addr = rdrq_packet_procsw2bank.rd_addr[16:0];
    rd_type_1 = proc;
  end
  else if ((rdrq_packet_pcfgdma2bank.rd_en == 1'h1) & (~cfg_pcfg_tile_connected_prev) & (~cfg_pcfg_tile_connected_next) & (rdrq_packet_pcfgdma2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_pcfgdma2bank.rd_addr[17] == 1'h1)) begin
    rdrq_packet_sw2bankarr_w[1].rd_en = rdrq_packet_pcfgdma2bank.rd_en;
    rdrq_packet_sw2bankarr_w[1].rd_addr = rdrq_packet_pcfgdma2bank.rd_addr[16:0];
    rd_type_1 = pcfg;
  end
  else if ((rdrq_packet_pcfgring2bank.rd_en == 1'h1) & (rdrq_packet_pcfgring2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_pcfgring2bank.rd_addr[17] == 1'h1)) begin
    rdrq_packet_sw2bankarr_w[1].rd_en = rdrq_packet_pcfgring2bank.rd_en;
    rdrq_packet_sw2bankarr_w[1].rd_addr = rdrq_packet_pcfgring2bank.rd_addr[16:0];
    rd_type_1 = pcfg;
  end
  else if ((rdrq_packet_dma2bank.rd_en == 1'h1) & (~cfg_tile_connected_prev) & (~cfg_tile_connected_next) & (rdrq_packet_dma2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_dma2bank.rd_addr[17] == 1'h1)) begin
    rdrq_packet_sw2bankarr_w[1].rd_en = rdrq_packet_dma2bank.rd_en;
    rdrq_packet_sw2bankarr_w[1].rd_addr = rdrq_packet_dma2bank.rd_addr[16:0];
    rd_type_1 = strm;
  end
  else if ((rdrq_packet_ring2bank.rd_en == 1'h1) & (rdrq_packet_ring2bank.rd_addr[18] == glb_tile_id) & (rdrq_packet_ring2bank.rd_addr[17] == 1'h1)) begin
    rdrq_packet_sw2bankarr_w[1].rd_en = rdrq_packet_ring2bank.rd_en;
    rdrq_packet_sw2bankarr_w[1].rd_addr = rdrq_packet_ring2bank.rd_addr[16:0];
    rd_type_1 = strm;
  end
  else begin
    rdrq_packet_sw2bankarr_w[1] = 18'h0;
    rd_type_1 = none;
  end
end
always_comb begin
  rdrs_packet_bank2dma = 65'h0;
  if ((~cfg_tile_connected_next) & (~cfg_tile_connected_prev)) begin
    if (rd_type_d_0 == strm) begin
      rdrs_packet_bank2dma = rdrs_packet_bankarr2sw_d[0];
    end
    if (rd_type_d_1 == strm) begin
      rdrs_packet_bank2dma = rdrs_packet_bankarr2sw_d[1];
    end
  end
end
always_comb begin
  rdrs_packet_bank2ring = 65'h0;
  if (cfg_tile_connected_next | cfg_tile_connected_prev) begin
    if (rd_type_d_0 == strm) begin
      rdrs_packet_bank2ring = rdrs_packet_bankarr2sw_d[0];
    end
    if (rd_type_d_1 == strm) begin
      rdrs_packet_bank2ring = rdrs_packet_bankarr2sw_d[1];
    end
  end
end
always_comb begin
  rdrs_packet_bank2procsw = 65'h0;
  if (rd_type_d_0 == proc) begin
    rdrs_packet_bank2procsw = rdrs_packet_bankarr2sw_d[0];
  end
  if (rd_type_d_1 == proc) begin
    rdrs_packet_bank2procsw = rdrs_packet_bankarr2sw_d[1];
  end
end
always_comb begin
  rdrs_packet_bank2pcfgdma = 65'h0;
  if ((~cfg_pcfg_tile_connected_next) & (~cfg_pcfg_tile_connected_prev)) begin
    if (rd_type_d_0 == pcfg) begin
      rdrs_packet_bank2pcfgdma = rdrs_packet_bankarr2sw_d[0];
    end
    if (rd_type_d_1 == pcfg) begin
      rdrs_packet_bank2pcfgdma = rdrs_packet_bankarr2sw_d[1];
    end
  end
end
always_comb begin
  rdrs_packet_bank2pcfgring = 65'h0;
  if (cfg_pcfg_tile_connected_next | cfg_pcfg_tile_connected_prev) begin
    if (rd_type_d_0 == pcfg) begin
      rdrs_packet_bank2pcfgring = rdrs_packet_bankarr2sw_d[0];
    end
    if (rd_type_d_1 == pcfg) begin
      rdrs_packet_bank2pcfgring = rdrs_packet_bankarr2sw_d[1];
    end
  end
end
pipeline_w_90_d_0 wr_sw2bank_pipeline_0 (
  .clk(clk),
  .clk_en(1'h1),
  .in_(wr_packet_sw2bankarr_w[0]),
  .reset(reset),
  .out_(wr_sw2bank_pipeline_0_out_)
);

pipeline_w_90_d_0 wr_sw2bank_pipeline_1 (
  .clk(clk),
  .clk_en(1'h1),
  .in_(wr_packet_sw2bankarr_w[1]),
  .reset(reset),
  .out_(wr_sw2bank_pipeline_1_out_)
);

pipeline_w_18_d_0 rdrq_sw2bank_pipeline_0 (
  .clk(clk),
  .clk_en(1'h1),
  .in_(rdrq_packet_sw2bankarr_w[0]),
  .reset(reset),
  .out_(rdrq_sw2bank_pipeline_0_out_)
);

pipeline_w_18_d_0 rdrq_sw2bank_pipeline_1 (
  .clk(clk),
  .clk_en(1'h1),
  .in_(rdrq_packet_sw2bankarr_w[1]),
  .reset(reset),
  .out_(rdrq_sw2bank_pipeline_1_out_)
);

pipeline_w_4_d_2 rd_type_pipeline_1 (
  .clk(clk),
  .clk_en(1'h1),
  .in_(rd_type_pipeline_1_in_),
  .reset(reset),
  .out_(rd_type_pipeline_1_out_)
);

pipeline_w_65_d_1 rdrs_bank2sw_pipeline_0 (
  .clk(clk),
  .clk_en(1'h1),
  .in_(rdrs_packet_bankarr2sw[0]),
  .reset(reset),
  .out_(rdrs_bank2sw_pipeline_0_out_)
);

pipeline_w_65_d_1 rdrs_bank2sw_pipeline_1 (
  .clk(clk),
  .clk_en(1'h1),
  .in_(rdrs_packet_bankarr2sw[1]),
  .reset(reset),
  .out_(rdrs_bank2sw_pipeline_1_out_)
);

endmodule   // glb_bank_mux

module glb_bank_sram_gen_14 (
  input logic [13:0] A,
  input logic [63:0] BW,
  input logic CEB,
  input logic CLK,
  input logic [63:0] D,
  input logic RESET,
  input logic WEB,
  output logic [63:0] Q
);

logic [11:0] A_SRAM;
logic [11:0] A_SRAM_d;
logic [63:0] BW_d;
logic [3:0] CEB_DEMUX;
logic [3:0] CEB_DEMUX_d;
logic CEB_d;
logic [63:0] D_d;
logic [1:0] Q_SEL;
logic [63:0] Q_SRAM2MUX [3:0];
logic [63:0] Q_w;
logic [1:0] SRAM_SEL;
logic [1:0] SRAM_SEL_d;
logic [3:0] WEB_DEMUX;
logic [3:0] WEB_DEMUX_d;
logic WEB_d;
logic [63:0] sram_array_0_Q;
logic [63:0] sram_array_1_Q;
logic [63:0] sram_array_2_Q;
logic [63:0] sram_array_3_Q;
logic [77:0] sram_signals_pipeline_in_;
logic [77:0] sram_signals_pipeline_out_;
logic [73:0] sram_signals_reset_high_pipeline_in_;
logic [73:0] sram_signals_reset_high_pipeline_out_;
assign SRAM_SEL = A[13:12];
assign A_SRAM = A[11:0];
assign sram_signals_reset_high_pipeline_in_ = {WEB, CEB, WEB_DEMUX, CEB_DEMUX, BW};
assign {WEB_d, CEB_d, WEB_DEMUX_d, CEB_DEMUX_d, BW_d} = sram_signals_reset_high_pipeline_out_;
assign sram_signals_pipeline_in_ = {A_SRAM, SRAM_SEL, D};
assign {A_SRAM_d, SRAM_SEL_d, D_d} = sram_signals_pipeline_out_;

always_ff @(posedge CLK, posedge RESET) begin
  if (RESET) begin
    Q_SEL <= 2'h0;
  end
  else if ((CEB_d == 1'h0) & (WEB_d == 1'h1)) begin
    Q_SEL <= SRAM_SEL_d;
  end
end
always_comb begin
  if (~WEB) begin
    WEB_DEMUX = ~(4'h1 << 4'(SRAM_SEL));
  end
  else WEB_DEMUX = 4'hF;
  if (~CEB) begin
    CEB_DEMUX = ~(4'h1 << 4'(SRAM_SEL));
  end
  else CEB_DEMUX = 4'hF;
end
assign Q_SRAM2MUX[0] = sram_array_0_Q;
assign Q_SRAM2MUX[1] = sram_array_1_Q;
assign Q_SRAM2MUX[2] = sram_array_2_Q;
assign Q_SRAM2MUX[3] = sram_array_3_Q;
assign Q_w = Q_SRAM2MUX[Q_SEL];
pipeline_w_74_d_0_reset_high sram_signals_reset_high_pipeline (
  .clk(CLK),
  .clk_en(1'h1),
  .in_(sram_signals_reset_high_pipeline_in_),
  .reset(RESET),
  .out_(sram_signals_reset_high_pipeline_out_)
);

pipeline_w_78_d_0 sram_signals_pipeline (
  .clk(CLK),
  .clk_en(1'h1),
  .in_(sram_signals_pipeline_in_),
  .reset(RESET),
  .out_(sram_signals_pipeline_out_)
);

pipeline_w_64_d_0 sram_signals_output_pipeline (
  .clk(CLK),
  .clk_en(1'h1),
  .in_(Q_w),
  .reset(RESET),
  .out_(Q)
);

IN12LP_S1DB_W04096B064M08S2_HB sram_array_0 (
  .A(A_SRAM_d),
  .BW(BW_d),
  .CEN(CEB_DEMUX_d[0]),
  .CLK(CLK),
  .D(D_d),
  .MA_SAWL0(1'h0),
  .MA_SAWL1(1'h0),
  .MA_STABAS0(1'h0),
  .MA_STABAS1(1'h0),
  .MA_VD0(1'h0),
  .MA_VD1(1'h0),
  .MA_WL0(1'h0),
  .MA_WL1(1'h0),
  .MA_WRAS0(1'h0),
  .MA_WRAS1(1'h0),
  .MA_WRT(1'h0),
  .RDWEN(WEB_DEMUX_d[0]),
  .T_LOGIC(1'h0),
  .T_Q_RST(1'h0),
  .Q(sram_array_0_Q)
);

IN12LP_S1DB_W04096B064M08S2_HB sram_array_1 (
  .A(A_SRAM_d),
  .BW(BW_d),
  .CEN(CEB_DEMUX_d[1]),
  .CLK(CLK),
  .D(D_d),
  .MA_SAWL0(1'h0),
  .MA_SAWL1(1'h0),
  .MA_STABAS0(1'h0),
  .MA_STABAS1(1'h0),
  .MA_VD0(1'h0),
  .MA_VD1(1'h0),
  .MA_WL0(1'h0),
  .MA_WL1(1'h0),
  .MA_WRAS0(1'h0),
  .MA_WRAS1(1'h0),
  .MA_WRT(1'h0),
  .RDWEN(WEB_DEMUX_d[1]),
  .T_LOGIC(1'h0),
  .T_Q_RST(1'h0),
  .Q(sram_array_1_Q)
);

IN12LP_S1DB_W04096B064M08S2_HB sram_array_2 (
  .A(A_SRAM_d),
  .BW(BW_d),
  .CEN(CEB_DEMUX_d[2]),
  .CLK(CLK),
  .D(D_d),
  .MA_SAWL0(1'h0),
  .MA_SAWL1(1'h0),
  .MA_STABAS0(1'h0),
  .MA_STABAS1(1'h0),
  .MA_VD0(1'h0),
  .MA_VD1(1'h0),
  .MA_WL0(1'h0),
  .MA_WL1(1'h0),
  .MA_WRAS0(1'h0),
  .MA_WRAS1(1'h0),
  .MA_WRT(1'h0),
  .RDWEN(WEB_DEMUX_d[2]),
  .T_LOGIC(1'h0),
  .T_Q_RST(1'h0),
  .Q(sram_array_2_Q)
);

IN12LP_S1DB_W04096B064M08S2_HB sram_array_3 (
  .A(A_SRAM_d),
  .BW(BW_d),
  .CEN(CEB_DEMUX_d[3]),
  .CLK(CLK),
  .D(D_d),
  .MA_SAWL0(1'h0),
  .MA_SAWL1(1'h0),
  .MA_STABAS0(1'h0),
  .MA_STABAS1(1'h0),
  .MA_VD0(1'h0),
  .MA_VD1(1'h0),
  .MA_WL0(1'h0),
  .MA_WL1(1'h0),
  .MA_WRAS0(1'h0),
  .MA_WRAS1(1'h0),
  .MA_WRT(1'h0),
  .RDWEN(WEB_DEMUX_d[3]),
  .T_LOGIC(1'h0),
  .T_Q_RST(1'h0),
  .Q(sram_array_3_Q)
);

endmodule   // glb_bank_sram_gen_14

module glb_cfg (
  glb_tile_ifc_A_12_D_32.master if_cfg_est_m,
  glb_tile_ifc_A_12_D_32.slave if_cfg_wst_s,
  input logic gclk,
  input logic glb_tile_id,
  input logic mclk,
  input logic reset,
  output cfg_data_network_t cfg_data_network,
  output load_dma_ctrl_t cfg_ld_dma_ctrl,
  output load_dma_header_t cfg_ld_dma_header,
  output pcfg_broadcast_mux_t cfg_pcfg_broadcast_mux,
  output pcfg_dma_ctrl_t cfg_pcfg_dma_ctrl,
  output pcfg_dma_header_t cfg_pcfg_dma_header,
  output cfg_pcfg_network_t cfg_pcfg_network,
  output store_dma_ctrl_t cfg_st_dma_ctrl,
  output store_dma_header_t cfg_st_dma_header,
  output logic [31:0] cfg_st_dma_num_blocks
);

logic [8:0] glb_cfg_ctrl_h2d_pio_dec_address;
logic glb_pio_d2h_dec_pio_ack;
logic glb_pio_d2h_dec_pio_nack;
logic [31:0] glb_pio_d2h_dec_pio_read_data;
logic [5:0] glb_pio_h2d_pio_dec_address;
logic glb_pio_h2d_pio_dec_read;
logic glb_pio_h2d_pio_dec_write;
logic [31:0] glb_pio_h2d_pio_dec_write_data;
logic glb_pio_l2h_data_network_ctrl_connected_r;
logic [5:0] glb_pio_l2h_data_network_latency_value_r;
logic [1:0] glb_pio_l2h_ld_dma_ctrl_data_mux_r;
logic glb_pio_l2h_ld_dma_ctrl_flush_mode_r;
logic [1:0] glb_pio_l2h_ld_dma_ctrl_mode_r;
logic glb_pio_l2h_ld_dma_ctrl_num_repeat_r;
logic [1:0] glb_pio_l2h_ld_dma_ctrl_valid_mode_r;
logic [15:0] glb_pio_l2h_ld_dma_header_0_cycle_start_addr_cycle_start_addr_r;
logic [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_0_cycle_stride_r;
logic [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_1_cycle_stride_r;
logic [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_2_cycle_stride_r;
logic [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_3_cycle_stride_r;
logic [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_4_cycle_stride_r;
logic [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_5_cycle_stride_r;
logic [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_6_cycle_stride_r;
logic [15:0] glb_pio_l2h_ld_dma_header_0_cycle_stride_7_cycle_stride_r;
logic [3:0] glb_pio_l2h_ld_dma_header_0_dim_dim_r;
logic [31:0] glb_pio_l2h_ld_dma_header_0_range_0_range_r;
logic [31:0] glb_pio_l2h_ld_dma_header_0_range_1_range_r;
logic [31:0] glb_pio_l2h_ld_dma_header_0_range_2_range_r;
logic [31:0] glb_pio_l2h_ld_dma_header_0_range_3_range_r;
logic [31:0] glb_pio_l2h_ld_dma_header_0_range_4_range_r;
logic [31:0] glb_pio_l2h_ld_dma_header_0_range_5_range_r;
logic [31:0] glb_pio_l2h_ld_dma_header_0_range_6_range_r;
logic [31:0] glb_pio_l2h_ld_dma_header_0_range_7_range_r;
logic [18:0] glb_pio_l2h_ld_dma_header_0_start_addr_start_addr_r;
logic [19:0] glb_pio_l2h_ld_dma_header_0_stride_0_stride_r;
logic [19:0] glb_pio_l2h_ld_dma_header_0_stride_1_stride_r;
logic [19:0] glb_pio_l2h_ld_dma_header_0_stride_2_stride_r;
logic [19:0] glb_pio_l2h_ld_dma_header_0_stride_3_stride_r;
logic [19:0] glb_pio_l2h_ld_dma_header_0_stride_4_stride_r;
logic [19:0] glb_pio_l2h_ld_dma_header_0_stride_5_stride_r;
logic [19:0] glb_pio_l2h_ld_dma_header_0_stride_6_stride_r;
logic [19:0] glb_pio_l2h_ld_dma_header_0_stride_7_stride_r;
logic [1:0] glb_pio_l2h_pcfg_broadcast_mux_east_r;
logic [1:0] glb_pio_l2h_pcfg_broadcast_mux_south_r;
logic [1:0] glb_pio_l2h_pcfg_broadcast_mux_west_r;
logic glb_pio_l2h_pcfg_dma_ctrl_mode_r;
logic glb_pio_l2h_pcfg_dma_ctrl_relocation_is_msb_r;
logic [15:0] glb_pio_l2h_pcfg_dma_ctrl_relocation_value_r;
logic [15:0] glb_pio_l2h_pcfg_dma_header_num_cfg_num_cfg_r;
logic [18:0] glb_pio_l2h_pcfg_dma_header_start_addr_start_addr_r;
logic glb_pio_l2h_pcfg_network_ctrl_connected_r;
logic [5:0] glb_pio_l2h_pcfg_network_latency_value_r;
logic [1:0] glb_pio_l2h_st_dma_ctrl_data_mux_r;
logic [1:0] glb_pio_l2h_st_dma_ctrl_mode_r;
logic glb_pio_l2h_st_dma_ctrl_num_repeat_r;
logic [1:0] glb_pio_l2h_st_dma_ctrl_valid_mode_r;
logic [15:0] glb_pio_l2h_st_dma_header_0_cycle_start_addr_cycle_start_addr_r;
logic [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_0_cycle_stride_r;
logic [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_1_cycle_stride_r;
logic [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_2_cycle_stride_r;
logic [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_3_cycle_stride_r;
logic [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_4_cycle_stride_r;
logic [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_5_cycle_stride_r;
logic [15:0] glb_pio_l2h_st_dma_header_0_cycle_stride_6_cycle_stride_r;
logic [3:0] glb_pio_l2h_st_dma_header_0_dim_dim_r;
logic [31:0] glb_pio_l2h_st_dma_header_0_range_0_range_r;
logic [31:0] glb_pio_l2h_st_dma_header_0_range_1_range_r;
logic [31:0] glb_pio_l2h_st_dma_header_0_range_2_range_r;
logic [31:0] glb_pio_l2h_st_dma_header_0_range_3_range_r;
logic [31:0] glb_pio_l2h_st_dma_header_0_range_4_range_r;
logic [31:0] glb_pio_l2h_st_dma_header_0_range_5_range_r;
logic [31:0] glb_pio_l2h_st_dma_header_0_range_6_range_r;
logic [18:0] glb_pio_l2h_st_dma_header_0_start_addr_start_addr_r;
logic [19:0] glb_pio_l2h_st_dma_header_0_stride_0_stride_r;
logic [19:0] glb_pio_l2h_st_dma_header_0_stride_1_stride_r;
logic [19:0] glb_pio_l2h_st_dma_header_0_stride_2_stride_r;
logic [19:0] glb_pio_l2h_st_dma_header_0_stride_3_stride_r;
logic [19:0] glb_pio_l2h_st_dma_header_0_stride_4_stride_r;
logic [19:0] glb_pio_l2h_st_dma_header_0_stride_5_stride_r;
logic [19:0] glb_pio_l2h_st_dma_header_0_stride_6_stride_r;
assign cfg_data_network.tile_connected = glb_pio_l2h_data_network_ctrl_connected_r;
assign cfg_data_network.latency = glb_pio_l2h_data_network_latency_value_r;
assign cfg_pcfg_network.tile_connected = glb_pio_l2h_pcfg_network_ctrl_connected_r;
assign cfg_pcfg_network.latency = glb_pio_l2h_pcfg_network_latency_value_r;
assign cfg_st_dma_ctrl.data_mux = glb_pio_l2h_st_dma_ctrl_data_mux_r;
assign cfg_st_dma_ctrl.mode = glb_pio_l2h_st_dma_ctrl_mode_r;
assign cfg_st_dma_ctrl.valid_mode = glb_pio_l2h_st_dma_ctrl_valid_mode_r;
assign cfg_st_dma_ctrl.num_repeat = glb_pio_l2h_st_dma_ctrl_num_repeat_r;
assign cfg_st_dma_header.start_addr = glb_pio_l2h_st_dma_header_0_start_addr_start_addr_r;
assign cfg_st_dma_header.cycle_start_addr = glb_pio_l2h_st_dma_header_0_cycle_start_addr_cycle_start_addr_r;
assign cfg_st_dma_header.dim = glb_pio_l2h_st_dma_header_0_dim_dim_r;
assign cfg_st_dma_header.cycle_stride_0 = glb_pio_l2h_st_dma_header_0_cycle_stride_0_cycle_stride_r;
assign cfg_st_dma_header.stride_0 = glb_pio_l2h_st_dma_header_0_stride_0_stride_r;
assign cfg_st_dma_header.range_0 = glb_pio_l2h_st_dma_header_0_range_0_range_r;
assign cfg_st_dma_header.cycle_stride_1 = glb_pio_l2h_st_dma_header_0_cycle_stride_1_cycle_stride_r;
assign cfg_st_dma_header.stride_1 = glb_pio_l2h_st_dma_header_0_stride_1_stride_r;
assign cfg_st_dma_header.range_1 = glb_pio_l2h_st_dma_header_0_range_1_range_r;
assign cfg_st_dma_header.cycle_stride_2 = glb_pio_l2h_st_dma_header_0_cycle_stride_2_cycle_stride_r;
assign cfg_st_dma_header.stride_2 = glb_pio_l2h_st_dma_header_0_stride_2_stride_r;
assign cfg_st_dma_header.range_2 = glb_pio_l2h_st_dma_header_0_range_2_range_r;
assign cfg_st_dma_header.cycle_stride_3 = glb_pio_l2h_st_dma_header_0_cycle_stride_3_cycle_stride_r;
assign cfg_st_dma_header.stride_3 = glb_pio_l2h_st_dma_header_0_stride_3_stride_r;
assign cfg_st_dma_header.range_3 = glb_pio_l2h_st_dma_header_0_range_3_range_r;
assign cfg_st_dma_header.cycle_stride_4 = glb_pio_l2h_st_dma_header_0_cycle_stride_4_cycle_stride_r;
assign cfg_st_dma_header.stride_4 = glb_pio_l2h_st_dma_header_0_stride_4_stride_r;
assign cfg_st_dma_header.range_4 = glb_pio_l2h_st_dma_header_0_range_4_range_r;
assign cfg_st_dma_header.cycle_stride_5 = glb_pio_l2h_st_dma_header_0_cycle_stride_5_cycle_stride_r;
assign cfg_st_dma_header.stride_5 = glb_pio_l2h_st_dma_header_0_stride_5_stride_r;
assign cfg_st_dma_header.range_5 = glb_pio_l2h_st_dma_header_0_range_5_range_r;
assign cfg_st_dma_header.cycle_stride_6 = glb_pio_l2h_st_dma_header_0_cycle_stride_6_cycle_stride_r;
assign cfg_st_dma_header.stride_6 = glb_pio_l2h_st_dma_header_0_stride_6_stride_r;
assign cfg_st_dma_header.range_6 = glb_pio_l2h_st_dma_header_0_range_6_range_r;
assign cfg_ld_dma_ctrl.data_mux = glb_pio_l2h_ld_dma_ctrl_data_mux_r;
assign cfg_ld_dma_ctrl.mode = glb_pio_l2h_ld_dma_ctrl_mode_r;
assign cfg_ld_dma_ctrl.valid_mode = glb_pio_l2h_ld_dma_ctrl_valid_mode_r;
assign cfg_ld_dma_ctrl.flush_mode = glb_pio_l2h_ld_dma_ctrl_flush_mode_r;
assign cfg_ld_dma_ctrl.num_repeat = glb_pio_l2h_ld_dma_ctrl_num_repeat_r;
assign cfg_ld_dma_header.start_addr = glb_pio_l2h_ld_dma_header_0_start_addr_start_addr_r;
assign cfg_ld_dma_header.cycle_start_addr = glb_pio_l2h_ld_dma_header_0_cycle_start_addr_cycle_start_addr_r;
assign cfg_ld_dma_header.dim = glb_pio_l2h_ld_dma_header_0_dim_dim_r;
assign cfg_ld_dma_header.cycle_stride_0 = glb_pio_l2h_ld_dma_header_0_cycle_stride_0_cycle_stride_r;
assign cfg_ld_dma_header.stride_0 = glb_pio_l2h_ld_dma_header_0_stride_0_stride_r;
assign cfg_ld_dma_header.range_0 = glb_pio_l2h_ld_dma_header_0_range_0_range_r;
assign cfg_ld_dma_header.cycle_stride_1 = glb_pio_l2h_ld_dma_header_0_cycle_stride_1_cycle_stride_r;
assign cfg_ld_dma_header.stride_1 = glb_pio_l2h_ld_dma_header_0_stride_1_stride_r;
assign cfg_ld_dma_header.range_1 = glb_pio_l2h_ld_dma_header_0_range_1_range_r;
assign cfg_ld_dma_header.cycle_stride_2 = glb_pio_l2h_ld_dma_header_0_cycle_stride_2_cycle_stride_r;
assign cfg_ld_dma_header.stride_2 = glb_pio_l2h_ld_dma_header_0_stride_2_stride_r;
assign cfg_ld_dma_header.range_2 = glb_pio_l2h_ld_dma_header_0_range_2_range_r;
assign cfg_ld_dma_header.cycle_stride_3 = glb_pio_l2h_ld_dma_header_0_cycle_stride_3_cycle_stride_r;
assign cfg_ld_dma_header.stride_3 = glb_pio_l2h_ld_dma_header_0_stride_3_stride_r;
assign cfg_ld_dma_header.range_3 = glb_pio_l2h_ld_dma_header_0_range_3_range_r;
assign cfg_ld_dma_header.cycle_stride_4 = glb_pio_l2h_ld_dma_header_0_cycle_stride_4_cycle_stride_r;
assign cfg_ld_dma_header.stride_4 = glb_pio_l2h_ld_dma_header_0_stride_4_stride_r;
assign cfg_ld_dma_header.range_4 = glb_pio_l2h_ld_dma_header_0_range_4_range_r;
assign cfg_ld_dma_header.cycle_stride_5 = glb_pio_l2h_ld_dma_header_0_cycle_stride_5_cycle_stride_r;
assign cfg_ld_dma_header.stride_5 = glb_pio_l2h_ld_dma_header_0_stride_5_stride_r;
assign cfg_ld_dma_header.range_5 = glb_pio_l2h_ld_dma_header_0_range_5_range_r;
assign cfg_ld_dma_header.cycle_stride_6 = glb_pio_l2h_ld_dma_header_0_cycle_stride_6_cycle_stride_r;
assign cfg_ld_dma_header.stride_6 = glb_pio_l2h_ld_dma_header_0_stride_6_stride_r;
assign cfg_ld_dma_header.range_6 = glb_pio_l2h_ld_dma_header_0_range_6_range_r;
assign cfg_ld_dma_header.cycle_stride_7 = glb_pio_l2h_ld_dma_header_0_cycle_stride_7_cycle_stride_r;
assign cfg_ld_dma_header.stride_7 = glb_pio_l2h_ld_dma_header_0_stride_7_stride_r;
assign cfg_ld_dma_header.range_7 = glb_pio_l2h_ld_dma_header_0_range_7_range_r;
assign cfg_pcfg_dma_ctrl.mode = glb_pio_l2h_pcfg_dma_ctrl_mode_r;
assign cfg_pcfg_dma_ctrl.relocation_value = glb_pio_l2h_pcfg_dma_ctrl_relocation_value_r;
assign cfg_pcfg_dma_ctrl.relocation_is_msb = glb_pio_l2h_pcfg_dma_ctrl_relocation_is_msb_r;
assign cfg_pcfg_dma_header.start_addr = glb_pio_l2h_pcfg_dma_header_start_addr_start_addr_r;
assign cfg_pcfg_dma_header.num_cfg = glb_pio_l2h_pcfg_dma_header_num_cfg_num_cfg_r;
assign cfg_pcfg_broadcast_mux.west = glb_pio_l2h_pcfg_broadcast_mux_west_r;
assign cfg_pcfg_broadcast_mux.east = glb_pio_l2h_pcfg_broadcast_mux_east_r;
assign cfg_pcfg_broadcast_mux.south = glb_pio_l2h_pcfg_broadcast_mux_south_r;
assign glb_pio_h2d_pio_dec_address = glb_cfg_ctrl_h2d_pio_dec_address[5:0];
glb_pio glb_pio (
  .clk(gclk),
  .h2d_pio_dec_address(glb_pio_h2d_pio_dec_address),
  .h2d_pio_dec_read(glb_pio_h2d_pio_dec_read),
  .h2d_pio_dec_write(glb_pio_h2d_pio_dec_write),
  .h2d_pio_dec_write_data(glb_pio_h2d_pio_dec_write_data),
  .reset(reset),
  .d2h_dec_pio_ack(glb_pio_d2h_dec_pio_ack),
  .d2h_dec_pio_nack(glb_pio_d2h_dec_pio_nack),
  .d2h_dec_pio_read_data(glb_pio_d2h_dec_pio_read_data),
  .l2h_data_network_ctrl_connected_r(glb_pio_l2h_data_network_ctrl_connected_r),
  .l2h_data_network_latency_value_r(glb_pio_l2h_data_network_latency_value_r),
  .l2h_ld_dma_ctrl_data_mux_r(glb_pio_l2h_ld_dma_ctrl_data_mux_r),
  .l2h_ld_dma_ctrl_flush_mode_r(glb_pio_l2h_ld_dma_ctrl_flush_mode_r),
  .l2h_ld_dma_ctrl_mode_r(glb_pio_l2h_ld_dma_ctrl_mode_r),
  .l2h_ld_dma_ctrl_num_repeat_r(glb_pio_l2h_ld_dma_ctrl_num_repeat_r),
  .l2h_ld_dma_ctrl_valid_mode_r(glb_pio_l2h_ld_dma_ctrl_valid_mode_r),
  .l2h_ld_dma_header_0_cycle_start_addr_cycle_start_addr_r(glb_pio_l2h_ld_dma_header_0_cycle_start_addr_cycle_start_addr_r),
  .l2h_ld_dma_header_0_cycle_stride_0_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_0_cycle_stride_r),
  .l2h_ld_dma_header_0_cycle_stride_1_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_1_cycle_stride_r),
  .l2h_ld_dma_header_0_cycle_stride_2_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_2_cycle_stride_r),
  .l2h_ld_dma_header_0_cycle_stride_3_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_3_cycle_stride_r),
  .l2h_ld_dma_header_0_cycle_stride_4_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_4_cycle_stride_r),
  .l2h_ld_dma_header_0_cycle_stride_5_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_5_cycle_stride_r),
  .l2h_ld_dma_header_0_cycle_stride_6_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_6_cycle_stride_r),
  .l2h_ld_dma_header_0_cycle_stride_7_cycle_stride_r(glb_pio_l2h_ld_dma_header_0_cycle_stride_7_cycle_stride_r),
  .l2h_ld_dma_header_0_dim_dim_r(glb_pio_l2h_ld_dma_header_0_dim_dim_r),
  .l2h_ld_dma_header_0_range_0_range_r(glb_pio_l2h_ld_dma_header_0_range_0_range_r),
  .l2h_ld_dma_header_0_range_1_range_r(glb_pio_l2h_ld_dma_header_0_range_1_range_r),
  .l2h_ld_dma_header_0_range_2_range_r(glb_pio_l2h_ld_dma_header_0_range_2_range_r),
  .l2h_ld_dma_header_0_range_3_range_r(glb_pio_l2h_ld_dma_header_0_range_3_range_r),
  .l2h_ld_dma_header_0_range_4_range_r(glb_pio_l2h_ld_dma_header_0_range_4_range_r),
  .l2h_ld_dma_header_0_range_5_range_r(glb_pio_l2h_ld_dma_header_0_range_5_range_r),
  .l2h_ld_dma_header_0_range_6_range_r(glb_pio_l2h_ld_dma_header_0_range_6_range_r),
  .l2h_ld_dma_header_0_range_7_range_r(glb_pio_l2h_ld_dma_header_0_range_7_range_r),
  .l2h_ld_dma_header_0_start_addr_start_addr_r(glb_pio_l2h_ld_dma_header_0_start_addr_start_addr_r),
  .l2h_ld_dma_header_0_stride_0_stride_r(glb_pio_l2h_ld_dma_header_0_stride_0_stride_r),
  .l2h_ld_dma_header_0_stride_1_stride_r(glb_pio_l2h_ld_dma_header_0_stride_1_stride_r),
  .l2h_ld_dma_header_0_stride_2_stride_r(glb_pio_l2h_ld_dma_header_0_stride_2_stride_r),
  .l2h_ld_dma_header_0_stride_3_stride_r(glb_pio_l2h_ld_dma_header_0_stride_3_stride_r),
  .l2h_ld_dma_header_0_stride_4_stride_r(glb_pio_l2h_ld_dma_header_0_stride_4_stride_r),
  .l2h_ld_dma_header_0_stride_5_stride_r(glb_pio_l2h_ld_dma_header_0_stride_5_stride_r),
  .l2h_ld_dma_header_0_stride_6_stride_r(glb_pio_l2h_ld_dma_header_0_stride_6_stride_r),
  .l2h_ld_dma_header_0_stride_7_stride_r(glb_pio_l2h_ld_dma_header_0_stride_7_stride_r),
  .l2h_pcfg_broadcast_mux_east_r(glb_pio_l2h_pcfg_broadcast_mux_east_r),
  .l2h_pcfg_broadcast_mux_south_r(glb_pio_l2h_pcfg_broadcast_mux_south_r),
  .l2h_pcfg_broadcast_mux_west_r(glb_pio_l2h_pcfg_broadcast_mux_west_r),
  .l2h_pcfg_dma_ctrl_mode_r(glb_pio_l2h_pcfg_dma_ctrl_mode_r),
  .l2h_pcfg_dma_ctrl_relocation_is_msb_r(glb_pio_l2h_pcfg_dma_ctrl_relocation_is_msb_r),
  .l2h_pcfg_dma_ctrl_relocation_value_r(glb_pio_l2h_pcfg_dma_ctrl_relocation_value_r),
  .l2h_pcfg_dma_header_num_cfg_num_cfg_r(glb_pio_l2h_pcfg_dma_header_num_cfg_num_cfg_r),
  .l2h_pcfg_dma_header_start_addr_start_addr_r(glb_pio_l2h_pcfg_dma_header_start_addr_start_addr_r),
  .l2h_pcfg_network_ctrl_connected_r(glb_pio_l2h_pcfg_network_ctrl_connected_r),
  .l2h_pcfg_network_latency_value_r(glb_pio_l2h_pcfg_network_latency_value_r),
  .l2h_st_dma_ctrl_data_mux_r(glb_pio_l2h_st_dma_ctrl_data_mux_r),
  .l2h_st_dma_ctrl_mode_r(glb_pio_l2h_st_dma_ctrl_mode_r),
  .l2h_st_dma_ctrl_num_repeat_r(glb_pio_l2h_st_dma_ctrl_num_repeat_r),
  .l2h_st_dma_ctrl_valid_mode_r(glb_pio_l2h_st_dma_ctrl_valid_mode_r),
  .l2h_st_dma_header_0_cycle_start_addr_cycle_start_addr_r(glb_pio_l2h_st_dma_header_0_cycle_start_addr_cycle_start_addr_r),
  .l2h_st_dma_header_0_cycle_stride_0_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_0_cycle_stride_r),
  .l2h_st_dma_header_0_cycle_stride_1_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_1_cycle_stride_r),
  .l2h_st_dma_header_0_cycle_stride_2_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_2_cycle_stride_r),
  .l2h_st_dma_header_0_cycle_stride_3_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_3_cycle_stride_r),
  .l2h_st_dma_header_0_cycle_stride_4_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_4_cycle_stride_r),
  .l2h_st_dma_header_0_cycle_stride_5_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_5_cycle_stride_r),
  .l2h_st_dma_header_0_cycle_stride_6_cycle_stride_r(glb_pio_l2h_st_dma_header_0_cycle_stride_6_cycle_stride_r),
  .l2h_st_dma_header_0_dim_dim_r(glb_pio_l2h_st_dma_header_0_dim_dim_r),
  .l2h_st_dma_header_0_range_0_range_r(glb_pio_l2h_st_dma_header_0_range_0_range_r),
  .l2h_st_dma_header_0_range_1_range_r(glb_pio_l2h_st_dma_header_0_range_1_range_r),
  .l2h_st_dma_header_0_range_2_range_r(glb_pio_l2h_st_dma_header_0_range_2_range_r),
  .l2h_st_dma_header_0_range_3_range_r(glb_pio_l2h_st_dma_header_0_range_3_range_r),
  .l2h_st_dma_header_0_range_4_range_r(glb_pio_l2h_st_dma_header_0_range_4_range_r),
  .l2h_st_dma_header_0_range_5_range_r(glb_pio_l2h_st_dma_header_0_range_5_range_r),
  .l2h_st_dma_header_0_range_6_range_r(glb_pio_l2h_st_dma_header_0_range_6_range_r),
  .l2h_st_dma_header_0_start_addr_start_addr_r(glb_pio_l2h_st_dma_header_0_start_addr_start_addr_r),
  .l2h_st_dma_header_0_stride_0_stride_r(glb_pio_l2h_st_dma_header_0_stride_0_stride_r),
  .l2h_st_dma_header_0_stride_1_stride_r(glb_pio_l2h_st_dma_header_0_stride_1_stride_r),
  .l2h_st_dma_header_0_stride_2_stride_r(glb_pio_l2h_st_dma_header_0_stride_2_stride_r),
  .l2h_st_dma_header_0_stride_3_stride_r(glb_pio_l2h_st_dma_header_0_stride_3_stride_r),
  .l2h_st_dma_header_0_stride_4_stride_r(glb_pio_l2h_st_dma_header_0_stride_4_stride_r),
  .l2h_st_dma_header_0_stride_5_stride_r(glb_pio_l2h_st_dma_header_0_stride_5_stride_r),
  .l2h_st_dma_header_0_stride_6_stride_r(glb_pio_l2h_st_dma_header_0_stride_6_stride_r),
  .l2h_st_dma_num_blocks_value_r(cfg_st_dma_num_blocks)
);

glb_cfg_ctrl glb_cfg_ctrl (
  .d2h_dec_pio_ack(glb_pio_d2h_dec_pio_ack),
  .d2h_dec_pio_nack(glb_pio_d2h_dec_pio_nack),
  .d2h_dec_pio_read_data(glb_pio_d2h_dec_pio_read_data),
  .gclk(gclk),
  .glb_tile_id(glb_tile_id),
  .mclk(mclk),
  .if_cfg_wst_s(if_cfg_wst_s),
  .if_cfg_est_m(if_cfg_est_m),
  .reset(reset),
  .h2d_pio_dec_address(glb_cfg_ctrl_h2d_pio_dec_address),
  .h2d_pio_dec_read(glb_pio_h2d_pio_dec_read),
  .h2d_pio_dec_write(glb_pio_h2d_pio_dec_write),
  .h2d_pio_dec_write_data(glb_pio_h2d_pio_dec_write_data)
);

endmodule   // glb_cfg

module glb_cfg_ctrl (
  glb_tile_ifc_A_12_D_32.master if_cfg_est_m,
  glb_tile_ifc_A_12_D_32.slave if_cfg_wst_s,
  input logic d2h_dec_pio_ack,
  input logic d2h_dec_pio_nack,
  input logic [31:0] d2h_dec_pio_read_data,
  input logic gclk,
  input logic glb_tile_id,
  input logic mclk,
  input logic reset,
  output logic [8:0] h2d_pio_dec_address,
  output logic h2d_pio_dec_read,
  output logic h2d_pio_dec_write,
  output logic [31:0] h2d_pio_dec_write_data
);

logic [8:0] addr_internal;
logic if_cfg_est_m_rd_clk_en_sel;
logic if_cfg_est_m_rd_clk_en_sel_first_cycle;
logic if_cfg_est_m_rd_clk_en_sel_latch;
logic if_cfg_est_m_wr_clk_en_sel;
logic if_cfg_est_m_wr_clk_en_sel_first_cycle;
logic if_cfg_est_m_wr_clk_en_sel_latch;
logic if_cfg_wst_s_rd_clk_en_d;
logic if_cfg_wst_s_wr_clk_en_d;
logic [31:0] rd_data_internal;
logic rd_data_valid_internal;
logic rd_en_d1;
logic rd_en_d2;
logic rd_tile_id_match;
logic read_internal;
logic [31:0] wr_data_internal;
logic wr_tile_id_match;
logic write_internal;
always_comb begin
  wr_tile_id_match = glb_tile_id == if_cfg_wst_s.wr_addr[11];
  rd_tile_id_match = glb_tile_id == if_cfg_wst_s.rd_addr[11];
end
always_comb begin
  wr_data_internal = 32'h0;
  addr_internal = 9'h0;
  read_internal = 1'h0;
  write_internal = 1'h0;
  if (if_cfg_wst_s.rd_en && rd_tile_id_match) begin
    addr_internal = if_cfg_wst_s.rd_addr[10:2];
    read_internal = 1'h1;
  end
  if (if_cfg_wst_s.wr_en && wr_tile_id_match) begin
    addr_internal = if_cfg_wst_s.wr_addr[10:2];
    wr_data_internal = if_cfg_wst_s.wr_data;
    write_internal = 1'h1;
  end
end

always_ff @(posedge gclk, posedge reset) begin
  if (reset) begin
    if_cfg_est_m.wr_en <= 1'h0;
    if_cfg_est_m.wr_addr <= 12'h0;
    if_cfg_est_m.wr_data <= 32'h0;
  end
  else if (~(wr_tile_id_match && (if_cfg_wst_s.wr_en == 1'h1))) begin
    if_cfg_est_m.wr_en <= if_cfg_wst_s.wr_en;
    if_cfg_est_m.wr_addr <= if_cfg_wst_s.wr_addr;
    if_cfg_est_m.wr_data <= if_cfg_wst_s.wr_data;
  end
  else begin
    if_cfg_est_m.wr_en <= 1'h0;
    if_cfg_est_m.wr_addr <= 12'h0;
    if_cfg_est_m.wr_data <= 32'h0;
  end
end

always_ff @(posedge gclk, posedge reset) begin
  if (reset) begin
    if_cfg_est_m.rd_en <= 1'h0;
    if_cfg_est_m.rd_addr <= 12'h0;
  end
  else if (~(rd_tile_id_match && (if_cfg_wst_s.rd_en == 1'h1))) begin
    if_cfg_est_m.rd_en <= if_cfg_wst_s.rd_en;
    if_cfg_est_m.rd_addr <= if_cfg_wst_s.rd_addr;
  end
  else begin
    if_cfg_est_m.rd_en <= 1'h0;
    if_cfg_est_m.rd_addr <= 12'h0;
  end
end

always_ff @(posedge gclk, posedge reset) begin
  if (reset) begin
    if_cfg_wst_s.rd_data <= 32'h0;
    if_cfg_wst_s.rd_data_valid <= 1'h0;
  end
  else if (rd_data_valid_internal) begin
    if_cfg_wst_s.rd_data <= rd_data_internal;
    if_cfg_wst_s.rd_data_valid <= rd_data_valid_internal;
  end
  else begin
    if_cfg_wst_s.rd_data <= if_cfg_est_m.rd_data;
    if_cfg_wst_s.rd_data_valid <= if_cfg_est_m.rd_data_valid;
  end
end

always_ff @(posedge gclk, posedge reset) begin
  if (reset) begin
    rd_en_d1 <= 1'h0;
    rd_en_d2 <= 1'h0;
  end
  else begin
    rd_en_d1 <= read_internal;
    rd_en_d2 <= rd_en_d1;
  end
end

always_ff @(posedge gclk, posedge reset) begin
  if (reset) begin
    rd_data_valid_internal <= 1'h0;
    rd_data_internal <= 32'h0;
  end
  else if ((rd_en_d2 == 1'h1) & (d2h_dec_pio_ack | d2h_dec_pio_nack)) begin
    rd_data_valid_internal <= 1'h1;
    rd_data_internal <= d2h_dec_pio_read_data;
  end
  else begin
    rd_data_valid_internal <= 1'h0;
    rd_data_internal <= 32'h0;
  end
end

always_ff @(posedge mclk, posedge reset) begin
  if (reset) begin
    if_cfg_wst_s_wr_clk_en_d <= 1'h0;
    if_cfg_wst_s_rd_clk_en_d <= 1'h0;
  end
  else begin
    if_cfg_wst_s_wr_clk_en_d <= if_cfg_wst_s.wr_clk_en;
    if_cfg_wst_s_rd_clk_en_d <= if_cfg_wst_s.rd_clk_en;
  end
end
always_comb begin
  if_cfg_est_m_wr_clk_en_sel_first_cycle = if_cfg_wst_s.wr_en & (~wr_tile_id_match);
  if_cfg_est_m_rd_clk_en_sel_first_cycle = if_cfg_wst_s.rd_en & (~rd_tile_id_match);
end

always_ff @(posedge mclk, posedge reset) begin
  if (reset) begin
    if_cfg_est_m_wr_clk_en_sel_latch <= 1'h0;
  end
  else if (if_cfg_wst_s.wr_en == 1'h1) begin
    if (wr_tile_id_match) begin
      if_cfg_est_m_wr_clk_en_sel_latch <= 1'h0;
    end
    else if_cfg_est_m_wr_clk_en_sel_latch <= 1'h1;
  end
  else if (if_cfg_wst_s.wr_clk_en == 1'h0) begin
    if_cfg_est_m_wr_clk_en_sel_latch <= 1'h0;
  end
end

always_ff @(posedge mclk, posedge reset) begin
  if (reset) begin
    if_cfg_est_m_rd_clk_en_sel_latch <= 1'h0;
  end
  else if (if_cfg_wst_s.rd_en == 1'h1) begin
    if (rd_tile_id_match) begin
      if_cfg_est_m_rd_clk_en_sel_latch <= 1'h0;
    end
    else if_cfg_est_m_rd_clk_en_sel_latch <= 1'h1;
  end
  else if (if_cfg_wst_s.rd_clk_en == 1'h0) begin
    if_cfg_est_m_rd_clk_en_sel_latch <= 1'h0;
  end
end
always_comb begin
  if_cfg_est_m_wr_clk_en_sel = if_cfg_est_m_wr_clk_en_sel_first_cycle | if_cfg_est_m_wr_clk_en_sel_latch;
  if_cfg_est_m_rd_clk_en_sel = if_cfg_est_m_rd_clk_en_sel_first_cycle | if_cfg_est_m_rd_clk_en_sel_latch;
end
always_comb begin
  if (if_cfg_est_m_wr_clk_en_sel) begin
    if_cfg_est_m.wr_clk_en = if_cfg_wst_s_wr_clk_en_d;
  end
  else if_cfg_est_m.wr_clk_en = 1'h0;
end
always_comb begin
  if (if_cfg_est_m_rd_clk_en_sel) begin
    if_cfg_est_m.rd_clk_en = if_cfg_wst_s_rd_clk_en_d;
  end
  else if_cfg_est_m.rd_clk_en = 1'h0;
end
assign h2d_pio_dec_write_data = wr_data_internal;
assign h2d_pio_dec_address = addr_internal;
assign h2d_pio_dec_read = read_internal;
assign h2d_pio_dec_write = write_internal;
endmodule   // glb_cfg_ctrl

module glb_clk_en_gen_11 #(
  parameter cnt = 32'hB
)
(
  input logic clk,
  input logic enable,
  input logic reset,
  output logic clk_en
);

logic [31:0] clk_en_cnt;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    clk_en_cnt <= 32'h0;
  end
  else if (enable) begin
    clk_en_cnt <= cnt - 32'h1;
  end
  else if (clk_en_cnt > 32'h0) begin
    clk_en_cnt <= clk_en_cnt - 32'h1;
  end
end
assign clk_en = enable | (clk_en_cnt > 32'h0);
endmodule   // glb_clk_en_gen_11

module glb_clk_en_gen_4 #(
  parameter cnt = 32'h4
)
(
  input logic clk,
  input logic enable,
  input logic reset,
  output logic clk_en
);

logic [31:0] clk_en_cnt;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    clk_en_cnt <= 32'h0;
  end
  else if (enable) begin
    clk_en_cnt <= cnt - 32'h1;
  end
  else if (clk_en_cnt > 32'h0) begin
    clk_en_cnt <= clk_en_cnt - 32'h1;
  end
end
assign clk_en = enable | (clk_en_cnt > 32'h0);
endmodule   // glb_clk_en_gen_4

module glb_clk_en_gen_5 #(
  parameter cnt = 32'h5
)
(
  input logic clk,
  input logic enable,
  input logic reset,
  output logic clk_en
);

logic [31:0] clk_en_cnt;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    clk_en_cnt <= 32'h0;
  end
  else if (enable) begin
    clk_en_cnt <= cnt - 32'h1;
  end
  else if (clk_en_cnt > 32'h0) begin
    clk_en_cnt <= clk_en_cnt - 32'h1;
  end
end
assign clk_en = enable | (clk_en_cnt > 32'h0);
endmodule   // glb_clk_en_gen_5

module glb_clk_en_gen_6 #(
  parameter cnt = 32'h6
)
(
  input logic clk,
  input logic enable,
  input logic reset,
  output logic clk_en
);

logic [31:0] clk_en_cnt;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    clk_en_cnt <= 32'h0;
  end
  else if (enable) begin
    clk_en_cnt <= cnt - 32'h1;
  end
  else if (clk_en_cnt > 32'h0) begin
    clk_en_cnt <= clk_en_cnt - 32'h1;
  end
end
assign clk_en = enable | (clk_en_cnt > 32'h0);
endmodule   // glb_clk_en_gen_6

module glb_crossbar_I_2_O_1_W_1 (
  input logic [1:0] in_,
  input logic sel_,
  output logic out_
);

always_comb begin
  out_ = in_[sel_];
end
endmodule   // glb_crossbar_I_2_O_1_W_1

module glb_load_dma (
  input logic [1:0] cfg_data_network_g2f_mux,
  input logic [5:0] cfg_data_network_latency,
  input logic cfg_ld_dma_ctrl_flush_mode,
  input logic [1:0] cfg_ld_dma_ctrl_mode,
  input logic [1:0] cfg_ld_dma_ctrl_valid_mode,
  input load_dma_header_t cfg_ld_dma_header,
  input logic cfg_ld_dma_num_repeat,
  input logic cfg_tile_connected_next,
  input logic cfg_tile_connected_prev,
  input logic clk,
  input logic [1:0] data_g2f_rdy,
  input logic glb_tile_id,
  input logic ld_dma_start_pulse,
  input rdrs_packet_t rdrs_packet_bank2dma,
  input rdrs_packet_t rdrs_packet_ring2dma,
  input logic reset,
  output logic clk_en_dma2bank,
  output logic [1:0] ctrl_g2f,
  output logic data_flush,
  output logic [1:0] [15:0] data_g2f,
  output logic [1:0] data_g2f_vld,
  output logic ld_dma_done_interrupt,
  output rdrq_packet_t rdrq_packet_dma2bank,
  output rdrq_packet_t rdrq_packet_dma2ring
);

logic all_skid_empty;
logic [18:0] bank_rdrq_rd_addr;
logic bank_rdrq_rd_en;
logic [63:0] bank_rdrs_data_cache_r;
logic [1:0] ctrl_g2f_w;
load_dma_header_t current_dma_header;
logic [15:0] cycle_count;
logic cycle_counter_en;
logic [15:0] cycle_current_addr;
logic [7:0][15:0] cycle_stride_addr_gen_strides;
logic cycle_valid;
logic [19:0] data_current_addr;
logic [15:0] data_dma2fifo;
logic [15:0] data_fifo2cgra;
logic data_flush_w;
logic [1:0] data_g2f_rdy_muxed;
logic [15:0] data_g2f_skid_0_data_out;
logic data_g2f_skid_0_empty;
logic data_g2f_skid_0_full;
logic [15:0] data_g2f_skid_1_data_out;
logic data_g2f_skid_1_empty;
logic data_g2f_skid_1_full;
logic [19:0] data_stride_addr_gen_start_addr;
logic [7:0][19:0] data_stride_addr_gen_strides;
logic dma2bank_clk_en;
logic [1:0] fifo2skid_rdy;
logic fifo2skid_rdy_muxed;
logic [1:0] fifo2skid_vld;
logic fifo2skid_vld_muxed;
logic fifo_almost_full;
logic [4:0] fifo_almost_full_diff;
logic fifo_empty;
logic fifo_full;
logic fifo_pop;
logic fifo_push;
logic fifo_push_ready;
logic is_cached;
logic is_first;
logic iter_step_valid;
logic [18:0] last_strm_rd_addr_r;
logic ld_dma_done_pulse;
logic ld_dma_done_pulse_anded;
logic ld_dma_done_pulse_d_arr [23:0];
logic ld_dma_done_pulse_last;
logic ld_dma_done_pulse_latch;
logic ld_dma_done_pulse_pipeline_out;
logic ld_dma_done_pulse_w;
logic ld_dma_start_pulse_next;
logic ld_dma_start_pulse_r;
logic loop_done;
logic [7:0][31:0] loop_iter_ranges;
logic [2:0] loop_mux_sel;
logic [1:0] pipeline_ctrl_in;
logic [1:0] pipeline_ctrl_out;
rdrq_packet_t rdrq_packet_dma2bank_w;
rdrq_packet_t rdrq_packet_dma2ring_w;
rdrs_packet_t rdrs_packet;
logic repeat_cnt;
logic [1:0] skid_empty;
logic [1:0] skid_full;
logic [1:0][15:0] skid_in;
logic [1:0][15:0] skid_out;
logic [1:0] skid_pop;
logic [1:0] skid_push;
logic strm_ctrl_muxed;
logic [15:0] strm_data;
logic [1:0] strm_data_sel_arr [21:0];
logic [1:0] strm_data_sel_w;
logic strm_data_start_pulse;
logic strm_data_start_pulse_d_arr [21:0];
logic strm_data_valid;
logic [18:0] strm_rd_addr_w;
logic strm_rd_en_d_arr [21:0];
logic strm_rd_en_w;
logic strm_run;
assign fifo_push_ready = ~fifo_almost_full;
assign data_dma2fifo = strm_data;
assign fifo_push = (~fifo_full) & strm_data_valid;
assign fifo2skid_vld_muxed = ~fifo_empty;
assign fifo_pop = fifo2skid_vld_muxed & fifo2skid_rdy_muxed;
always_comb begin
  fifo_almost_full_diff = 5'(6'h5 + cfg_data_network_latency);
end
assign skid_out[0] = data_g2f_skid_0_data_out;
assign skid_full[0] = data_g2f_skid_0_full;
assign skid_empty[0] = data_g2f_skid_0_empty;
assign data_g2f[0] = skid_out[0];
assign fifo2skid_rdy[0] = ~skid_full[0];
assign skid_push[0] = fifo2skid_rdy[0] & fifo2skid_vld[0];
assign data_g2f_vld[0] = ~skid_empty[0];
assign skid_pop[0] = (~skid_empty[0]) & data_g2f_rdy_muxed[0];
assign skid_out[1] = data_g2f_skid_1_data_out;
assign skid_full[1] = data_g2f_skid_1_full;
assign skid_empty[1] = data_g2f_skid_1_empty;
assign data_g2f[1] = skid_out[1];
assign fifo2skid_rdy[1] = ~skid_full[1];
assign skid_push[1] = fifo2skid_rdy[1] & fifo2skid_vld[1];
assign data_g2f_vld[1] = ~skid_empty[1];
assign skid_pop[1] = (~skid_empty[1]) & data_g2f_rdy_muxed[1];
always_comb begin
  fifo2skid_rdy_muxed = 1'h0;
  if (cfg_data_network_g2f_mux[0] == 1'h1) begin
    fifo2skid_rdy_muxed = fifo2skid_rdy[0];
    fifo2skid_vld[0] = fifo2skid_vld_muxed;
    skid_in[0] = data_fifo2cgra;
  end
  else begin
    fifo2skid_rdy_muxed = fifo2skid_rdy_muxed;
    fifo2skid_vld[0] = 1'h0;
    skid_in[0] = 16'h0;
  end
  if (cfg_data_network_g2f_mux[1] == 1'h1) begin
    fifo2skid_rdy_muxed = fifo2skid_rdy[1];
    fifo2skid_vld[1] = fifo2skid_vld_muxed;
    skid_in[1] = data_fifo2cgra;
  end
  else begin
    fifo2skid_rdy_muxed = fifo2skid_rdy_muxed;
    fifo2skid_vld[1] = 1'h0;
    skid_in[1] = 16'h0;
  end
end
always_comb begin
  if (cfg_ld_dma_ctrl_valid_mode == 2'h2) begin
    data_g2f_rdy_muxed[0] = data_g2f_rdy[0];
  end
  else data_g2f_rdy_muxed[0] = 1'h1;
  if (cfg_ld_dma_ctrl_valid_mode == 2'h2) begin
    data_g2f_rdy_muxed[1] = data_g2f_rdy[1];
  end
  else data_g2f_rdy_muxed[1] = 1'h1;
end
always_comb begin
  all_skid_empty = 1'h1;
  if (cfg_data_network_g2f_mux[0]) begin
    all_skid_empty = all_skid_empty & skid_empty[0];
  end
  else all_skid_empty = all_skid_empty;
  if (cfg_data_network_g2f_mux[1]) begin
    all_skid_empty = all_skid_empty & skid_empty[1];
  end
  else all_skid_empty = all_skid_empty;
end
assign current_dma_header = cfg_ld_dma_header;
always_comb begin
  if (cycle_counter_en) begin
    iter_step_valid = cycle_valid;
  end
  else iter_step_valid = strm_run & fifo_push_ready;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    repeat_cnt <= 1'h0;
  end
  else if (cfg_ld_dma_ctrl_mode == 2'h2) begin
    if (ld_dma_done_pulse) begin
      if ((repeat_cnt + 1'h1) < cfg_ld_dma_num_repeat) begin
        repeat_cnt <= repeat_cnt + 1'h1;
      end
    end
  end
  else if (cfg_ld_dma_ctrl_mode == 2'h3) begin
    if (ld_dma_done_pulse) begin
      if (((repeat_cnt + 1'h1) < cfg_ld_dma_num_repeat) & ((repeat_cnt + 1'h1) < 1'h1)) begin
        repeat_cnt <= repeat_cnt + 1'h1;
      end
    end
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    cycle_count <= 16'h0;
  end
  else if (ld_dma_start_pulse_r) begin
    cycle_count <= 16'h0;
  end
  else if (loop_done) begin
    cycle_count <= 16'h0;
  end
  else if (cycle_counter_en & strm_run) begin
    cycle_count <= cycle_count + 16'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    is_first <= 1'h0;
  end
  else if (ld_dma_start_pulse_r) begin
    is_first <= 1'h1;
  end
  else if (bank_rdrq_rd_en) begin
    is_first <= 1'h0;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    strm_run <= 1'h0;
  end
  else if (ld_dma_start_pulse_r) begin
    strm_run <= 1'h1;
  end
  else if (loop_done) begin
    strm_run <= 1'h0;
  end
end
assign strm_data_start_pulse = strm_data_start_pulse_d_arr[5'(cfg_data_network_latency) + 5'h3];
assign strm_data_valid = strm_rd_en_d_arr[5'(cfg_data_network_latency) + 5'h3];
assign strm_data_sel_w = strm_rd_addr_w[2:1];
always_comb begin
  if (cfg_ld_dma_ctrl_mode == 2'h0) begin
    ld_dma_start_pulse_next = 1'h0;
  end
  else if (cfg_ld_dma_ctrl_mode == 2'h1) begin
    ld_dma_start_pulse_next = (~strm_run) & ld_dma_start_pulse;
  end
  else if ((cfg_ld_dma_ctrl_mode == 2'h2) | (cfg_ld_dma_ctrl_mode == 2'h3)) begin
    ld_dma_start_pulse_next = ((~strm_run) & ld_dma_start_pulse) | (ld_dma_done_pulse & ((repeat_cnt + 1'h1) <
        cfg_ld_dma_num_repeat));
  end
  else ld_dma_start_pulse_next = 1'h0;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    ld_dma_start_pulse_r <= 1'h0;
  end
  else if (ld_dma_start_pulse_r) begin
    ld_dma_start_pulse_r <= 1'h0;
  end
  else ld_dma_start_pulse_r <= ld_dma_start_pulse_next;
end
always_comb begin
  if (cfg_ld_dma_ctrl_flush_mode == 1'h0) begin
    data_flush_w = strm_data_start_pulse;
    if (cfg_ld_dma_ctrl_valid_mode == 2'h1) begin
      strm_ctrl_muxed = strm_data_valid;
    end
    else strm_ctrl_muxed = 1'h0;
  end
  else begin
    data_flush_w = 1'h0;
    if (cfg_ld_dma_ctrl_valid_mode == 2'h1) begin
      strm_ctrl_muxed = strm_data_valid;
    end
    else strm_ctrl_muxed = strm_data_start_pulse;
  end
end
always_comb begin
  if (cfg_data_network_g2f_mux[0] == 1'h1) begin
    if (cfg_ld_dma_ctrl_valid_mode != 2'h2) begin
      ctrl_g2f_w[0] = strm_ctrl_muxed;
    end
    else ctrl_g2f_w[0] = 1'h0;
  end
  else ctrl_g2f_w[0] = 1'h0;
  if (cfg_data_network_g2f_mux[1] == 1'h1) begin
    if (cfg_ld_dma_ctrl_valid_mode != 2'h2) begin
      ctrl_g2f_w[1] = strm_ctrl_muxed;
    end
    else ctrl_g2f_w[1] = 1'h0;
  end
  else ctrl_g2f_w[1] = 1'h0;
end
always_comb begin
  ld_dma_done_pulse_w = strm_run & loop_done;
end
always_comb begin
  strm_rd_en_w = iter_step_valid;
  strm_rd_addr_w = 19'(data_current_addr);
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    last_strm_rd_addr_r <= 19'h0;
  end
  else if (strm_rd_en_w) begin
    last_strm_rd_addr_r <= strm_rd_addr_w;
  end
end
always_comb begin
  if (cfg_tile_connected_next | cfg_tile_connected_prev) begin
    rdrq_packet_dma2bank_w = 20'h0;
    rdrq_packet_dma2ring_w.rd_en = bank_rdrq_rd_en;
    rdrq_packet_dma2ring_w.rd_addr = bank_rdrq_rd_addr;
  end
  else begin
    rdrq_packet_dma2bank_w.rd_en = bank_rdrq_rd_en;
    rdrq_packet_dma2bank_w.rd_addr = bank_rdrq_rd_addr;
    rdrq_packet_dma2ring_w = 20'h0;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    rdrq_packet_dma2bank <= 20'h0;
    rdrq_packet_dma2ring <= 20'h0;
  end
  else begin
    rdrq_packet_dma2bank <= rdrq_packet_dma2bank_w;
    rdrq_packet_dma2ring <= rdrq_packet_dma2ring_w;
  end
end
always_comb begin
  is_cached = strm_rd_addr_w[18:3] == last_strm_rd_addr_r[18:3];
  bank_rdrq_rd_en = strm_rd_en_w & (is_first | (~is_cached));
  bank_rdrq_rd_addr = strm_rd_addr_w;
end
always_comb begin
  if (cfg_tile_connected_next | cfg_tile_connected_prev) begin
    rdrs_packet = rdrs_packet_ring2dma;
  end
  else rdrs_packet = rdrs_packet_bank2dma;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    bank_rdrs_data_cache_r <= 64'h0;
  end
  else if (rdrs_packet.rd_data_valid) begin
    bank_rdrs_data_cache_r <= rdrs_packet.rd_data;
  end
end
always_comb begin
  unique case (strm_data_sel_arr[5'(cfg_data_network_latency) + 5'h3])
    2'h0: strm_data = bank_rdrs_data_cache_r[15:0];
    2'h1: strm_data = bank_rdrs_data_cache_r[31:16];
    2'h2: strm_data = bank_rdrs_data_cache_r[47:32];
    2'h3: strm_data = bank_rdrs_data_cache_r[63:48];
    default: strm_data = bank_rdrs_data_cache_r[15:0];
  endcase
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    ld_dma_done_pulse_latch <= 1'h0;
  end
  else if (ld_dma_done_pulse_pipeline_out) begin
    ld_dma_done_pulse_latch <= 1'h1;
  end
  else if (ld_dma_done_pulse_latch & all_skid_empty) begin
    ld_dma_done_pulse_latch <= 1'h0;
  end
end
always_comb begin
  if (cfg_ld_dma_ctrl_valid_mode != 2'h2) begin
    ld_dma_done_pulse = ld_dma_done_pulse_pipeline_out;
  end
  else ld_dma_done_pulse = ld_dma_done_pulse_anded;
end
always_comb begin
  ld_dma_done_pulse_anded = ld_dma_done_pulse_latch & all_skid_empty;
end
assign ld_dma_done_pulse_pipeline_out = ld_dma_done_pulse_d_arr[5'(cfg_data_network_latency) + 5'h3 + 5'h2];

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    ld_dma_done_interrupt <= 1'h0;
  end
  else if (ld_dma_done_pulse) begin
    ld_dma_done_interrupt <= 1'h1;
  end
  else if (ld_dma_done_pulse_last) begin
    ld_dma_done_interrupt <= 1'h0;
  end
end
assign clk_en_dma2bank = dma2bank_clk_en;
assign pipeline_ctrl_in[0] = ctrl_g2f_w[0];
assign pipeline_ctrl_in[1] = ctrl_g2f_w[1];
assign ctrl_g2f[0] = pipeline_ctrl_out[0];
assign ctrl_g2f[1] = pipeline_ctrl_out[1];
assign loop_iter_ranges[0] = current_dma_header.range_0;
assign loop_iter_ranges[1] = current_dma_header.range_1;
assign loop_iter_ranges[2] = current_dma_header.range_2;
assign loop_iter_ranges[3] = current_dma_header.range_3;
assign loop_iter_ranges[4] = current_dma_header.range_4;
assign loop_iter_ranges[5] = current_dma_header.range_5;
assign loop_iter_ranges[6] = current_dma_header.range_6;
assign loop_iter_ranges[7] = current_dma_header.range_7;
assign cycle_counter_en = cfg_ld_dma_ctrl_valid_mode != 2'h2;
assign cycle_stride_addr_gen_strides[0] = current_dma_header.cycle_stride_0;
assign cycle_stride_addr_gen_strides[1] = current_dma_header.cycle_stride_1;
assign cycle_stride_addr_gen_strides[2] = current_dma_header.cycle_stride_2;
assign cycle_stride_addr_gen_strides[3] = current_dma_header.cycle_stride_3;
assign cycle_stride_addr_gen_strides[4] = current_dma_header.cycle_stride_4;
assign cycle_stride_addr_gen_strides[5] = current_dma_header.cycle_stride_5;
assign cycle_stride_addr_gen_strides[6] = current_dma_header.cycle_stride_6;
assign cycle_stride_addr_gen_strides[7] = current_dma_header.cycle_stride_7;
assign data_stride_addr_gen_start_addr = 20'(current_dma_header.start_addr);
assign data_stride_addr_gen_strides[0] = current_dma_header.stride_0;
assign data_stride_addr_gen_strides[1] = current_dma_header.stride_1;
assign data_stride_addr_gen_strides[2] = current_dma_header.stride_2;
assign data_stride_addr_gen_strides[3] = current_dma_header.stride_3;
assign data_stride_addr_gen_strides[4] = current_dma_header.stride_4;
assign data_stride_addr_gen_strides[5] = current_dma_header.stride_5;
assign data_stride_addr_gen_strides[6] = current_dma_header.stride_6;
assign data_stride_addr_gen_strides[7] = current_dma_header.stride_7;
reg_fifo_d_19_w_16 #(
  .data_width(16'h10))
data_g2f_fifo (
  .almost_empty_diff(5'h2),
  .almost_full_diff(fifo_almost_full_diff),
  .clk(clk),
  .clk_en(1'h1),
  .data_in(data_dma2fifo),
  .flush(ld_dma_start_pulse_r),
  .pop(fifo_pop),
  .push(fifo_push),
  .reset(reset),
  .almost_full(fifo_almost_full),
  .data_out(data_fifo2cgra),
  .empty(fifo_empty),
  .full(fifo_full)
);

reg_fifo_d_2_w_16 #(
  .data_width(16'h10))
data_g2f_skid_0 (
  .almost_empty_diff(1'h0),
  .almost_full_diff(1'h0),
  .clk(clk),
  .clk_en(1'h1),
  .data_in(skid_in[0]),
  .flush(ld_dma_start_pulse_r),
  .pop(skid_pop[0]),
  .push(skid_push[0]),
  .reset(reset),
  .data_out(data_g2f_skid_0_data_out),
  .empty(data_g2f_skid_0_empty),
  .full(data_g2f_skid_0_full)
);

reg_fifo_d_2_w_16 #(
  .data_width(16'h10))
data_g2f_skid_1 (
  .almost_empty_diff(1'h0),
  .almost_full_diff(1'h0),
  .clk(clk),
  .clk_en(1'h1),
  .data_in(skid_in[1]),
  .flush(ld_dma_start_pulse_r),
  .pop(skid_pop[1]),
  .push(skid_push[1]),
  .reset(reset),
  .data_out(data_g2f_skid_1_data_out),
  .empty(data_g2f_skid_1_empty),
  .full(data_g2f_skid_1_full)
);

pipeline_w_1_d_22_array strm_dma_start_pulse_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(ld_dma_start_pulse_r),
  .reset(reset),
  .out_(strm_data_start_pulse_d_arr)
);

pipeline_w_1_d_22_array strm_rd_en_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(strm_rd_en_w),
  .reset(reset),
  .out_(strm_rd_en_d_arr)
);

pipeline_w_2_d_22_array strm_data_sel_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(strm_data_sel_w),
  .reset(reset),
  .out_(strm_data_sel_arr)
);

pipeline_w_1_d_24_array ld_dma_done_pulse_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(ld_dma_done_pulse_w),
  .reset(reset),
  .out_(ld_dma_done_pulse_d_arr)
);

pipeline_w_1_d_5 ld_dma_interrupt_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(ld_dma_done_pulse),
  .reset(reset),
  .out_(ld_dma_done_pulse_last)
);

glb_clk_en_gen_6 #(
  .cnt(32'h6))
dma2bank_clk_en_gen (
  .clk(clk),
  .enable(rdrq_packet_dma2bank_w.rd_en),
  .reset(reset),
  .clk_en(dma2bank_clk_en)
);

pipeline_w_2_d_2 pipeline_ctrl (
  .clk(clk),
  .clk_en(1'h1),
  .in_(pipeline_ctrl_in),
  .reset(reset),
  .out_(pipeline_ctrl_out)
);

pipeline_w_1_d_0 pipeline_flush (
  .clk(clk),
  .clk_en(1'h1),
  .in_(data_flush_w),
  .reset(reset),
  .out_(data_flush)
);

glb_loop_iter_8 loop_iter (
  .clk(clk),
  .clk_en(1'h1),
  .dim(current_dma_header.dim),
  .ranges(loop_iter_ranges),
  .reset(reset),
  .step(iter_step_valid),
  .mux_sel_out(loop_mux_sel),
  .restart(loop_done)
);

glb_sched_gen cycle_stride_sched_gen (
  .clk(clk),
  .clk_en(cycle_counter_en),
  .current_addr(cycle_current_addr),
  .cycle_count(cycle_count),
  .finished(loop_done),
  .reset(reset),
  .restart(ld_dma_start_pulse_r),
  .valid_output(cycle_valid)
);

glb_addr_gen_8 #(
  .addr_width(32'h10),
  .loop_level(32'h8))
cycle_stride_addr_gen (
  .clk(clk),
  .clk_en(cycle_counter_en),
  .mux_sel(loop_mux_sel),
  .reset(reset),
  .restart(ld_dma_start_pulse_r),
  .start_addr(current_dma_header.cycle_start_addr),
  .step(iter_step_valid),
  .strides(cycle_stride_addr_gen_strides),
  .addr_out(cycle_current_addr)
);

glb_addr_gen_8 #(
  .addr_width(32'h14),
  .loop_level(32'h8))
data_stride_addr_gen (
  .clk(clk),
  .clk_en(1'h1),
  .mux_sel(loop_mux_sel),
  .reset(reset),
  .restart(ld_dma_start_pulse_r),
  .start_addr(data_stride_addr_gen_start_addr),
  .step(iter_step_valid),
  .strides(data_stride_addr_gen_strides),
  .addr_out(data_current_addr)
);

endmodule   // glb_load_dma

module glb_loop_iter_7 (
  input logic clk,
  input logic clk_en,
  input logic [3:0] dim,
  input logic [6:0] [31:0] ranges,
  input logic reset,
  input logic step,
  output logic [2:0] mux_sel_out,
  output logic restart
);

logic [6:0] clear;
logic [6:0][31:0] dim_counter;
logic [6:0] inc;
logic is_maxed;
logic [6:0] max_value;
logic [2:0] mux_sel;
logic not_done;
assign mux_sel_out = mux_sel;
assign is_maxed = (dim_counter[mux_sel] == ranges[mux_sel]) & inc[mux_sel];
always_comb begin
  mux_sel = 3'h0;
  not_done = 1'h0;
  for (int unsigned i = 0; i < 7; i += 1) begin
      if (~not_done) begin
        if ((~max_value[3'(i)]) & (4'(i) < dim)) begin
          mux_sel = 3'(i);
          not_done = 1'h1;
        end
      end
    end
end
always_comb begin
  clear[0] = 1'h0;
  if (((mux_sel > 3'h0) | (~not_done)) & step) begin
    clear[0] = 1'h1;
  end
end
always_comb begin
  inc[0] = 1'h0;
  if ((5'h0 == 5'h0) & step & (dim > 4'h0)) begin
    inc[0] = 1'h1;
  end
  else if ((mux_sel == 3'h0) & step & (dim > 4'h0)) begin
    inc[0] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[0] <= 32'h0;
  end
  else if (clear[0]) begin
    dim_counter[0] <= 32'h0;
  end
  else if (inc[0]) begin
    dim_counter[0] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[0] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[0]) begin
      max_value[0] <= 1'h0;
    end
    else if (inc[0]) begin
      max_value[0] <= is_maxed;
    end
  end
end
always_comb begin
  clear[1] = 1'h0;
  if (((mux_sel > 3'h1) | (~not_done)) & step) begin
    clear[1] = 1'h1;
  end
end
always_comb begin
  inc[1] = 1'h0;
  if ((5'h1 == 5'h0) & step & (dim > 4'h1)) begin
    inc[1] = 1'h1;
  end
  else if ((mux_sel == 3'h1) & step & (dim > 4'h1)) begin
    inc[1] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[1] <= 32'h0;
  end
  else if (clear[1]) begin
    dim_counter[1] <= 32'h0;
  end
  else if (inc[1]) begin
    dim_counter[1] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[1] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[1]) begin
      max_value[1] <= 1'h0;
    end
    else if (inc[1]) begin
      max_value[1] <= is_maxed;
    end
  end
end
always_comb begin
  clear[2] = 1'h0;
  if (((mux_sel > 3'h2) | (~not_done)) & step) begin
    clear[2] = 1'h1;
  end
end
always_comb begin
  inc[2] = 1'h0;
  if ((5'h2 == 5'h0) & step & (dim > 4'h2)) begin
    inc[2] = 1'h1;
  end
  else if ((mux_sel == 3'h2) & step & (dim > 4'h2)) begin
    inc[2] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[2] <= 32'h0;
  end
  else if (clear[2]) begin
    dim_counter[2] <= 32'h0;
  end
  else if (inc[2]) begin
    dim_counter[2] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[2] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[2]) begin
      max_value[2] <= 1'h0;
    end
    else if (inc[2]) begin
      max_value[2] <= is_maxed;
    end
  end
end
always_comb begin
  clear[3] = 1'h0;
  if (((mux_sel > 3'h3) | (~not_done)) & step) begin
    clear[3] = 1'h1;
  end
end
always_comb begin
  inc[3] = 1'h0;
  if ((5'h3 == 5'h0) & step & (dim > 4'h3)) begin
    inc[3] = 1'h1;
  end
  else if ((mux_sel == 3'h3) & step & (dim > 4'h3)) begin
    inc[3] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[3] <= 32'h0;
  end
  else if (clear[3]) begin
    dim_counter[3] <= 32'h0;
  end
  else if (inc[3]) begin
    dim_counter[3] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[3] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[3]) begin
      max_value[3] <= 1'h0;
    end
    else if (inc[3]) begin
      max_value[3] <= is_maxed;
    end
  end
end
always_comb begin
  clear[4] = 1'h0;
  if (((mux_sel > 3'h4) | (~not_done)) & step) begin
    clear[4] = 1'h1;
  end
end
always_comb begin
  inc[4] = 1'h0;
  if ((5'h4 == 5'h0) & step & (dim > 4'h4)) begin
    inc[4] = 1'h1;
  end
  else if ((mux_sel == 3'h4) & step & (dim > 4'h4)) begin
    inc[4] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[4] <= 32'h0;
  end
  else if (clear[4]) begin
    dim_counter[4] <= 32'h0;
  end
  else if (inc[4]) begin
    dim_counter[4] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[4] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[4]) begin
      max_value[4] <= 1'h0;
    end
    else if (inc[4]) begin
      max_value[4] <= is_maxed;
    end
  end
end
always_comb begin
  clear[5] = 1'h0;
  if (((mux_sel > 3'h5) | (~not_done)) & step) begin
    clear[5] = 1'h1;
  end
end
always_comb begin
  inc[5] = 1'h0;
  if ((5'h5 == 5'h0) & step & (dim > 4'h5)) begin
    inc[5] = 1'h1;
  end
  else if ((mux_sel == 3'h5) & step & (dim > 4'h5)) begin
    inc[5] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[5] <= 32'h0;
  end
  else if (clear[5]) begin
    dim_counter[5] <= 32'h0;
  end
  else if (inc[5]) begin
    dim_counter[5] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[5] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[5]) begin
      max_value[5] <= 1'h0;
    end
    else if (inc[5]) begin
      max_value[5] <= is_maxed;
    end
  end
end
always_comb begin
  clear[6] = 1'h0;
  if (((mux_sel > 3'h6) | (~not_done)) & step) begin
    clear[6] = 1'h1;
  end
end
always_comb begin
  inc[6] = 1'h0;
  if ((5'h6 == 5'h0) & step & (dim > 4'h6)) begin
    inc[6] = 1'h1;
  end
  else if ((mux_sel == 3'h6) & step & (dim > 4'h6)) begin
    inc[6] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[6] <= 32'h0;
  end
  else if (clear[6]) begin
    dim_counter[6] <= 32'h0;
  end
  else if (inc[6]) begin
    dim_counter[6] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[6] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[6]) begin
      max_value[6] <= 1'h0;
    end
    else if (inc[6]) begin
      max_value[6] <= is_maxed;
    end
  end
end
assign restart = step & (~not_done);
endmodule   // glb_loop_iter_7

module glb_loop_iter_8 (
  input logic clk,
  input logic clk_en,
  input logic [3:0] dim,
  input logic [7:0] [31:0] ranges,
  input logic reset,
  input logic step,
  output logic [2:0] mux_sel_out,
  output logic restart
);

logic [7:0] clear;
logic [7:0][31:0] dim_counter;
logic [7:0] inc;
logic is_maxed;
logic [7:0] max_value;
logic [2:0] mux_sel;
logic not_done;
assign mux_sel_out = mux_sel;
assign is_maxed = (dim_counter[mux_sel] == ranges[mux_sel]) & inc[mux_sel];
always_comb begin
  mux_sel = 3'h0;
  not_done = 1'h0;
  for (int unsigned i = 0; i < 8; i += 1) begin
      if (~not_done) begin
        if ((~max_value[3'(i)]) & (4'(i) < dim)) begin
          mux_sel = 3'(i);
          not_done = 1'h1;
        end
      end
    end
end
always_comb begin
  clear[0] = 1'h0;
  if (((mux_sel > 3'h0) | (~not_done)) & step) begin
    clear[0] = 1'h1;
  end
end
always_comb begin
  inc[0] = 1'h0;
  if ((5'h0 == 5'h0) & step & (dim > 4'h0)) begin
    inc[0] = 1'h1;
  end
  else if ((mux_sel == 3'h0) & step & (dim > 4'h0)) begin
    inc[0] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[0] <= 32'h0;
  end
  else if (clear[0]) begin
    dim_counter[0] <= 32'h0;
  end
  else if (inc[0]) begin
    dim_counter[0] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[0] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[0]) begin
      max_value[0] <= 1'h0;
    end
    else if (inc[0]) begin
      max_value[0] <= is_maxed;
    end
  end
end
always_comb begin
  clear[1] = 1'h0;
  if (((mux_sel > 3'h1) | (~not_done)) & step) begin
    clear[1] = 1'h1;
  end
end
always_comb begin
  inc[1] = 1'h0;
  if ((5'h1 == 5'h0) & step & (dim > 4'h1)) begin
    inc[1] = 1'h1;
  end
  else if ((mux_sel == 3'h1) & step & (dim > 4'h1)) begin
    inc[1] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[1] <= 32'h0;
  end
  else if (clear[1]) begin
    dim_counter[1] <= 32'h0;
  end
  else if (inc[1]) begin
    dim_counter[1] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[1] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[1]) begin
      max_value[1] <= 1'h0;
    end
    else if (inc[1]) begin
      max_value[1] <= is_maxed;
    end
  end
end
always_comb begin
  clear[2] = 1'h0;
  if (((mux_sel > 3'h2) | (~not_done)) & step) begin
    clear[2] = 1'h1;
  end
end
always_comb begin
  inc[2] = 1'h0;
  if ((5'h2 == 5'h0) & step & (dim > 4'h2)) begin
    inc[2] = 1'h1;
  end
  else if ((mux_sel == 3'h2) & step & (dim > 4'h2)) begin
    inc[2] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[2] <= 32'h0;
  end
  else if (clear[2]) begin
    dim_counter[2] <= 32'h0;
  end
  else if (inc[2]) begin
    dim_counter[2] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[2] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[2]) begin
      max_value[2] <= 1'h0;
    end
    else if (inc[2]) begin
      max_value[2] <= is_maxed;
    end
  end
end
always_comb begin
  clear[3] = 1'h0;
  if (((mux_sel > 3'h3) | (~not_done)) & step) begin
    clear[3] = 1'h1;
  end
end
always_comb begin
  inc[3] = 1'h0;
  if ((5'h3 == 5'h0) & step & (dim > 4'h3)) begin
    inc[3] = 1'h1;
  end
  else if ((mux_sel == 3'h3) & step & (dim > 4'h3)) begin
    inc[3] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[3] <= 32'h0;
  end
  else if (clear[3]) begin
    dim_counter[3] <= 32'h0;
  end
  else if (inc[3]) begin
    dim_counter[3] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[3] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[3]) begin
      max_value[3] <= 1'h0;
    end
    else if (inc[3]) begin
      max_value[3] <= is_maxed;
    end
  end
end
always_comb begin
  clear[4] = 1'h0;
  if (((mux_sel > 3'h4) | (~not_done)) & step) begin
    clear[4] = 1'h1;
  end
end
always_comb begin
  inc[4] = 1'h0;
  if ((5'h4 == 5'h0) & step & (dim > 4'h4)) begin
    inc[4] = 1'h1;
  end
  else if ((mux_sel == 3'h4) & step & (dim > 4'h4)) begin
    inc[4] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[4] <= 32'h0;
  end
  else if (clear[4]) begin
    dim_counter[4] <= 32'h0;
  end
  else if (inc[4]) begin
    dim_counter[4] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[4] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[4]) begin
      max_value[4] <= 1'h0;
    end
    else if (inc[4]) begin
      max_value[4] <= is_maxed;
    end
  end
end
always_comb begin
  clear[5] = 1'h0;
  if (((mux_sel > 3'h5) | (~not_done)) & step) begin
    clear[5] = 1'h1;
  end
end
always_comb begin
  inc[5] = 1'h0;
  if ((5'h5 == 5'h0) & step & (dim > 4'h5)) begin
    inc[5] = 1'h1;
  end
  else if ((mux_sel == 3'h5) & step & (dim > 4'h5)) begin
    inc[5] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[5] <= 32'h0;
  end
  else if (clear[5]) begin
    dim_counter[5] <= 32'h0;
  end
  else if (inc[5]) begin
    dim_counter[5] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[5] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[5]) begin
      max_value[5] <= 1'h0;
    end
    else if (inc[5]) begin
      max_value[5] <= is_maxed;
    end
  end
end
always_comb begin
  clear[6] = 1'h0;
  if (((mux_sel > 3'h6) | (~not_done)) & step) begin
    clear[6] = 1'h1;
  end
end
always_comb begin
  inc[6] = 1'h0;
  if ((5'h6 == 5'h0) & step & (dim > 4'h6)) begin
    inc[6] = 1'h1;
  end
  else if ((mux_sel == 3'h6) & step & (dim > 4'h6)) begin
    inc[6] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[6] <= 32'h0;
  end
  else if (clear[6]) begin
    dim_counter[6] <= 32'h0;
  end
  else if (inc[6]) begin
    dim_counter[6] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[6] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[6]) begin
      max_value[6] <= 1'h0;
    end
    else if (inc[6]) begin
      max_value[6] <= is_maxed;
    end
  end
end
always_comb begin
  clear[7] = 1'h0;
  if (((mux_sel > 3'h7) | (~not_done)) & step) begin
    clear[7] = 1'h1;
  end
end
always_comb begin
  inc[7] = 1'h0;
  if ((5'h7 == 5'h0) & step & (dim > 4'h7)) begin
    inc[7] = 1'h1;
  end
  else if ((mux_sel == 3'h7) & step & (dim > 4'h7)) begin
    inc[7] = 1'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    dim_counter[7] <= 32'h0;
  end
  else if (clear[7]) begin
    dim_counter[7] <= 32'h0;
  end
  else if (inc[7]) begin
    dim_counter[7] <= dim_counter[mux_sel] + 32'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    max_value[7] <= 1'h0;
  end
  else if (clk_en) begin
    if (clear[7]) begin
      max_value[7] <= 1'h0;
    end
    else if (inc[7]) begin
      max_value[7] <= is_maxed;
    end
  end
end
assign restart = step & (~not_done);
endmodule   // glb_loop_iter_8

module glb_pcfg_broadcast (
  input pcfg_broadcast_mux_t cfg_pcfg_broadcast_mux,
  input cgra_cfg_t cgra_cfg_dma2mux,
  input logic [31:0] cgra_cfg_jtag_addr_bypass_wsti,
  input logic cgra_cfg_jtag_rd_en_bypass_wsti,
  input cgra_cfg_t cgra_cfg_jtag_wsti,
  input cgra_cfg_t cgra_cfg_pcfg_esti,
  input cgra_cfg_t cgra_cfg_pcfg_wsti,
  input logic clk,
  input logic reset,
  output cgra_cfg_t [1:0] cgra_cfg_g2f,
  output logic [31:0] cgra_cfg_jtag_addr_bypass_esto,
  output cgra_cfg_t cgra_cfg_jtag_esto,
  output logic cgra_cfg_jtag_rd_en_bypass_esto,
  output cgra_cfg_t cgra_cfg_pcfg_esto,
  output cgra_cfg_t cgra_cfg_pcfg_wsto
);

cgra_cfg_t [1:0] cgra_cfg_g2f_w;
cgra_cfg_t pcfg_east_muxed;
cgra_cfg_t pcfg_south_muxed;
cgra_cfg_t pcfg_west_muxed;
always_comb begin
  cgra_cfg_jtag_rd_en_bypass_esto = cgra_cfg_jtag_rd_en_bypass_wsti;
  cgra_cfg_jtag_addr_bypass_esto = cgra_cfg_jtag_addr_bypass_wsti;
end
always_comb begin
  if (cfg_pcfg_broadcast_mux.south == 2'h0) begin
    pcfg_south_muxed = 66'h0;
  end
  else if (cfg_pcfg_broadcast_mux.south == 2'h1) begin
    pcfg_south_muxed = cgra_cfg_dma2mux;
  end
  else if (cfg_pcfg_broadcast_mux.south == 2'h2) begin
    pcfg_south_muxed = cgra_cfg_pcfg_wsti;
  end
  else if (cfg_pcfg_broadcast_mux.south == 2'h3) begin
    pcfg_south_muxed = cgra_cfg_pcfg_esti;
  end
  else pcfg_south_muxed = 66'h0;
end
always_comb begin
  if (cfg_pcfg_broadcast_mux.west == 2'h0) begin
    pcfg_west_muxed = 66'h0;
  end
  else if (cfg_pcfg_broadcast_mux.west == 2'h1) begin
    pcfg_west_muxed = cgra_cfg_dma2mux;
  end
  else if (cfg_pcfg_broadcast_mux.west == 2'h2) begin
    pcfg_west_muxed = cgra_cfg_pcfg_esti;
  end
  else pcfg_west_muxed = 66'h0;
end
always_comb begin
  if (cfg_pcfg_broadcast_mux.east == 2'h0) begin
    pcfg_east_muxed = 66'h0;
  end
  else if (cfg_pcfg_broadcast_mux.east == 2'h1) begin
    pcfg_east_muxed = cgra_cfg_dma2mux;
  end
  else if (cfg_pcfg_broadcast_mux.east == 2'h2) begin
    pcfg_east_muxed = cgra_cfg_pcfg_wsti;
  end
  else pcfg_east_muxed = 66'h0;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    cgra_cfg_jtag_esto <= 66'h0;
  end
  else cgra_cfg_jtag_esto <= cgra_cfg_jtag_wsti;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    cgra_cfg_pcfg_esto <= 66'h0;
    cgra_cfg_pcfg_wsto <= 66'h0;
  end
  else begin
    cgra_cfg_pcfg_esto <= pcfg_east_muxed;
    cgra_cfg_pcfg_wsto <= pcfg_west_muxed;
  end
end
always_comb begin
  if (cgra_cfg_jtag_rd_en_bypass_esto) begin
    cgra_cfg_g2f_w[0].wr_en = 1'h0;
    cgra_cfg_g2f_w[0].rd_en = 1'h1;
    cgra_cfg_g2f_w[0].addr = cgra_cfg_jtag_addr_bypass_esto;
    cgra_cfg_g2f_w[0].data = 32'h0;
  end
  else cgra_cfg_g2f_w[0] = cgra_cfg_jtag_wsti | pcfg_south_muxed;
end
always_comb begin
  if (cgra_cfg_jtag_rd_en_bypass_esto) begin
    cgra_cfg_g2f_w[1].wr_en = 1'h0;
    cgra_cfg_g2f_w[1].rd_en = 1'h1;
    cgra_cfg_g2f_w[1].addr = cgra_cfg_jtag_addr_bypass_esto;
    cgra_cfg_g2f_w[1].data = 32'h0;
  end
  else cgra_cfg_g2f_w[1] = cgra_cfg_jtag_wsti | pcfg_south_muxed;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    for (int unsigned i = 0; i < 2; i += 1) begin
        cgra_cfg_g2f[1'(i)] <= 66'h0;
      end
  end
  else begin
    for (int unsigned i = 0; i < 2; i += 1) begin
        cgra_cfg_g2f[1'(i)] <= cgra_cfg_g2f_w[1'(i)];
      end
  end
end
endmodule   // glb_pcfg_broadcast

module glb_pcfg_dma (
  input logic cfg_pcfg_dma_ctrl_mode,
  input logic cfg_pcfg_dma_ctrl_relocation_is_msb,
  input logic [15:0] cfg_pcfg_dma_ctrl_relocation_value,
  input pcfg_dma_header_t cfg_pcfg_dma_header,
  input logic [5:0] cfg_pcfg_network_latency,
  input logic cfg_pcfg_tile_connected_next,
  input logic cfg_pcfg_tile_connected_prev,
  input logic clk,
  input logic glb_tile_id,
  input logic pcfg_dma_start_pulse,
  input rdrs_packet_t rdrs_packet_bank2dma,
  input rdrs_packet_t rdrs_packet_ring2dma,
  input logic reset,
  output cgra_cfg_t cgra_cfg_pcfg,
  output logic clk_en_dma2bank,
  output logic pcfg_dma_done_interrupt,
  output rdrq_packet_t rdrq_packet_dma2bank,
  output rdrq_packet_t rdrq_packet_dma2ring
);

logic [18:0] addr_next;
logic [18:0] addr_r;
logic dma2bank_clk_en;
logic done_pulse_d_arr [11:0];
logic done_pulse_r;
logic is_running_r;
logic [15:0] num_cfg_cnt_next;
logic [15:0] num_cfg_cnt_r;
logic pcfg_done_pulse;
logic pcfg_done_pulse_last;
rdrq_packet_t rdrq_packet_dma2bank_w;
rdrq_packet_t rdrq_packet_dma2ring_w;
logic [18:0] rdrq_packet_rd_addr_next;
logic rdrq_packet_rd_en_next;
rdrs_packet_t rdrs_packet;
logic [63:0] rdrs_packet_rd_data_r;
logic rdrs_packet_rd_data_valid_r;
logic start_pulse_r;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    start_pulse_r <= 1'h0;
  end
  else if ((cfg_pcfg_dma_ctrl_mode == 1'h1) & (~is_running_r) & pcfg_dma_start_pulse) begin
    start_pulse_r <= 1'h1;
  end
  else start_pulse_r <= 1'h0;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    done_pulse_r <= 1'h0;
  end
  else if (is_running_r & (num_cfg_cnt_r == 16'h0)) begin
    done_pulse_r <= 1'h1;
  end
  else done_pulse_r <= 1'h0;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    is_running_r <= 1'h0;
  end
  else if (start_pulse_r) begin
    is_running_r <= 1'h1;
  end
  else if ((is_running_r == 1'h1) & (num_cfg_cnt_r == 16'h0)) begin
    is_running_r <= 1'h0;
  end
end
always_comb begin
  if (start_pulse_r) begin
    num_cfg_cnt_next = cfg_pcfg_dma_header.num_cfg;
    addr_next = cfg_pcfg_dma_header.start_addr;
  end
  else if ((is_running_r == 1'h1) & (num_cfg_cnt_r > 16'h0)) begin
    num_cfg_cnt_next = num_cfg_cnt_r - 16'h1;
    addr_next = addr_r + 19'h8;
  end
  else begin
    num_cfg_cnt_next = 16'h0;
    addr_next = 19'h0;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    num_cfg_cnt_r <= 16'h0;
    addr_r <= 19'h0;
  end
  else begin
    num_cfg_cnt_r <= num_cfg_cnt_next;
    addr_r <= addr_next;
  end
end
always_comb begin
  if (is_running_r & (num_cfg_cnt_r > 16'h0)) begin
    rdrq_packet_rd_en_next = 1'h1;
    rdrq_packet_rd_addr_next = addr_r;
  end
  else begin
    rdrq_packet_rd_en_next = 1'h0;
    rdrq_packet_rd_addr_next = 19'h0;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    rdrq_packet_dma2ring <= 20'h0;
    rdrq_packet_dma2bank <= 20'h0;
  end
  else begin
    rdrq_packet_dma2ring <= rdrq_packet_dma2ring_w;
    rdrq_packet_dma2bank <= rdrq_packet_dma2bank_w;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    rdrs_packet_rd_data_r <= 64'h0;
    rdrs_packet_rd_data_valid_r <= 1'h0;
  end
  else if (rdrs_packet.rd_data_valid) begin
    rdrs_packet_rd_data_r <= rdrs_packet.rd_data;
    rdrs_packet_rd_data_valid_r <= 1'h1;
  end
  else begin
    rdrs_packet_rd_data_r <= 64'h0;
    rdrs_packet_rd_data_valid_r <= 1'h0;
  end
end
always_comb begin
  if (cfg_pcfg_tile_connected_next | cfg_pcfg_tile_connected_prev) begin
    rdrq_packet_dma2ring_w.rd_en = rdrq_packet_rd_en_next;
    rdrq_packet_dma2ring_w.rd_addr = rdrq_packet_rd_addr_next;
    rdrq_packet_dma2bank_w.rd_en = 1'h0;
    rdrq_packet_dma2bank_w.rd_addr = 19'h0;
  end
  else begin
    rdrq_packet_dma2ring_w.rd_en = 1'h0;
    rdrq_packet_dma2ring_w.rd_addr = 19'h0;
    rdrq_packet_dma2bank_w.rd_en = rdrq_packet_rd_en_next;
    rdrq_packet_dma2bank_w.rd_addr = rdrq_packet_rd_addr_next;
  end
end
always_comb begin
  if (cfg_pcfg_tile_connected_next | cfg_pcfg_tile_connected_prev) begin
    rdrs_packet = rdrs_packet_ring2dma;
  end
  else rdrs_packet = rdrs_packet_bank2dma;
end
always_comb begin
  cgra_cfg_pcfg.rd_en = 1'h0;
  cgra_cfg_pcfg.wr_en = rdrs_packet_rd_data_valid_r;
  cgra_cfg_pcfg.data = rdrs_packet_rd_data_r[31:0];
  if (cfg_pcfg_dma_ctrl_relocation_is_msb) begin
    cgra_cfg_pcfg.addr = rdrs_packet_rd_data_r[63:32] + 32'(cfg_pcfg_dma_ctrl_relocation_value << 16'h10);
  end
  else cgra_cfg_pcfg.addr = rdrs_packet_rd_data_r[63:32] + 32'(cfg_pcfg_dma_ctrl_relocation_value);
end
assign pcfg_done_pulse = done_pulse_d_arr[4'(cfg_pcfg_network_latency) + 4'h3 + 4'h2];

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    pcfg_dma_done_interrupt <= 1'h0;
  end
  else if (pcfg_done_pulse) begin
    pcfg_dma_done_interrupt <= 1'h1;
  end
  else if (pcfg_done_pulse_last) begin
    pcfg_dma_done_interrupt <= 1'h0;
  end
end
assign clk_en_dma2bank = dma2bank_clk_en;
pipeline_w_1_d_12_array done_pulse_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(done_pulse_r),
  .reset(reset),
  .out_(done_pulse_d_arr)
);

pipeline_w_1_d_5 pcfg_dma_interrupt_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(pcfg_done_pulse),
  .reset(reset),
  .out_(pcfg_done_pulse_last)
);

glb_clk_en_gen_6 #(
  .cnt(32'h6))
dma2bank_clk_en_gen (
  .clk(clk),
  .enable(rdrq_packet_dma2bank_w.rd_en),
  .reset(reset),
  .clk_en(dma2bank_clk_en)
);

endmodule   // glb_pcfg_dma

module glb_ring_switch_RD (
  input logic cfg_ld_dma_on,
  input logic cfg_tile_connected_next,
  input logic cfg_tile_connected_prev,
  input logic clk,
  input logic glb_tile_id,
  input rdrq_packet_t rdrq_packet_dma2ring,
  input rdrq_packet_t rdrq_packet_e2w_esti,
  input rdrq_packet_t rdrq_packet_w2e_wsti,
  input rdrs_packet_t rdrs_packet_bank2ring,
  input rdrs_packet_t rdrs_packet_e2w_esti,
  input rdrs_packet_t rdrs_packet_w2e_wsti,
  input logic reset,
  output logic clk_en_ring2bank,
  output rdrq_packet_t rdrq_packet_e2w_wsto,
  output rdrq_packet_t rdrq_packet_ring2bank,
  output rdrq_packet_t rdrq_packet_w2e_esto,
  output rdrs_packet_t rdrs_packet_e2w_wsto,
  output rdrs_packet_t rdrs_packet_ring2dma,
  output rdrs_packet_t rdrs_packet_w2e_esto
);

rdrq_packet_t rdrq_packet_e2w_esti_muxed;
rdrq_packet_t rdrq_packet_e2w_wsto_w;
rdrq_packet_t rdrq_packet_ring2bank_w;
rdrq_packet_t rdrq_packet_w2e_esto_w;
rdrq_packet_t rdrq_packet_w2e_wsti_muxed;
rdrs_packet_t rdrs_packet_e2w_esti_muxed;
rdrs_packet_t rdrs_packet_e2w_wsto_w;
rdrs_packet_t rdrs_packet_ring2dma_w;
rdrs_packet_t rdrs_packet_w2e_esto_w;
rdrs_packet_t rdrs_packet_w2e_wsti_muxed;
logic ring2bank_rd_clk_en;
always_comb begin
  if (cfg_tile_connected_prev) begin
    rdrq_packet_w2e_wsti_muxed = rdrq_packet_w2e_wsti;
    rdrs_packet_w2e_wsti_muxed = rdrs_packet_w2e_wsti;
  end
  else begin
    rdrq_packet_w2e_wsti_muxed = rdrq_packet_e2w_wsto;
    rdrs_packet_w2e_wsti_muxed = rdrs_packet_e2w_wsto;
  end
end
always_comb begin
  if (cfg_tile_connected_next) begin
    rdrq_packet_e2w_esti_muxed = rdrq_packet_e2w_esti;
    rdrs_packet_e2w_esti_muxed = rdrs_packet_e2w_esti;
  end
  else begin
    rdrq_packet_e2w_esti_muxed = rdrq_packet_w2e_esto;
    rdrs_packet_e2w_esti_muxed = rdrs_packet_w2e_esto;
  end
end
always_comb begin
  if (rdrq_packet_dma2ring.rd_en == 1'h1) begin
    if (rdrq_packet_dma2ring.rd_addr[18] == glb_tile_id) begin
      rdrq_packet_ring2bank_w = rdrq_packet_dma2ring;
      rdrq_packet_w2e_esto_w = 20'h0;
    end
    else begin
      rdrq_packet_ring2bank_w = 20'h0;
      rdrq_packet_w2e_esto_w = rdrq_packet_dma2ring;
    end
  end
  else if (rdrq_packet_w2e_wsti_muxed.rd_en == 1'h1) begin
    if (rdrq_packet_w2e_wsti_muxed.rd_addr[18] == glb_tile_id) begin
      rdrq_packet_ring2bank_w = rdrq_packet_w2e_wsti_muxed;
      rdrq_packet_w2e_esto_w = 20'h0;
    end
    else begin
      rdrq_packet_ring2bank_w = 20'h0;
      rdrq_packet_w2e_esto_w = rdrq_packet_w2e_wsti_muxed;
    end
  end
  else begin
    rdrq_packet_ring2bank_w = 20'h0;
    rdrq_packet_w2e_esto_w = 20'h0;
  end
  rdrq_packet_e2w_wsto_w = rdrq_packet_e2w_esti_muxed;
end
always_comb begin
  if (rdrs_packet_bank2ring.rd_data_valid == 1'h1) begin
    rdrs_packet_w2e_esto_w = rdrs_packet_bank2ring;
  end
  else if (rdrs_packet_w2e_wsti_muxed.rd_data_valid & cfg_ld_dma_on) begin
    rdrs_packet_w2e_esto_w = 65'h0;
  end
  else rdrs_packet_w2e_esto_w = rdrs_packet_w2e_wsti_muxed;
  if (rdrs_packet_w2e_wsti_muxed.rd_data_valid & cfg_ld_dma_on) begin
    rdrs_packet_ring2dma_w = rdrs_packet_w2e_wsti_muxed;
  end
  else rdrs_packet_ring2dma_w = 65'h0;
  rdrs_packet_e2w_wsto_w = rdrs_packet_e2w_esti_muxed;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    rdrq_packet_w2e_esto <= 20'h0;
    rdrq_packet_e2w_wsto <= 20'h0;
    rdrq_packet_ring2bank <= 20'h0;
    rdrs_packet_w2e_esto <= 65'h0;
    rdrs_packet_e2w_wsto <= 65'h0;
  end
  else begin
    rdrq_packet_w2e_esto <= rdrq_packet_w2e_esto_w;
    rdrq_packet_e2w_wsto <= rdrq_packet_e2w_wsto_w;
    rdrq_packet_ring2bank <= rdrq_packet_ring2bank_w;
    rdrs_packet_w2e_esto <= rdrs_packet_w2e_esto_w;
    rdrs_packet_e2w_wsto <= rdrs_packet_e2w_wsto_w;
  end
end
always_comb begin
  rdrs_packet_ring2dma = rdrs_packet_ring2dma_w;
end
assign clk_en_ring2bank = ring2bank_rd_clk_en;
glb_clk_en_gen_6 #(
  .cnt(32'h6))
ring2bank_rd_clk_en_gen (
  .clk(clk),
  .enable(rdrq_packet_ring2bank_w.rd_en),
  .reset(reset),
  .clk_en(ring2bank_rd_clk_en)
);

endmodule   // glb_ring_switch_RD

module glb_ring_switch_WR_RD (
  input logic cfg_ld_dma_on,
  input logic cfg_tile_connected_next,
  input logic cfg_tile_connected_prev,
  input logic clk,
  input logic glb_tile_id,
  input rdrq_packet_t rdrq_packet_dma2ring,
  input rdrq_packet_t rdrq_packet_e2w_esti,
  input rdrq_packet_t rdrq_packet_w2e_wsti,
  input rdrs_packet_t rdrs_packet_bank2ring,
  input rdrs_packet_t rdrs_packet_e2w_esti,
  input rdrs_packet_t rdrs_packet_w2e_wsti,
  input logic reset,
  input wr_packet_t wr_packet_dma2ring,
  input wr_packet_t wr_packet_e2w_esti,
  input wr_packet_t wr_packet_w2e_wsti,
  output logic clk_en_ring2bank,
  output rdrq_packet_t rdrq_packet_e2w_wsto,
  output rdrq_packet_t rdrq_packet_ring2bank,
  output rdrq_packet_t rdrq_packet_w2e_esto,
  output rdrs_packet_t rdrs_packet_e2w_wsto,
  output rdrs_packet_t rdrs_packet_ring2dma,
  output rdrs_packet_t rdrs_packet_w2e_esto,
  output wr_packet_t wr_packet_e2w_wsto,
  output wr_packet_t wr_packet_ring2bank,
  output wr_packet_t wr_packet_w2e_esto
);

rdrq_packet_t rdrq_packet_e2w_esti_muxed;
rdrq_packet_t rdrq_packet_e2w_wsto_w;
rdrq_packet_t rdrq_packet_ring2bank_w;
rdrq_packet_t rdrq_packet_w2e_esto_w;
rdrq_packet_t rdrq_packet_w2e_wsti_muxed;
rdrs_packet_t rdrs_packet_e2w_esti_muxed;
rdrs_packet_t rdrs_packet_e2w_wsto_w;
rdrs_packet_t rdrs_packet_ring2dma_w;
rdrs_packet_t rdrs_packet_w2e_esto_w;
rdrs_packet_t rdrs_packet_w2e_wsti_muxed;
logic ring2bank_rd_clk_en;
logic ring2bank_wr_clk_en;
wr_packet_t wr_packet_e2w_esti_muxed;
wr_packet_t wr_packet_e2w_wsto_w;
wr_packet_t wr_packet_ring2bank_w;
wr_packet_t wr_packet_w2e_esto_w;
wr_packet_t wr_packet_w2e_wsti_muxed;
always_comb begin
  if (cfg_tile_connected_prev) begin
    wr_packet_w2e_wsti_muxed = wr_packet_w2e_wsti;
    rdrq_packet_w2e_wsti_muxed = rdrq_packet_w2e_wsti;
    rdrs_packet_w2e_wsti_muxed = rdrs_packet_w2e_wsti;
  end
  else begin
    wr_packet_w2e_wsti_muxed = wr_packet_e2w_wsto;
    rdrq_packet_w2e_wsti_muxed = rdrq_packet_e2w_wsto;
    rdrs_packet_w2e_wsti_muxed = rdrs_packet_e2w_wsto;
  end
end
always_comb begin
  if (cfg_tile_connected_next) begin
    wr_packet_e2w_esti_muxed = wr_packet_e2w_esti;
    rdrq_packet_e2w_esti_muxed = rdrq_packet_e2w_esti;
    rdrs_packet_e2w_esti_muxed = rdrs_packet_e2w_esti;
  end
  else begin
    wr_packet_e2w_esti_muxed = wr_packet_w2e_esto;
    rdrq_packet_e2w_esti_muxed = rdrq_packet_w2e_esto;
    rdrs_packet_e2w_esti_muxed = rdrs_packet_w2e_esto;
  end
end
always_comb begin
  if (wr_packet_dma2ring.wr_en == 1'h1) begin
    if (wr_packet_dma2ring.wr_addr[18] == glb_tile_id) begin
      wr_packet_ring2bank_w = wr_packet_dma2ring;
      wr_packet_w2e_esto_w = 92'h0;
    end
    else begin
      wr_packet_ring2bank_w = 92'h0;
      wr_packet_w2e_esto_w = wr_packet_dma2ring;
    end
  end
  else if (wr_packet_w2e_wsti_muxed.wr_en == 1'h1) begin
    if (wr_packet_w2e_wsti_muxed.wr_addr[18] == glb_tile_id) begin
      wr_packet_ring2bank_w = wr_packet_w2e_wsti_muxed;
      wr_packet_w2e_esto_w = 92'h0;
    end
    else begin
      wr_packet_ring2bank_w = 92'h0;
      wr_packet_w2e_esto_w = wr_packet_w2e_wsti_muxed;
    end
  end
  else begin
    wr_packet_ring2bank_w = 92'h0;
    wr_packet_w2e_esto_w = 92'h0;
  end
  wr_packet_e2w_wsto_w = wr_packet_e2w_esti_muxed;
end
always_comb begin
  if (rdrq_packet_dma2ring.rd_en == 1'h1) begin
    if (rdrq_packet_dma2ring.rd_addr[18] == glb_tile_id) begin
      rdrq_packet_ring2bank_w = rdrq_packet_dma2ring;
      rdrq_packet_w2e_esto_w = 20'h0;
    end
    else begin
      rdrq_packet_ring2bank_w = 20'h0;
      rdrq_packet_w2e_esto_w = rdrq_packet_dma2ring;
    end
  end
  else if (rdrq_packet_w2e_wsti_muxed.rd_en == 1'h1) begin
    if (rdrq_packet_w2e_wsti_muxed.rd_addr[18] == glb_tile_id) begin
      rdrq_packet_ring2bank_w = rdrq_packet_w2e_wsti_muxed;
      rdrq_packet_w2e_esto_w = 20'h0;
    end
    else begin
      rdrq_packet_ring2bank_w = 20'h0;
      rdrq_packet_w2e_esto_w = rdrq_packet_w2e_wsti_muxed;
    end
  end
  else begin
    rdrq_packet_ring2bank_w = 20'h0;
    rdrq_packet_w2e_esto_w = 20'h0;
  end
  rdrq_packet_e2w_wsto_w = rdrq_packet_e2w_esti_muxed;
end
always_comb begin
  if (rdrs_packet_bank2ring.rd_data_valid == 1'h1) begin
    rdrs_packet_w2e_esto_w = rdrs_packet_bank2ring;
  end
  else if (rdrs_packet_w2e_wsti_muxed.rd_data_valid & cfg_ld_dma_on) begin
    rdrs_packet_w2e_esto_w = 65'h0;
  end
  else rdrs_packet_w2e_esto_w = rdrs_packet_w2e_wsti_muxed;
  if (rdrs_packet_w2e_wsti_muxed.rd_data_valid & cfg_ld_dma_on) begin
    rdrs_packet_ring2dma_w = rdrs_packet_w2e_wsti_muxed;
  end
  else rdrs_packet_ring2dma_w = 65'h0;
  rdrs_packet_e2w_wsto_w = rdrs_packet_e2w_esti_muxed;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    wr_packet_w2e_esto <= 92'h0;
    wr_packet_e2w_wsto <= 92'h0;
    wr_packet_ring2bank <= 92'h0;
    rdrq_packet_w2e_esto <= 20'h0;
    rdrq_packet_e2w_wsto <= 20'h0;
    rdrq_packet_ring2bank <= 20'h0;
    rdrs_packet_w2e_esto <= 65'h0;
    rdrs_packet_e2w_wsto <= 65'h0;
  end
  else begin
    wr_packet_w2e_esto <= wr_packet_w2e_esto_w;
    wr_packet_e2w_wsto <= wr_packet_e2w_wsto_w;
    wr_packet_ring2bank <= wr_packet_ring2bank_w;
    rdrq_packet_w2e_esto <= rdrq_packet_w2e_esto_w;
    rdrq_packet_e2w_wsto <= rdrq_packet_e2w_wsto_w;
    rdrq_packet_ring2bank <= rdrq_packet_ring2bank_w;
    rdrs_packet_w2e_esto <= rdrs_packet_w2e_esto_w;
    rdrs_packet_e2w_wsto <= rdrs_packet_e2w_wsto_w;
  end
end
always_comb begin
  rdrs_packet_ring2dma = rdrs_packet_ring2dma_w;
end
assign clk_en_ring2bank = ring2bank_wr_clk_en | ring2bank_rd_clk_en;
glb_clk_en_gen_4 #(
  .cnt(32'h4))
ring2bank_wr_clk_en_gen (
  .clk(clk),
  .enable(wr_packet_ring2bank_w.wr_en),
  .reset(reset),
  .clk_en(ring2bank_wr_clk_en)
);

glb_clk_en_gen_6 #(
  .cnt(32'h6))
ring2bank_rd_clk_en_gen (
  .clk(clk),
  .enable(rdrq_packet_ring2bank_w.rd_en),
  .reset(reset),
  .clk_en(ring2bank_rd_clk_en)
);

endmodule   // glb_ring_switch_WR_RD

module glb_sched_gen (
  input logic clk,
  input logic clk_en,
  input logic [15:0] current_addr,
  input logic [15:0] cycle_count,
  input logic finished,
  input logic reset,
  input logic restart,
  output logic valid_output
);

logic valid_gate;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    valid_gate <= 1'h1;
  end
  else if (clk_en) begin
    if (restart) begin
      valid_gate <= 1'h0;
    end
    else if (finished) begin
      valid_gate <= 1'h1;
    end
  end
end
always_comb begin
  valid_output = (cycle_count == current_addr) & (~valid_gate);
end
endmodule   // glb_sched_gen

module glb_store_dma (
  input logic [1:0] cfg_data_network_f2g_mux,
  input logic [5:0] cfg_data_network_latency,
  input logic [1:0] cfg_st_dma_ctrl_mode,
  input logic [1:0] cfg_st_dma_ctrl_valid_mode,
  input store_dma_header_t cfg_st_dma_header,
  input logic [31:0] cfg_st_dma_num_blocks,
  input logic cfg_st_dma_num_repeat,
  input logic cfg_tile_connected_next,
  input logic cfg_tile_connected_prev,
  input logic clk,
  input logic [1:0] ctrl_f2g,
  input logic [1:0] [15:0] data_f2g,
  input logic [1:0] data_f2g_vld,
  input logic reset,
  input logic st_dma_start_pulse,
  output logic clk_en_dma2bank,
  output logic [1:0] data_f2g_rdy,
  output logic st_dma_done_interrupt,
  output wr_packet_t wr_packet_dma2bank,
  output wr_packet_t wr_packet_dma2ring
);

logic bank_addr_match;
logic [18:0] bank_wr_addr;
logic [63:0] bank_wr_data_cache_r;
logic [63:0] bank_wr_data_cache_w;
logic bank_wr_en;
logic [7:0] bank_wr_strb_cache_r;
logic [7:0] bank_wr_strb_cache_w;
logic block_done;
logic [1:0] ctrl_f2g_r;
store_dma_header_t current_dma_header;
logic [15:0] cycle_count;
logic cycle_counter_en;
logic [15:0] cycle_current_addr;
logic [6:0][15:0] cycle_stride_addr_gen_strides;
logic cycle_valid;
logic [15:0] data_cgra2fifo;
logic [19:0] data_current_addr;
logic [1:0][15:0] data_f2g_r;
logic [1:0] data_f2g_vld_r;
logic [15:0] data_fifo2dma;
logic data_ready_g2f_w;
logic [19:0] data_stride_addr_gen_start_addr;
logic [6:0][19:0] data_stride_addr_gen_strides;
logic dma2bank_clk_en;
logic done_pulse_d_arr [19:0];
logic done_pulse_w;
logic fifo2cgra_ready;
logic fifo_almost_full;
logic fifo_empty;
logic fifo_full;
logic fifo_pop;
logic fifo_pop_ready;
logic fifo_push;
logic is_first;
logic is_last;
logic is_last_block;
logic iter_step_valid;
logic [18:0] last_strm_wr_addr_r;
logic loop_done;
logic loop_done_muxed;
logic [6:0][31:0] loop_iter_ranges;
logic [2:0] loop_mux_sel;
logic repeat_cnt;
logic rv_is_metadata;
logic rv_mode_on;
logic [31:0] rv_num_blocks_cnt;
logic [15:0] rv_num_data_cnt;
logic st_dma_done_pulse;
logic st_dma_done_pulse_last;
logic st_dma_start_pulse_next;
logic st_dma_start_pulse_r;
logic [15:0] strm_data;
logic [1:0] strm_data_sel;
logic strm_data_valid;
logic strm_run;
logic [18:0] strm_wr_addr_w;
logic [15:0] strm_wr_data_w;
logic strm_wr_en_w;
wr_packet_t wr_packet_dma2bank_w;
wr_packet_t wr_packet_dma2ring_w;
assign current_dma_header = cfg_st_dma_header;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    repeat_cnt <= 1'h0;
  end
  else if (cfg_st_dma_ctrl_mode == 2'h2) begin
    if (st_dma_done_pulse) begin
      if ((repeat_cnt + 1'h1) < cfg_st_dma_num_repeat) begin
        repeat_cnt <= repeat_cnt + 1'h1;
      end
    end
  end
  else if (cfg_st_dma_ctrl_mode == 2'h3) begin
    if (st_dma_done_pulse) begin
      if (((repeat_cnt + 1'h1) < cfg_st_dma_num_repeat) & ((repeat_cnt + 1'h1) < 1'h1)) begin
        repeat_cnt <= repeat_cnt + 1'h1;
      end
    end
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    is_first <= 1'h0;
  end
  else if (st_dma_start_pulse_r) begin
    is_first <= 1'h1;
  end
  else if (strm_wr_en_w) begin
    is_first <= 1'h0;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    is_last <= 1'h0;
  end
  else if (loop_done_muxed) begin
    is_last <= 1'h1;
  end
  else if (bank_wr_en) begin
    is_last <= 1'h0;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    strm_run <= 1'h0;
  end
  else if (st_dma_start_pulse_r) begin
    strm_run <= 1'h1;
  end
  else if (loop_done_muxed) begin
    strm_run <= 1'h0;
  end
end
always_comb begin
  if (cfg_st_dma_ctrl_mode == 2'h0) begin
    st_dma_start_pulse_next = 1'h0;
  end
  else if (cfg_st_dma_ctrl_mode == 2'h1) begin
    st_dma_start_pulse_next = (~strm_run) & st_dma_start_pulse;
  end
  else if ((cfg_st_dma_ctrl_mode == 2'h2) | (cfg_st_dma_ctrl_mode == 2'h3)) begin
    st_dma_start_pulse_next = ((~strm_run) & st_dma_start_pulse) | (st_dma_done_pulse & ((repeat_cnt + 1'h1) <
        cfg_st_dma_num_repeat));
  end
  else st_dma_start_pulse_next = 1'h0;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    st_dma_start_pulse_r <= 1'h0;
  end
  else if (st_dma_start_pulse_r) begin
    st_dma_start_pulse_r <= 1'h0;
  end
  else st_dma_start_pulse_r <= st_dma_start_pulse_next;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    cycle_count <= 16'h0;
  end
  else if (st_dma_start_pulse_r) begin
    cycle_count <= 16'h0;
  end
  else if (loop_done_muxed) begin
    cycle_count <= 16'h0;
  end
  else if (cycle_counter_en & strm_run) begin
    cycle_count <= cycle_count + 16'h1;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    data_f2g_r <= 32'h0;
    data_f2g_vld_r <= 2'h0;
    ctrl_f2g_r <= 2'h0;
  end
  else begin
    data_f2g_r[0] <= data_f2g[0];
    data_f2g_r[1] <= data_f2g[1];
    data_f2g_vld_r <= data_f2g_vld;
    ctrl_f2g_r <= ctrl_f2g;
  end
end
always_comb begin
  strm_data = 16'h0;
  strm_data_valid = 1'h0;
  if (cfg_data_network_f2g_mux[0] == 1'h1) begin
    strm_data = data_f2g_r[0];
    data_f2g_rdy[0] = data_ready_g2f_w;
    if (rv_mode_on) begin
      strm_data_valid = data_f2g_vld_r[0];
    end
    else strm_data_valid = ctrl_f2g_r[0];
  end
  else begin
    strm_data = strm_data;
    strm_data_valid = strm_data_valid;
    data_f2g_rdy[0] = 1'h0;
  end
  if (cfg_data_network_f2g_mux[1] == 1'h1) begin
    strm_data = data_f2g_r[1];
    data_f2g_rdy[1] = data_ready_g2f_w;
    if (rv_mode_on) begin
      strm_data_valid = data_f2g_vld_r[1];
    end
    else strm_data_valid = ctrl_f2g_r[1];
  end
  else begin
    strm_data = strm_data;
    strm_data_valid = strm_data_valid;
    data_f2g_rdy[1] = 1'h0;
  end
end
always_comb begin
  if (cycle_counter_en) begin
    iter_step_valid = cycle_valid;
  end
  else if (rv_mode_on) begin
    iter_step_valid = strm_run & fifo_pop_ready;
  end
  else iter_step_valid = strm_data_valid;
end
always_comb begin
  strm_wr_en_w = iter_step_valid;
  if (rv_mode_on) begin
    strm_wr_addr_w = 19'(data_current_addr);
    strm_wr_data_w = data_fifo2dma;
  end
  else begin
    strm_wr_addr_w = 19'(data_current_addr);
    strm_wr_data_w = strm_data;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    last_strm_wr_addr_r <= 19'h0;
  end
  else if (strm_wr_en_w) begin
    last_strm_wr_addr_r <= strm_wr_addr_w;
  end
end
always_comb begin
  strm_data_sel = strm_wr_addr_w[2:1];
end
always_comb begin
  bank_wr_strb_cache_w = bank_wr_strb_cache_r;
  bank_wr_data_cache_w = bank_wr_data_cache_r;
  if (bank_wr_en) begin
    bank_wr_strb_cache_w = 8'h0;
    bank_wr_data_cache_w = 64'h0;
  end
  if (strm_wr_en_w) begin
    if (strm_data_sel == 2'h0) begin
      bank_wr_strb_cache_w[1:0] = 2'h3;
      bank_wr_data_cache_w[15:0] = strm_wr_data_w;
    end
    else if (strm_data_sel == 2'h1) begin
      bank_wr_strb_cache_w[3:2] = 2'h3;
      bank_wr_data_cache_w[31:16] = strm_wr_data_w;
    end
    else if (strm_data_sel == 2'h2) begin
      bank_wr_strb_cache_w[5:4] = 2'h3;
      bank_wr_data_cache_w[47:32] = strm_wr_data_w;
    end
    else if (strm_data_sel == 2'h3) begin
      bank_wr_strb_cache_w[7:6] = 2'h3;
      bank_wr_data_cache_w[63:48] = strm_wr_data_w;
    end
    else begin
      bank_wr_strb_cache_w = bank_wr_strb_cache_r;
      bank_wr_data_cache_w = bank_wr_data_cache_r;
    end
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    bank_wr_strb_cache_r <= 8'h0;
    bank_wr_data_cache_r <= 64'h0;
  end
  else begin
    bank_wr_strb_cache_r <= bank_wr_strb_cache_w;
    bank_wr_data_cache_r <= bank_wr_data_cache_w;
  end
end
always_comb begin
  bank_addr_match = strm_wr_addr_w[18:3] == last_strm_wr_addr_r[18:3];
  bank_wr_en = (strm_wr_en_w & (~bank_addr_match) & (~is_first)) | is_last;
  bank_wr_addr = last_strm_wr_addr_r;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    wr_packet_dma2bank <= 92'h0;
    wr_packet_dma2ring <= 92'h0;
  end
  else begin
    wr_packet_dma2bank <= wr_packet_dma2bank_w;
    wr_packet_dma2ring <= wr_packet_dma2ring_w;
  end
end
always_comb begin
  if (cfg_tile_connected_next | cfg_tile_connected_prev) begin
    wr_packet_dma2bank_w = 92'h0;
    wr_packet_dma2ring_w.wr_en = bank_wr_en;
    wr_packet_dma2ring_w.wr_strb = bank_wr_strb_cache_r;
    wr_packet_dma2ring_w.wr_data = bank_wr_data_cache_r;
    wr_packet_dma2ring_w.wr_addr = bank_wr_addr;
  end
  else begin
    wr_packet_dma2bank_w.wr_en = bank_wr_en;
    wr_packet_dma2bank_w.wr_strb = bank_wr_strb_cache_r;
    wr_packet_dma2bank_w.wr_data = bank_wr_data_cache_r;
    wr_packet_dma2bank_w.wr_addr = bank_wr_addr;
    wr_packet_dma2ring_w = 92'h0;
  end
end
assign clk_en_dma2bank = dma2bank_clk_en;
always_comb begin
  done_pulse_w = loop_done_muxed & strm_run;
end
assign st_dma_done_pulse = done_pulse_d_arr[5'(cfg_data_network_latency) + 5'h1];

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    st_dma_done_interrupt <= 1'h0;
  end
  else if (st_dma_done_pulse) begin
    st_dma_done_interrupt <= 1'h1;
  end
  else if (st_dma_done_pulse_last) begin
    st_dma_done_interrupt <= 1'h0;
  end
end
always_comb begin
  if (rv_mode_on) begin
    block_done = strm_run & (~rv_is_metadata) & (((rv_num_data_cnt == 16'h1) & fifo_pop_ready) |
        (rv_num_data_cnt == 16'h0));
  end
  else block_done = 1'h0;
end
always_comb begin
  if (rv_mode_on) begin
    loop_done_muxed = block_done & is_last_block;
  end
  else loop_done_muxed = loop_done;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    rv_num_blocks_cnt <= 32'h0;
  end
  else if (rv_mode_on) begin
    if (st_dma_start_pulse_r) begin
      rv_num_blocks_cnt <= cfg_st_dma_num_blocks;
    end
    else if (block_done & (rv_num_blocks_cnt > 32'h0)) begin
      rv_num_blocks_cnt <= rv_num_blocks_cnt - 32'h1;
    end
  end
end
always_comb begin
  is_last_block = rv_num_blocks_cnt == 32'h1;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    rv_is_metadata <= 1'h0;
  end
  else if (rv_mode_on) begin
    if (st_dma_start_pulse_r) begin
      rv_is_metadata <= 1'h1;
    end
    else if (rv_mode_on & block_done & (~is_last_block)) begin
      rv_is_metadata <= 1'h1;
    end
    else if (rv_is_metadata & fifo_pop_ready) begin
      rv_is_metadata <= 1'h0;
    end
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    rv_num_data_cnt <= 16'h0;
  end
  else if (st_dma_start_pulse_r) begin
    rv_num_data_cnt <= 16'h0;
  end
  else if (strm_run & rv_is_metadata & fifo_pop_ready) begin
    rv_num_data_cnt <= data_fifo2dma;
  end
  else if ((rv_num_data_cnt > 16'h0) & fifo_pop_ready) begin
    rv_num_data_cnt <= rv_num_data_cnt - 16'h1;
  end
end
always_comb begin
  if (rv_mode_on) begin
    data_ready_g2f_w = fifo2cgra_ready;
  end
  else data_ready_g2f_w = 1'h0;
end
assign rv_mode_on = cfg_st_dma_ctrl_valid_mode == 2'h1;
assign data_cgra2fifo = strm_data;
assign fifo_pop_ready = ~fifo_empty;
assign fifo_pop = (~fifo_empty) & strm_run;
assign fifo_push = (~fifo_full) & strm_data_valid;
assign fifo2cgra_ready = ~fifo_almost_full;
assign loop_iter_ranges[0] = current_dma_header.range_0;
assign loop_iter_ranges[1] = current_dma_header.range_1;
assign loop_iter_ranges[2] = current_dma_header.range_2;
assign loop_iter_ranges[3] = current_dma_header.range_3;
assign loop_iter_ranges[4] = current_dma_header.range_4;
assign loop_iter_ranges[5] = current_dma_header.range_5;
assign loop_iter_ranges[6] = current_dma_header.range_6;
assign cycle_counter_en = cfg_st_dma_ctrl_valid_mode == 2'h2;
assign cycle_stride_addr_gen_strides[0] = current_dma_header.cycle_stride_0;
assign cycle_stride_addr_gen_strides[1] = current_dma_header.cycle_stride_1;
assign cycle_stride_addr_gen_strides[2] = current_dma_header.cycle_stride_2;
assign cycle_stride_addr_gen_strides[3] = current_dma_header.cycle_stride_3;
assign cycle_stride_addr_gen_strides[4] = current_dma_header.cycle_stride_4;
assign cycle_stride_addr_gen_strides[5] = current_dma_header.cycle_stride_5;
assign cycle_stride_addr_gen_strides[6] = current_dma_header.cycle_stride_6;
assign data_stride_addr_gen_start_addr = 20'(current_dma_header.start_addr);
assign data_stride_addr_gen_strides[0] = current_dma_header.stride_0;
assign data_stride_addr_gen_strides[1] = current_dma_header.stride_1;
assign data_stride_addr_gen_strides[2] = current_dma_header.stride_2;
assign data_stride_addr_gen_strides[3] = current_dma_header.stride_3;
assign data_stride_addr_gen_strides[4] = current_dma_header.stride_4;
assign data_stride_addr_gen_strides[5] = current_dma_header.stride_5;
assign data_stride_addr_gen_strides[6] = current_dma_header.stride_6;
glb_clk_en_gen_4 #(
  .cnt(32'h4))
dma2bank_clk_en_gen (
  .clk(clk),
  .enable(wr_packet_dma2bank_w.wr_en),
  .reset(reset),
  .clk_en(dma2bank_clk_en)
);

pipeline_w_1_d_20_array done_pulse_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(done_pulse_w),
  .reset(reset),
  .out_(done_pulse_d_arr)
);

pipeline_w_1_d_5 st_dma_interrupt_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(st_dma_done_pulse),
  .reset(reset),
  .out_(st_dma_done_pulse_last)
);

reg_fifo_d_4_w_16 #(
  .data_width(16'h10))
data_f2g_fifo (
  .almost_empty_diff(2'h2),
  .almost_full_diff(2'h2),
  .clk(clk),
  .clk_en(rv_mode_on),
  .data_in(data_cgra2fifo),
  .flush(st_dma_start_pulse_r),
  .pop(fifo_pop),
  .push(fifo_push),
  .reset(reset),
  .almost_full(fifo_almost_full),
  .data_out(data_fifo2dma),
  .empty(fifo_empty),
  .full(fifo_full)
);

glb_loop_iter_7 loop_iter (
  .clk(clk),
  .clk_en(1'h1),
  .dim(current_dma_header.dim),
  .ranges(loop_iter_ranges),
  .reset(reset),
  .step(iter_step_valid),
  .mux_sel_out(loop_mux_sel),
  .restart(loop_done)
);

glb_sched_gen cycle_stride_sched_gen (
  .clk(clk),
  .clk_en(cycle_counter_en),
  .current_addr(cycle_current_addr),
  .cycle_count(cycle_count),
  .finished(loop_done_muxed),
  .reset(reset),
  .restart(st_dma_start_pulse_r),
  .valid_output(cycle_valid)
);

glb_addr_gen_7 #(
  .addr_width(32'h10),
  .loop_level(32'h7))
cycle_stride_addr_gen (
  .clk(clk),
  .clk_en(cycle_counter_en),
  .mux_sel(loop_mux_sel),
  .reset(reset),
  .restart(st_dma_start_pulse_r),
  .start_addr(current_dma_header.cycle_start_addr),
  .step(iter_step_valid),
  .strides(cycle_stride_addr_gen_strides),
  .addr_out(cycle_current_addr)
);

glb_addr_gen_7 #(
  .addr_width(32'h14),
  .loop_level(32'h7))
data_stride_addr_gen (
  .clk(clk),
  .clk_en(1'h1),
  .mux_sel(loop_mux_sel),
  .reset(reset),
  .restart(st_dma_start_pulse_r),
  .start_addr(data_stride_addr_gen_start_addr),
  .step(iter_step_valid),
  .strides(data_stride_addr_gen_strides),
  .addr_out(data_current_addr)
);

endmodule   // glb_store_dma

module glb_switch (
  glb_tile_ifc_A_19_D_64.master if_est_m,
  glb_tile_ifc_A_19_D_64.slave if_wst_s,
  input logic gclk,
  input logic glb_tile_id,
  input logic mclk,
  input rdrs_packet_t rdrs_packet,
  input logic reset,
  output logic clk_en_sw2bank,
  output rdrq_packet_t rdrq_packet,
  output wr_packet_t wr_packet
);

logic [18:0] bank_rd_addr;
logic bank_rd_en;
logic [18:0] bank_wr_addr;
logic [63:0] bank_wr_data;
logic bank_wr_en;
logic [7:0] bank_wr_strb;
logic [18:0] if_est_m_rd_addr_w;
logic if_est_m_rd_clk_en_sel;
logic if_est_m_rd_clk_en_sel_first_cycle;
logic if_est_m_rd_clk_en_sel_latch;
logic if_est_m_rd_en_w;
logic [18:0] if_est_m_wr_addr_w;
logic if_est_m_wr_clk_en_sel;
logic if_est_m_wr_clk_en_sel_first_cycle;
logic if_est_m_wr_clk_en_sel_latch;
logic [63:0] if_est_m_wr_data_w;
logic if_est_m_wr_en_w;
logic [7:0] if_est_m_wr_strb_w;
logic if_wst_s_rd_clk_en_d;
logic if_wst_s_wr_clk_en_d;
logic rd_data_valid_w;
logic [63:0] rd_data_w;
logic rd_tile_id_match;
logic sw2bank_rd_clk_en;
logic sw2bank_rd_clk_en_gen_enable;
logic sw2bank_wr_clk_en;
logic sw2bank_wr_clk_en_gen_enable;
logic wr_tile_id_match;
always_comb begin
  wr_tile_id_match = glb_tile_id == if_wst_s.wr_addr[18];
  rd_tile_id_match = glb_tile_id == if_wst_s.rd_addr[18];
end
always_comb begin
  if (if_wst_s.wr_en) begin
    if (wr_tile_id_match) begin
      if_est_m_wr_en_w = 1'h0;
      if_est_m_wr_addr_w = 19'h0;
      if_est_m_wr_data_w = 64'h0;
      if_est_m_wr_strb_w = 8'h0;
      bank_wr_en = 1'h1;
      bank_wr_addr = if_wst_s.wr_addr;
      bank_wr_data = if_wst_s.wr_data;
      bank_wr_strb = if_wst_s.wr_strb;
    end
    else begin
      if_est_m_wr_en_w = if_wst_s.wr_en;
      if_est_m_wr_addr_w = if_wst_s.wr_addr;
      if_est_m_wr_data_w = if_wst_s.wr_data;
      if_est_m_wr_strb_w = if_wst_s.wr_strb;
      bank_wr_en = 1'h0;
      bank_wr_addr = 19'h0;
      bank_wr_data = 64'h0;
      bank_wr_strb = 8'h0;
    end
  end
  else begin
    if_est_m_wr_en_w = 1'h0;
    if_est_m_wr_addr_w = 19'h0;
    if_est_m_wr_data_w = 64'h0;
    if_est_m_wr_strb_w = 8'h0;
    bank_wr_en = 1'h0;
    bank_wr_addr = 19'h0;
    bank_wr_data = 64'h0;
    bank_wr_strb = 8'h0;
  end
end
always_comb begin
  if (if_wst_s.rd_en) begin
    if (rd_tile_id_match) begin
      if_est_m_rd_en_w = 1'h0;
      if_est_m_rd_addr_w = 19'h0;
      bank_rd_en = 1'h1;
      bank_rd_addr = if_wst_s.rd_addr;
    end
    else begin
      if_est_m_rd_en_w = if_wst_s.rd_en;
      if_est_m_rd_addr_w = if_wst_s.rd_addr;
      bank_rd_en = 1'h0;
      bank_rd_addr = 19'h0;
    end
  end
  else begin
    if_est_m_rd_en_w = 1'h0;
    if_est_m_rd_addr_w = 19'h0;
    bank_rd_en = 1'h0;
    bank_rd_addr = 19'h0;
  end
end
always_comb begin
  rd_data_w = 64'h0;
  rd_data_valid_w = 1'h0;
  if (rdrs_packet.rd_data_valid == 1'h1) begin
    rd_data_w = rdrs_packet.rd_data;
    rd_data_valid_w = 1'h1;
  end
  else if (if_est_m.rd_data_valid == 1'h1) begin
    rd_data_w = if_est_m.rd_data;
    rd_data_valid_w = 1'h1;
  end
end

always_ff @(posedge gclk, posedge reset) begin
  if (reset) begin
    if_est_m.wr_en <= 1'h0;
    if_est_m.wr_strb <= 8'h0;
    if_est_m.wr_addr <= 19'h0;
    if_est_m.wr_data <= 64'h0;
    if_est_m.rd_en <= 1'h0;
    if_est_m.rd_addr <= 19'h0;
    if_wst_s.rd_data <= 64'h0;
    if_wst_s.rd_data_valid <= 1'h0;
    wr_packet.wr_en <= 1'h0;
    wr_packet.wr_strb <= 8'h0;
    wr_packet.wr_addr <= 19'h0;
    wr_packet.wr_data <= 64'h0;
    rdrq_packet.rd_en <= 1'h0;
    rdrq_packet.rd_addr <= 19'h0;
  end
  else begin
    if_est_m.wr_en <= if_est_m_wr_en_w;
    if_est_m.wr_strb <= if_est_m_wr_strb_w;
    if_est_m.wr_addr <= if_est_m_wr_addr_w;
    if_est_m.wr_data <= if_est_m_wr_data_w;
    if_est_m.rd_en <= if_est_m_rd_en_w;
    if_est_m.rd_addr <= if_est_m_rd_addr_w;
    if_wst_s.rd_data <= rd_data_w;
    if_wst_s.rd_data_valid <= rd_data_valid_w;
    wr_packet.wr_en <= bank_wr_en;
    wr_packet.wr_strb <= bank_wr_strb;
    wr_packet.wr_addr <= bank_wr_addr;
    wr_packet.wr_data <= bank_wr_data;
    rdrq_packet.rd_en <= bank_rd_en;
    rdrq_packet.rd_addr <= bank_rd_addr;
  end
end

always_ff @(posedge mclk, posedge reset) begin
  if (reset) begin
    if_wst_s_wr_clk_en_d <= 1'h0;
    if_wst_s_rd_clk_en_d <= 1'h0;
  end
  else begin
    if_wst_s_wr_clk_en_d <= if_wst_s.wr_clk_en;
    if_wst_s_rd_clk_en_d <= if_wst_s.rd_clk_en;
  end
end
always_comb begin
  if_est_m_wr_clk_en_sel_first_cycle = if_wst_s.wr_en & (~wr_tile_id_match);
  if_est_m_rd_clk_en_sel_first_cycle = if_wst_s.rd_en & (~rd_tile_id_match);
end

always_ff @(posedge mclk, posedge reset) begin
  if (reset) begin
    if_est_m_wr_clk_en_sel_latch <= 1'h0;
  end
  else if (if_wst_s.wr_en == 1'h1) begin
    if (wr_tile_id_match) begin
      if_est_m_wr_clk_en_sel_latch <= 1'h0;
    end
    else if_est_m_wr_clk_en_sel_latch <= 1'h1;
  end
  else if (if_wst_s.wr_clk_en == 1'h0) begin
    if_est_m_wr_clk_en_sel_latch <= 1'h0;
  end
end

always_ff @(posedge mclk, posedge reset) begin
  if (reset) begin
    if_est_m_rd_clk_en_sel_latch <= 1'h0;
  end
  else if (if_wst_s.rd_en == 1'h1) begin
    if (rd_tile_id_match) begin
      if_est_m_rd_clk_en_sel_latch <= 1'h0;
    end
    else if_est_m_rd_clk_en_sel_latch <= 1'h1;
  end
  else if (if_wst_s.rd_clk_en == 1'h0) begin
    if_est_m_rd_clk_en_sel_latch <= 1'h0;
  end
end
always_comb begin
  if_est_m_wr_clk_en_sel = if_est_m_wr_clk_en_sel_first_cycle | if_est_m_wr_clk_en_sel_latch;
  if_est_m_rd_clk_en_sel = if_est_m_rd_clk_en_sel_first_cycle | if_est_m_rd_clk_en_sel_latch;
end
always_comb begin
  if (if_est_m_wr_clk_en_sel) begin
    if_est_m.wr_clk_en = if_wst_s_wr_clk_en_d;
  end
  else if_est_m.wr_clk_en = 1'h0;
end
always_comb begin
  if (if_est_m_rd_clk_en_sel) begin
    if_est_m.rd_clk_en = if_wst_s_rd_clk_en_d;
  end
  else if_est_m.rd_clk_en = 1'h0;
end
assign sw2bank_wr_clk_en_gen_enable = if_wst_s.wr_en & wr_tile_id_match;
assign sw2bank_rd_clk_en_gen_enable = if_wst_s.rd_en & rd_tile_id_match;
assign clk_en_sw2bank = sw2bank_wr_clk_en | sw2bank_rd_clk_en;
glb_clk_en_gen_4 #(
  .cnt(32'h4))
sw2bank_wr_clk_en_gen (
  .clk(mclk),
  .enable(sw2bank_wr_clk_en_gen_enable),
  .reset(reset),
  .clk_en(sw2bank_wr_clk_en)
);

glb_clk_en_gen_6 #(
  .cnt(32'h6))
sw2bank_rd_clk_en_gen (
  .clk(mclk),
  .enable(sw2bank_rd_clk_en_gen_enable),
  .reset(reset),
  .clk_en(sw2bank_rd_clk_en)
);

endmodule   // glb_switch

module glb_tile (
  input logic cfg_pcfg_tile_connected_wsti,
  input logic cfg_tile_connected_wsti,
  input logic [31:0] cgra_cfg_jtag_addr_bypass_wsti,
  input logic [31:0] cgra_cfg_jtag_addr_wsti,
  input logic [31:0] cgra_cfg_jtag_data_wsti,
  input logic cgra_cfg_jtag_rd_en_bypass_wsti,
  input logic cgra_cfg_jtag_rd_en_wsti,
  input logic cgra_cfg_jtag_wr_en_wsti,
  input logic [31:0] cgra_cfg_pcfg_addr_e2w_esti,
  input logic [31:0] cgra_cfg_pcfg_addr_w2e_wsti,
  input logic [31:0] cgra_cfg_pcfg_data_e2w_esti,
  input logic [31:0] cgra_cfg_pcfg_data_w2e_wsti,
  input logic cgra_cfg_pcfg_rd_en_e2w_esti,
  input logic cgra_cfg_pcfg_rd_en_w2e_wsti,
  input logic cgra_cfg_pcfg_wr_en_e2w_esti,
  input logic cgra_cfg_pcfg_wr_en_w2e_wsti,
  input logic clk,
  input logic clk_en_bank_master,
  input logic clk_en_master,
  input logic clk_en_pcfg_broadcast,
  input logic glb_tile_id,
  input logic [31:0] if_cfg_est_m_rd_data,
  input logic if_cfg_est_m_rd_data_valid,
  input logic [11:0] if_cfg_wst_s_rd_addr,
  input logic if_cfg_wst_s_rd_clk_en,
  input logic if_cfg_wst_s_rd_en,
  input logic [11:0] if_cfg_wst_s_wr_addr,
  input logic if_cfg_wst_s_wr_clk_en,
  input logic [31:0] if_cfg_wst_s_wr_data,
  input logic if_cfg_wst_s_wr_en,
  input logic [63:0] if_proc_est_m_rd_data,
  input logic if_proc_est_m_rd_data_valid,
  input logic [18:0] if_proc_wst_s_rd_addr,
  input logic if_proc_wst_s_rd_clk_en,
  input logic if_proc_wst_s_rd_en,
  input logic [18:0] if_proc_wst_s_wr_addr,
  input logic if_proc_wst_s_wr_clk_en,
  input logic [63:0] if_proc_wst_s_wr_data,
  input logic if_proc_wst_s_wr_en,
  input logic [7:0] if_proc_wst_s_wr_strb,
  input logic [18:0] pcfg_rd_addr_e2w_esti,
  input logic [18:0] pcfg_rd_addr_w2e_wsti,
  input logic [63:0] pcfg_rd_data_e2w_esti,
  input logic pcfg_rd_data_valid_e2w_esti,
  input logic pcfg_rd_data_valid_w2e_wsti,
  input logic [63:0] pcfg_rd_data_w2e_wsti,
  input logic pcfg_rd_en_e2w_esti,
  input logic pcfg_rd_en_w2e_wsti,
  input logic pcfg_start_pulse,
  input logic reset,
  input logic [1:0] strm_ctrl_f2g,
  input logic [1:0] [15:0] strm_data_f2g,
  input logic [1:0] strm_data_f2g_vld,
  input logic [1:0] strm_data_g2f_rdy,
  input logic strm_f2g_start_pulse,
  input logic strm_g2f_start_pulse,
  input logic [18:0] strm_rd_addr_e2w_esti,
  input logic [18:0] strm_rd_addr_w2e_wsti,
  input logic [63:0] strm_rd_data_e2w_esti,
  input logic strm_rd_data_valid_e2w_esti,
  input logic strm_rd_data_valid_w2e_wsti,
  input logic [63:0] strm_rd_data_w2e_wsti,
  input logic strm_rd_en_e2w_esti,
  input logic strm_rd_en_w2e_wsti,
  input logic [18:0] strm_wr_addr_e2w_esti,
  input logic [18:0] strm_wr_addr_w2e_wsti,
  input logic [63:0] strm_wr_data_e2w_esti,
  input logic [63:0] strm_wr_data_w2e_wsti,
  input logic strm_wr_en_e2w_esti,
  input logic strm_wr_en_w2e_wsti,
  input logic [7:0] strm_wr_strb_e2w_esti,
  input logic [7:0] strm_wr_strb_w2e_wsti,
  output logic cfg_pcfg_tile_connected_esto,
  output logic cfg_tile_connected_esto,
  output logic [1:0] [31:0] cgra_cfg_g2f_cfg_addr,
  output logic [1:0] [31:0] cgra_cfg_g2f_cfg_data,
  output logic [1:0] cgra_cfg_g2f_cfg_rd_en,
  output logic [1:0] cgra_cfg_g2f_cfg_wr_en,
  output logic [31:0] cgra_cfg_jtag_addr_bypass_esto,
  output logic [31:0] cgra_cfg_jtag_addr_esto,
  output logic [31:0] cgra_cfg_jtag_data_esto,
  output logic cgra_cfg_jtag_rd_en_bypass_esto,
  output logic cgra_cfg_jtag_rd_en_esto,
  output logic cgra_cfg_jtag_wr_en_esto,
  output logic [31:0] cgra_cfg_pcfg_addr_e2w_wsto,
  output logic [31:0] cgra_cfg_pcfg_addr_w2e_esto,
  output logic [31:0] cgra_cfg_pcfg_data_e2w_wsto,
  output logic [31:0] cgra_cfg_pcfg_data_w2e_esto,
  output logic cgra_cfg_pcfg_rd_en_e2w_wsto,
  output logic cgra_cfg_pcfg_rd_en_w2e_esto,
  output logic cgra_cfg_pcfg_wr_en_e2w_wsto,
  output logic cgra_cfg_pcfg_wr_en_w2e_esto,
  output logic data_flush,
  output logic [11:0] if_cfg_est_m_rd_addr,
  output logic if_cfg_est_m_rd_clk_en,
  output logic if_cfg_est_m_rd_en,
  output logic [11:0] if_cfg_est_m_wr_addr,
  output logic if_cfg_est_m_wr_clk_en,
  output logic [31:0] if_cfg_est_m_wr_data,
  output logic if_cfg_est_m_wr_en,
  output logic [31:0] if_cfg_wst_s_rd_data,
  output logic if_cfg_wst_s_rd_data_valid,
  output logic [18:0] if_proc_est_m_rd_addr,
  output logic if_proc_est_m_rd_clk_en,
  output logic if_proc_est_m_rd_en,
  output logic [18:0] if_proc_est_m_wr_addr,
  output logic if_proc_est_m_wr_clk_en,
  output logic [63:0] if_proc_est_m_wr_data,
  output logic if_proc_est_m_wr_en,
  output logic [7:0] if_proc_est_m_wr_strb,
  output logic [63:0] if_proc_wst_s_rd_data,
  output logic if_proc_wst_s_rd_data_valid,
  output logic pcfg_g2f_interrupt_pulse,
  output logic [18:0] pcfg_rd_addr_e2w_wsto,
  output logic [18:0] pcfg_rd_addr_w2e_esto,
  output logic [63:0] pcfg_rd_data_e2w_wsto,
  output logic pcfg_rd_data_valid_e2w_wsto,
  output logic pcfg_rd_data_valid_w2e_esto,
  output logic [63:0] pcfg_rd_data_w2e_esto,
  output logic pcfg_rd_en_e2w_wsto,
  output logic pcfg_rd_en_w2e_esto,
  output logic [1:0] strm_ctrl_g2f,
  output logic [1:0] strm_data_f2g_rdy,
  output logic [1:0] [15:0] strm_data_g2f,
  output logic [1:0] strm_data_g2f_vld,
  output logic strm_f2g_interrupt_pulse,
  output logic strm_g2f_interrupt_pulse,
  output logic [18:0] strm_rd_addr_e2w_wsto,
  output logic [18:0] strm_rd_addr_w2e_esto,
  output logic [63:0] strm_rd_data_e2w_wsto,
  output logic strm_rd_data_valid_e2w_wsto,
  output logic strm_rd_data_valid_w2e_esto,
  output logic [63:0] strm_rd_data_w2e_esto,
  output logic strm_rd_en_e2w_wsto,
  output logic strm_rd_en_w2e_esto,
  output logic [18:0] strm_wr_addr_e2w_wsto,
  output logic [18:0] strm_wr_addr_w2e_esto,
  output logic [63:0] strm_wr_data_e2w_wsto,
  output logic [63:0] strm_wr_data_w2e_esto,
  output logic strm_wr_en_e2w_wsto,
  output logic strm_wr_en_w2e_esto,
  output logic [7:0] strm_wr_strb_e2w_wsto,
  output logic [7:0] strm_wr_strb_w2e_esto
);

load_dma_ctrl_t cfg_ld_dma_ctrl;
load_dma_header_t cfg_ld_dma_header;
pcfg_broadcast_mux_t cfg_pcfg_broadcast_mux;
pcfg_dma_ctrl_t cfg_pcfg_dma_ctrl;
pcfg_dma_header_t cfg_pcfg_dma_header;
logic cfg_pcfg_tile_connected_next;
logic cfg_pcfg_tile_connected_prev;
store_dma_ctrl_t cfg_st_dma_ctrl;
store_dma_header_t cfg_st_dma_header;
logic [31:0] cfg_st_dma_num_blocks;
logic cfg_tile_connected_next;
logic cfg_tile_connected_prev;
cgra_cfg_t [1:0] cgra_cfg_g2f_cfg_w;
cgra_cfg_t cgra_cfg_pcfgdma2mux;
logic clk_en_bank;
logic clk_en_cfg;
logic clk_en_ld_dma;
logic clk_en_lddma2bank;
logic clk_en_pcfg_dma;
logic clk_en_pcfg_switch;
logic clk_en_pcfgdma2bank;
logic clk_en_pcfgring2bank;
logic clk_en_proc_switch;
logic clk_en_procsw2bank;
logic clk_en_ring2bank;
logic clk_en_st_dma;
logic clk_en_stdma2bank;
logic clk_en_strm_switch;
logic gclk_bank;
logic gclk_cfg;
logic gclk_ld_dma;
logic gclk_pcfg_broadcast;
logic gclk_pcfg_dma;
logic gclk_pcfg_switch;
logic gclk_proc_switch;
logic gclk_st_dma;
logic gclk_strm_switch;
rdrs_packet_t glb_bank_0_rdrs_packet;
rdrs_packet_t glb_bank_1_rdrs_packet;
cfg_data_network_t glb_cfg_cfg_data_network;
cfg_pcfg_network_t glb_cfg_cfg_pcfg_network;
logic glb_clk_gate_bank_enable;
logic glb_clk_gate_cfg_enable;
logic glb_clk_gate_ld_dma_enable;
logic glb_clk_gate_pcfg_broadcast_enable;
logic glb_clk_gate_pcfg_dma_enable;
logic glb_clk_gate_pcfg_switch_enable;
logic glb_clk_gate_proc_switch_enable;
logic glb_clk_gate_st_dma_enable;
logic glb_clk_gate_strm_switch_enable;
cgra_cfg_t glb_pcfg_broadcast_cgra_cfg_jtag_esto;
cgra_cfg_t glb_pcfg_broadcast_cgra_cfg_jtag_wsti;
cgra_cfg_t glb_pcfg_broadcast_cgra_cfg_pcfg_esti;
cgra_cfg_t glb_pcfg_broadcast_cgra_cfg_pcfg_esto;
cgra_cfg_t glb_pcfg_broadcast_cgra_cfg_pcfg_wsti;
cgra_cfg_t glb_pcfg_broadcast_cgra_cfg_pcfg_wsto;
logic glb_pcfg_ring_switch_cfg_ld_dma_on;
logic glb_strm_ring_switch_cfg_ld_dma_on;
rdrq_packet_t pcfg_rdrq_packet_e2w_esti;
rdrq_packet_t pcfg_rdrq_packet_e2w_wsto;
rdrq_packet_t pcfg_rdrq_packet_w2e_esto;
rdrq_packet_t pcfg_rdrq_packet_w2e_wsti;
rdrs_packet_t pcfg_rdrs_packet_e2w_esti;
rdrs_packet_t pcfg_rdrs_packet_e2w_wsto;
rdrs_packet_t pcfg_rdrs_packet_w2e_esto;
rdrs_packet_t pcfg_rdrs_packet_w2e_wsti;
rdrq_packet_t rdrq_packet_dma2bank;
rdrq_packet_t rdrq_packet_dma2ring;
rdrq_packet_t rdrq_packet_pcfgdma2bank;
rdrq_packet_t rdrq_packet_pcfgdma2ring;
rdrq_packet_t rdrq_packet_pcfgring2bank;
rdrq_packet_t rdrq_packet_procsw2bank;
rdrq_packet_t rdrq_packet_ring2bank;
rdrq_bank_packet_t [1:0] rdrq_packet_sw2bankarr;
rdrs_packet_t rdrs_packet_bank2dma;
rdrs_packet_t rdrs_packet_bank2pcfgdma;
rdrs_packet_t rdrs_packet_bank2pcfgring;
rdrs_packet_t rdrs_packet_bank2procsw;
rdrs_packet_t rdrs_packet_bank2ring;
rdrs_packet_t [1:0] rdrs_packet_bankarr2sw;
rdrs_packet_t rdrs_packet_pcfgring2dma;
rdrs_packet_t rdrs_packet_ring2dma;
rdrq_packet_t strm_rdrq_packet_e2w_esti;
rdrq_packet_t strm_rdrq_packet_e2w_wsto;
rdrq_packet_t strm_rdrq_packet_w2e_esto;
rdrq_packet_t strm_rdrq_packet_w2e_wsti;
rdrs_packet_t strm_rdrs_packet_e2w_esti;
rdrs_packet_t strm_rdrs_packet_e2w_wsto;
rdrs_packet_t strm_rdrs_packet_w2e_esto;
rdrs_packet_t strm_rdrs_packet_w2e_wsti;
wr_packet_t strm_wr_packet_e2w_esti;
wr_packet_t strm_wr_packet_e2w_wsto;
wr_packet_t strm_wr_packet_w2e_esto;
wr_packet_t strm_wr_packet_w2e_wsti;
wr_packet_t wr_packet_dma2bank;
wr_packet_t wr_packet_dma2ring;
wr_packet_t wr_packet_procsw2bank;
wr_packet_t wr_packet_ring2bank;
wr_bank_packet_t [1:0] wr_packet_sw2bankarr;
glb_tile_ifc_A_12_D_32 if_cfg_est_m();
glb_tile_ifc_A_12_D_32 if_cfg_wst_s();
glb_tile_ifc_A_19_D_64 if_proc_est_m();
glb_tile_ifc_A_19_D_64 if_proc_wst_s();
assign if_proc_est_m_wr_en = if_proc_est_m.wr_en;
assign if_proc_wst_s.wr_en = if_proc_wst_s_wr_en;
assign if_proc_est_m_wr_addr = if_proc_est_m.wr_addr;
assign if_proc_wst_s.wr_addr = if_proc_wst_s_wr_addr;
assign if_proc_est_m_wr_data = if_proc_est_m.wr_data;
assign if_proc_wst_s.wr_data = if_proc_wst_s_wr_data;
assign if_proc_est_m_rd_en = if_proc_est_m.rd_en;
assign if_proc_wst_s.rd_en = if_proc_wst_s_rd_en;
assign if_proc_est_m_rd_addr = if_proc_est_m.rd_addr;
assign if_proc_wst_s.rd_addr = if_proc_wst_s_rd_addr;
assign if_proc_est_m_wr_strb = if_proc_est_m.wr_strb;
assign if_proc_wst_s.wr_strb = if_proc_wst_s_wr_strb;
assign if_proc_est_m_wr_clk_en = if_proc_est_m.wr_clk_en;
assign if_proc_wst_s.wr_clk_en = if_proc_wst_s_wr_clk_en;
assign if_proc_est_m_rd_clk_en = if_proc_est_m.rd_clk_en;
assign if_proc_wst_s.rd_clk_en = if_proc_wst_s_rd_clk_en;
assign if_proc_est_m.rd_data = if_proc_est_m_rd_data;
assign if_proc_wst_s_rd_data = if_proc_wst_s.rd_data;
assign if_proc_est_m.rd_data_valid = if_proc_est_m_rd_data_valid;
assign if_proc_wst_s_rd_data_valid = if_proc_wst_s.rd_data_valid;
assign if_cfg_est_m_wr_en = if_cfg_est_m.wr_en;
assign if_cfg_wst_s.wr_en = if_cfg_wst_s_wr_en;
assign if_cfg_est_m_wr_addr = if_cfg_est_m.wr_addr;
assign if_cfg_wst_s.wr_addr = if_cfg_wst_s_wr_addr;
assign if_cfg_est_m_wr_data = if_cfg_est_m.wr_data;
assign if_cfg_wst_s.wr_data = if_cfg_wst_s_wr_data;
assign if_cfg_est_m_rd_en = if_cfg_est_m.rd_en;
assign if_cfg_wst_s.rd_en = if_cfg_wst_s_rd_en;
assign if_cfg_est_m_rd_addr = if_cfg_est_m.rd_addr;
assign if_cfg_wst_s.rd_addr = if_cfg_wst_s_rd_addr;
assign if_cfg_est_m_wr_clk_en = if_cfg_est_m.wr_clk_en;
assign if_cfg_wst_s.wr_clk_en = if_cfg_wst_s_wr_clk_en;
assign if_cfg_est_m_rd_clk_en = if_cfg_est_m.rd_clk_en;
assign if_cfg_wst_s.rd_clk_en = if_cfg_wst_s_rd_clk_en;
assign if_cfg_est_m.rd_data = if_cfg_est_m_rd_data;
assign if_cfg_wst_s_rd_data = if_cfg_wst_s.rd_data;
assign if_cfg_est_m.rd_data_valid = if_cfg_est_m_rd_data_valid;
assign if_cfg_wst_s_rd_data_valid = if_cfg_wst_s.rd_data_valid;
assign strm_wr_packet_w2e_wsti.wr_en = strm_wr_en_w2e_wsti;
assign strm_wr_packet_w2e_wsti.wr_strb = strm_wr_strb_w2e_wsti;
assign strm_wr_packet_w2e_wsti.wr_addr = strm_wr_addr_w2e_wsti;
assign strm_wr_packet_w2e_wsti.wr_data = strm_wr_data_w2e_wsti;
assign strm_wr_en_w2e_esto = strm_wr_packet_w2e_esto.wr_en;
assign strm_wr_strb_w2e_esto = strm_wr_packet_w2e_esto.wr_strb;
assign strm_wr_addr_w2e_esto = strm_wr_packet_w2e_esto.wr_addr;
assign strm_wr_data_w2e_esto = strm_wr_packet_w2e_esto.wr_data;
assign strm_wr_packet_e2w_esti.wr_en = strm_wr_en_e2w_esti;
assign strm_wr_packet_e2w_esti.wr_strb = strm_wr_strb_e2w_esti;
assign strm_wr_packet_e2w_esti.wr_addr = strm_wr_addr_e2w_esti;
assign strm_wr_packet_e2w_esti.wr_data = strm_wr_data_e2w_esti;
assign strm_wr_en_e2w_wsto = strm_wr_packet_e2w_wsto.wr_en;
assign strm_wr_strb_e2w_wsto = strm_wr_packet_e2w_wsto.wr_strb;
assign strm_wr_addr_e2w_wsto = strm_wr_packet_e2w_wsto.wr_addr;
assign strm_wr_data_e2w_wsto = strm_wr_packet_e2w_wsto.wr_data;
assign strm_rdrq_packet_w2e_wsti.rd_en = strm_rd_en_w2e_wsti;
assign strm_rdrq_packet_w2e_wsti.rd_addr = strm_rd_addr_w2e_wsti;
assign strm_rd_en_w2e_esto = strm_rdrq_packet_w2e_esto.rd_en;
assign strm_rd_addr_w2e_esto = strm_rdrq_packet_w2e_esto.rd_addr;
assign strm_rdrq_packet_e2w_esti.rd_en = strm_rd_en_e2w_esti;
assign strm_rdrq_packet_e2w_esti.rd_addr = strm_rd_addr_e2w_esti;
assign strm_rd_en_e2w_wsto = strm_rdrq_packet_e2w_wsto.rd_en;
assign strm_rd_addr_e2w_wsto = strm_rdrq_packet_e2w_wsto.rd_addr;
assign strm_rd_data_e2w_wsto = strm_rdrs_packet_e2w_wsto.rd_data;
assign strm_rd_data_valid_e2w_wsto = strm_rdrs_packet_e2w_wsto.rd_data_valid;
assign strm_rdrs_packet_e2w_esti.rd_data = strm_rd_data_e2w_esti;
assign strm_rdrs_packet_e2w_esti.rd_data_valid = strm_rd_data_valid_e2w_esti;
assign strm_rdrs_packet_w2e_wsti.rd_data = strm_rd_data_w2e_wsti;
assign strm_rdrs_packet_w2e_wsti.rd_data_valid = strm_rd_data_valid_w2e_wsti;
assign strm_rd_data_w2e_esto = strm_rdrs_packet_w2e_esto.rd_data;
assign strm_rd_data_valid_w2e_esto = strm_rdrs_packet_w2e_esto.rd_data_valid;
assign pcfg_rdrq_packet_w2e_wsti.rd_en = pcfg_rd_en_w2e_wsti;
assign pcfg_rdrq_packet_w2e_wsti.rd_addr = pcfg_rd_addr_w2e_wsti;
assign pcfg_rd_en_w2e_esto = pcfg_rdrq_packet_w2e_esto.rd_en;
assign pcfg_rd_addr_w2e_esto = pcfg_rdrq_packet_w2e_esto.rd_addr;
assign pcfg_rdrq_packet_e2w_esti.rd_en = pcfg_rd_en_e2w_esti;
assign pcfg_rdrq_packet_e2w_esti.rd_addr = pcfg_rd_addr_e2w_esti;
assign pcfg_rd_en_e2w_wsto = pcfg_rdrq_packet_e2w_wsto.rd_en;
assign pcfg_rd_addr_e2w_wsto = pcfg_rdrq_packet_e2w_wsto.rd_addr;
assign pcfg_rd_data_e2w_wsto = pcfg_rdrs_packet_e2w_wsto.rd_data;
assign pcfg_rd_data_valid_e2w_wsto = pcfg_rdrs_packet_e2w_wsto.rd_data_valid;
assign pcfg_rdrs_packet_e2w_esti.rd_data = pcfg_rd_data_e2w_esti;
assign pcfg_rdrs_packet_e2w_esti.rd_data_valid = pcfg_rd_data_valid_e2w_esti;
assign pcfg_rdrs_packet_w2e_wsti.rd_data = pcfg_rd_data_w2e_wsti;
assign pcfg_rdrs_packet_w2e_wsti.rd_data_valid = pcfg_rd_data_valid_w2e_wsti;
assign pcfg_rd_data_w2e_esto = pcfg_rdrs_packet_w2e_esto.rd_data;
assign pcfg_rd_data_valid_w2e_esto = pcfg_rdrs_packet_w2e_esto.rd_data_valid;
assign clk_en_cfg = if_cfg_wst_s.wr_clk_en | if_cfg_wst_s.rd_clk_en;
assign glb_clk_gate_cfg_enable = clk_en_cfg | clk_en_master;
assign glb_clk_gate_pcfg_broadcast_enable = clk_en_pcfg_broadcast | clk_en_master;
assign clk_en_ld_dma = cfg_ld_dma_ctrl.mode != 2'h0;
assign glb_clk_gate_ld_dma_enable = clk_en_ld_dma | clk_en_master;
assign clk_en_st_dma = cfg_st_dma_ctrl.mode != 2'h0;
assign glb_clk_gate_st_dma_enable = clk_en_st_dma | clk_en_master;
assign clk_en_proc_switch = if_proc_wst_s.wr_clk_en | if_proc_wst_s.rd_clk_en;
assign glb_clk_gate_proc_switch_enable = clk_en_proc_switch | clk_en_master;
assign clk_en_pcfg_dma = cfg_pcfg_dma_ctrl.mode != 1'h0;
assign glb_clk_gate_pcfg_dma_enable = clk_en_pcfg_dma | clk_en_master;
assign clk_en_strm_switch = cfg_tile_connected_next | cfg_tile_connected_prev;
assign glb_clk_gate_strm_switch_enable = clk_en_strm_switch | clk_en_master;
assign clk_en_pcfg_switch = cfg_pcfg_tile_connected_next | cfg_pcfg_tile_connected_prev;
assign glb_clk_gate_pcfg_switch_enable = clk_en_pcfg_switch | clk_en_master;
assign clk_en_bank = clk_en_lddma2bank | clk_en_stdma2bank | clk_en_pcfgdma2bank | clk_en_ring2bank |
    clk_en_pcfgring2bank | clk_en_procsw2bank;
assign glb_clk_gate_bank_enable = clk_en_bank | clk_en_master | clk_en_bank_master;
assign cfg_tile_connected_next = glb_cfg_cfg_data_network.tile_connected;
assign cfg_tile_connected_prev = cfg_tile_connected_wsti;
assign cfg_tile_connected_esto = cfg_tile_connected_next;
assign cfg_pcfg_tile_connected_next = glb_cfg_cfg_pcfg_network.tile_connected;
assign cfg_pcfg_tile_connected_prev = cfg_pcfg_tile_connected_wsti;
assign cfg_pcfg_tile_connected_esto = cfg_pcfg_tile_connected_next;
assign glb_strm_ring_switch_cfg_ld_dma_on = cfg_ld_dma_ctrl.mode != 2'h0;
assign glb_pcfg_ring_switch_cfg_ld_dma_on = cfg_pcfg_dma_ctrl.mode != 1'h0;
assign rdrs_packet_bankarr2sw[0] = glb_bank_0_rdrs_packet;
assign rdrs_packet_bankarr2sw[1] = glb_bank_1_rdrs_packet;
assign cgra_cfg_g2f_cfg_wr_en[0] = cgra_cfg_g2f_cfg_w[0].wr_en;
assign cgra_cfg_g2f_cfg_rd_en[0] = cgra_cfg_g2f_cfg_w[0].rd_en;
assign cgra_cfg_g2f_cfg_addr[0] = cgra_cfg_g2f_cfg_w[0].addr;
assign cgra_cfg_g2f_cfg_data[0] = cgra_cfg_g2f_cfg_w[0].data;
assign cgra_cfg_g2f_cfg_wr_en[1] = cgra_cfg_g2f_cfg_w[1].wr_en;
assign cgra_cfg_g2f_cfg_rd_en[1] = cgra_cfg_g2f_cfg_w[1].rd_en;
assign cgra_cfg_g2f_cfg_addr[1] = cgra_cfg_g2f_cfg_w[1].addr;
assign cgra_cfg_g2f_cfg_data[1] = cgra_cfg_g2f_cfg_w[1].data;
assign glb_pcfg_broadcast_cgra_cfg_jtag_wsti.wr_en = cgra_cfg_jtag_wr_en_wsti;
assign glb_pcfg_broadcast_cgra_cfg_jtag_wsti.rd_en = cgra_cfg_jtag_rd_en_wsti;
assign glb_pcfg_broadcast_cgra_cfg_jtag_wsti.addr = cgra_cfg_jtag_addr_wsti;
assign glb_pcfg_broadcast_cgra_cfg_jtag_wsti.data = cgra_cfg_jtag_data_wsti;
assign cgra_cfg_jtag_wr_en_esto = glb_pcfg_broadcast_cgra_cfg_jtag_esto.wr_en;
assign cgra_cfg_jtag_rd_en_esto = glb_pcfg_broadcast_cgra_cfg_jtag_esto.rd_en;
assign cgra_cfg_jtag_addr_esto = glb_pcfg_broadcast_cgra_cfg_jtag_esto.addr;
assign cgra_cfg_jtag_data_esto = glb_pcfg_broadcast_cgra_cfg_jtag_esto.data;
assign glb_pcfg_broadcast_cgra_cfg_pcfg_wsti.wr_en = cgra_cfg_pcfg_wr_en_w2e_wsti;
assign glb_pcfg_broadcast_cgra_cfg_pcfg_wsti.rd_en = cgra_cfg_pcfg_rd_en_w2e_wsti;
assign glb_pcfg_broadcast_cgra_cfg_pcfg_wsti.addr = cgra_cfg_pcfg_addr_w2e_wsti;
assign glb_pcfg_broadcast_cgra_cfg_pcfg_wsti.data = cgra_cfg_pcfg_data_w2e_wsti;
assign cgra_cfg_pcfg_wr_en_w2e_esto = glb_pcfg_broadcast_cgra_cfg_pcfg_esto.wr_en;
assign cgra_cfg_pcfg_rd_en_w2e_esto = glb_pcfg_broadcast_cgra_cfg_pcfg_esto.rd_en;
assign cgra_cfg_pcfg_addr_w2e_esto = glb_pcfg_broadcast_cgra_cfg_pcfg_esto.addr;
assign cgra_cfg_pcfg_data_w2e_esto = glb_pcfg_broadcast_cgra_cfg_pcfg_esto.data;
assign glb_pcfg_broadcast_cgra_cfg_pcfg_esti.wr_en = cgra_cfg_pcfg_wr_en_e2w_esti;
assign glb_pcfg_broadcast_cgra_cfg_pcfg_esti.rd_en = cgra_cfg_pcfg_rd_en_e2w_esti;
assign glb_pcfg_broadcast_cgra_cfg_pcfg_esti.addr = cgra_cfg_pcfg_addr_e2w_esti;
assign glb_pcfg_broadcast_cgra_cfg_pcfg_esti.data = cgra_cfg_pcfg_data_e2w_esti;
assign cgra_cfg_pcfg_wr_en_e2w_wsto = glb_pcfg_broadcast_cgra_cfg_pcfg_wsto.wr_en;
assign cgra_cfg_pcfg_rd_en_e2w_wsto = glb_pcfg_broadcast_cgra_cfg_pcfg_wsto.rd_en;
assign cgra_cfg_pcfg_addr_e2w_wsto = glb_pcfg_broadcast_cgra_cfg_pcfg_wsto.addr;
assign cgra_cfg_pcfg_data_e2w_wsto = glb_pcfg_broadcast_cgra_cfg_pcfg_wsto.data;
clk_gate glb_clk_gate_cfg (
  .clk(clk),
  .enable(glb_clk_gate_cfg_enable),
  .gclk(gclk_cfg)
);

clk_gate glb_clk_gate_pcfg_broadcast (
  .clk(clk),
  .enable(glb_clk_gate_pcfg_broadcast_enable),
  .gclk(gclk_pcfg_broadcast)
);

clk_gate glb_clk_gate_ld_dma (
  .clk(clk),
  .enable(glb_clk_gate_ld_dma_enable),
  .gclk(gclk_ld_dma)
);

clk_gate glb_clk_gate_st_dma (
  .clk(clk),
  .enable(glb_clk_gate_st_dma_enable),
  .gclk(gclk_st_dma)
);

clk_gate glb_clk_gate_proc_switch (
  .clk(clk),
  .enable(glb_clk_gate_proc_switch_enable),
  .gclk(gclk_proc_switch)
);

clk_gate glb_clk_gate_pcfg_dma (
  .clk(clk),
  .enable(glb_clk_gate_pcfg_dma_enable),
  .gclk(gclk_pcfg_dma)
);

clk_gate glb_clk_gate_strm_switch (
  .clk(clk),
  .enable(glb_clk_gate_strm_switch_enable),
  .gclk(gclk_strm_switch)
);

clk_gate glb_clk_gate_pcfg_switch (
  .clk(clk),
  .enable(glb_clk_gate_pcfg_switch_enable),
  .gclk(gclk_pcfg_switch)
);

clk_gate glb_clk_gate_bank (
  .clk(clk),
  .enable(glb_clk_gate_bank_enable),
  .gclk(gclk_bank)
);

glb_cfg glb_cfg (
  .gclk(gclk_cfg),
  .glb_tile_id(glb_tile_id),
  .mclk(clk),
  .if_cfg_wst_s(if_cfg_wst_s.slave),
  .if_cfg_est_m(if_cfg_est_m.master),
  .reset(reset),
  .cfg_data_network(glb_cfg_cfg_data_network),
  .cfg_ld_dma_ctrl(cfg_ld_dma_ctrl),
  .cfg_ld_dma_header(cfg_ld_dma_header),
  .cfg_pcfg_broadcast_mux(cfg_pcfg_broadcast_mux),
  .cfg_pcfg_dma_ctrl(cfg_pcfg_dma_ctrl),
  .cfg_pcfg_dma_header(cfg_pcfg_dma_header),
  .cfg_pcfg_network(glb_cfg_cfg_pcfg_network),
  .cfg_st_dma_ctrl(cfg_st_dma_ctrl),
  .cfg_st_dma_header(cfg_st_dma_header),
  .cfg_st_dma_num_blocks(cfg_st_dma_num_blocks)
);

glb_pcfg_broadcast glb_pcfg_broadcast (
  .cfg_pcfg_broadcast_mux(cfg_pcfg_broadcast_mux),
  .cgra_cfg_dma2mux(cgra_cfg_pcfgdma2mux),
  .cgra_cfg_jtag_addr_bypass_wsti(cgra_cfg_jtag_addr_bypass_wsti),
  .cgra_cfg_jtag_rd_en_bypass_wsti(cgra_cfg_jtag_rd_en_bypass_wsti),
  .cgra_cfg_jtag_wsti(glb_pcfg_broadcast_cgra_cfg_jtag_wsti),
  .cgra_cfg_pcfg_esti(glb_pcfg_broadcast_cgra_cfg_pcfg_esti),
  .cgra_cfg_pcfg_wsti(glb_pcfg_broadcast_cgra_cfg_pcfg_wsti),
  .clk(gclk_pcfg_broadcast),
  .reset(reset),
  .cgra_cfg_g2f(cgra_cfg_g2f_cfg_w),
  .cgra_cfg_jtag_addr_bypass_esto(cgra_cfg_jtag_addr_bypass_esto),
  .cgra_cfg_jtag_esto(glb_pcfg_broadcast_cgra_cfg_jtag_esto),
  .cgra_cfg_jtag_rd_en_bypass_esto(cgra_cfg_jtag_rd_en_bypass_esto),
  .cgra_cfg_pcfg_esto(glb_pcfg_broadcast_cgra_cfg_pcfg_esto),
  .cgra_cfg_pcfg_wsto(glb_pcfg_broadcast_cgra_cfg_pcfg_wsto)
);

glb_store_dma glb_store_dma (
  .cfg_data_network_f2g_mux(cfg_st_dma_ctrl.data_mux),
  .cfg_data_network_latency(glb_cfg_cfg_data_network.latency),
  .cfg_st_dma_ctrl_mode(cfg_st_dma_ctrl.mode),
  .cfg_st_dma_ctrl_valid_mode(cfg_st_dma_ctrl.valid_mode),
  .cfg_st_dma_header(cfg_st_dma_header),
  .cfg_st_dma_num_blocks(cfg_st_dma_num_blocks),
  .cfg_st_dma_num_repeat(cfg_st_dma_ctrl.num_repeat),
  .cfg_tile_connected_next(cfg_tile_connected_next),
  .cfg_tile_connected_prev(cfg_tile_connected_prev),
  .clk(gclk_st_dma),
  .ctrl_f2g(strm_ctrl_f2g),
  .data_f2g(strm_data_f2g),
  .data_f2g_vld(strm_data_f2g_vld),
  .reset(reset),
  .st_dma_start_pulse(strm_f2g_start_pulse),
  .clk_en_dma2bank(clk_en_stdma2bank),
  .data_f2g_rdy(strm_data_f2g_rdy),
  .st_dma_done_interrupt(strm_f2g_interrupt_pulse),
  .wr_packet_dma2bank(wr_packet_dma2bank),
  .wr_packet_dma2ring(wr_packet_dma2ring)
);

glb_load_dma glb_load_dma (
  .cfg_data_network_g2f_mux(cfg_ld_dma_ctrl.data_mux),
  .cfg_data_network_latency(glb_cfg_cfg_data_network.latency),
  .cfg_ld_dma_ctrl_flush_mode(cfg_ld_dma_ctrl.flush_mode),
  .cfg_ld_dma_ctrl_mode(cfg_ld_dma_ctrl.mode),
  .cfg_ld_dma_ctrl_valid_mode(cfg_ld_dma_ctrl.valid_mode),
  .cfg_ld_dma_header(cfg_ld_dma_header),
  .cfg_ld_dma_num_repeat(cfg_ld_dma_ctrl.num_repeat),
  .cfg_tile_connected_next(cfg_tile_connected_next),
  .cfg_tile_connected_prev(cfg_tile_connected_prev),
  .clk(gclk_ld_dma),
  .data_g2f_rdy(strm_data_g2f_rdy),
  .glb_tile_id(glb_tile_id),
  .ld_dma_start_pulse(strm_g2f_start_pulse),
  .rdrs_packet_bank2dma(rdrs_packet_bank2dma),
  .rdrs_packet_ring2dma(rdrs_packet_ring2dma),
  .reset(reset),
  .clk_en_dma2bank(clk_en_lddma2bank),
  .ctrl_g2f(strm_ctrl_g2f),
  .data_flush(data_flush),
  .data_g2f(strm_data_g2f),
  .data_g2f_vld(strm_data_g2f_vld),
  .ld_dma_done_interrupt(strm_g2f_interrupt_pulse),
  .rdrq_packet_dma2bank(rdrq_packet_dma2bank),
  .rdrq_packet_dma2ring(rdrq_packet_dma2ring)
);

glb_pcfg_dma glb_pcfg_dma (
  .cfg_pcfg_dma_ctrl_mode(cfg_pcfg_dma_ctrl.mode),
  .cfg_pcfg_dma_ctrl_relocation_is_msb(cfg_pcfg_dma_ctrl.relocation_is_msb),
  .cfg_pcfg_dma_ctrl_relocation_value(cfg_pcfg_dma_ctrl.relocation_value),
  .cfg_pcfg_dma_header(cfg_pcfg_dma_header),
  .cfg_pcfg_network_latency(glb_cfg_cfg_pcfg_network.latency),
  .cfg_pcfg_tile_connected_next(cfg_pcfg_tile_connected_next),
  .cfg_pcfg_tile_connected_prev(cfg_pcfg_tile_connected_prev),
  .clk(gclk_pcfg_dma),
  .glb_tile_id(glb_tile_id),
  .pcfg_dma_start_pulse(pcfg_start_pulse),
  .rdrs_packet_bank2dma(rdrs_packet_bank2pcfgdma),
  .rdrs_packet_ring2dma(rdrs_packet_pcfgring2dma),
  .reset(reset),
  .cgra_cfg_pcfg(cgra_cfg_pcfgdma2mux),
  .clk_en_dma2bank(clk_en_pcfgdma2bank),
  .pcfg_dma_done_interrupt(pcfg_g2f_interrupt_pulse),
  .rdrq_packet_dma2bank(rdrq_packet_pcfgdma2bank),
  .rdrq_packet_dma2ring(rdrq_packet_pcfgdma2ring)
);

glb_bank_mux glb_bank_mux (
  .cfg_pcfg_tile_connected_next(cfg_pcfg_tile_connected_next),
  .cfg_pcfg_tile_connected_prev(cfg_pcfg_tile_connected_prev),
  .cfg_tile_connected_next(cfg_tile_connected_next),
  .cfg_tile_connected_prev(cfg_tile_connected_prev),
  .clk(gclk_bank),
  .glb_tile_id(glb_tile_id),
  .rdrq_packet_dma2bank(rdrq_packet_dma2bank),
  .rdrq_packet_pcfgdma2bank(rdrq_packet_pcfgdma2bank),
  .rdrq_packet_pcfgring2bank(rdrq_packet_pcfgring2bank),
  .rdrq_packet_procsw2bank(rdrq_packet_procsw2bank),
  .rdrq_packet_ring2bank(rdrq_packet_ring2bank),
  .rdrs_packet_bankarr2sw(rdrs_packet_bankarr2sw),
  .reset(reset),
  .wr_packet_dma2bank(wr_packet_dma2bank),
  .wr_packet_procsw2bank(wr_packet_procsw2bank),
  .wr_packet_ring2bank(wr_packet_ring2bank),
  .rdrq_packet_sw2bankarr(rdrq_packet_sw2bankarr),
  .rdrs_packet_bank2dma(rdrs_packet_bank2dma),
  .rdrs_packet_bank2pcfgdma(rdrs_packet_bank2pcfgdma),
  .rdrs_packet_bank2pcfgring(rdrs_packet_bank2pcfgring),
  .rdrs_packet_bank2procsw(rdrs_packet_bank2procsw),
  .rdrs_packet_bank2ring(rdrs_packet_bank2ring),
  .wr_packet_sw2bankarr(wr_packet_sw2bankarr)
);

glb_switch glb_proc_switch (
  .gclk(gclk_proc_switch),
  .glb_tile_id(glb_tile_id),
  .mclk(clk),
  .if_wst_s(if_proc_wst_s.slave),
  .if_est_m(if_proc_est_m.master),
  .rdrs_packet(rdrs_packet_bank2procsw),
  .reset(reset),
  .clk_en_sw2bank(clk_en_procsw2bank),
  .rdrq_packet(rdrq_packet_procsw2bank),
  .wr_packet(wr_packet_procsw2bank)
);

glb_ring_switch_WR_RD glb_strm_ring_switch (
  .cfg_ld_dma_on(glb_strm_ring_switch_cfg_ld_dma_on),
  .cfg_tile_connected_next(cfg_tile_connected_next),
  .cfg_tile_connected_prev(cfg_tile_connected_prev),
  .clk(gclk_strm_switch),
  .glb_tile_id(glb_tile_id),
  .rdrq_packet_dma2ring(rdrq_packet_dma2ring),
  .rdrq_packet_e2w_esti(strm_rdrq_packet_e2w_esti),
  .rdrq_packet_w2e_wsti(strm_rdrq_packet_w2e_wsti),
  .rdrs_packet_bank2ring(rdrs_packet_bank2ring),
  .rdrs_packet_e2w_esti(strm_rdrs_packet_e2w_esti),
  .rdrs_packet_w2e_wsti(strm_rdrs_packet_w2e_wsti),
  .reset(reset),
  .wr_packet_dma2ring(wr_packet_dma2ring),
  .wr_packet_e2w_esti(strm_wr_packet_e2w_esti),
  .wr_packet_w2e_wsti(strm_wr_packet_w2e_wsti),
  .clk_en_ring2bank(clk_en_ring2bank),
  .rdrq_packet_e2w_wsto(strm_rdrq_packet_e2w_wsto),
  .rdrq_packet_ring2bank(rdrq_packet_ring2bank),
  .rdrq_packet_w2e_esto(strm_rdrq_packet_w2e_esto),
  .rdrs_packet_e2w_wsto(strm_rdrs_packet_e2w_wsto),
  .rdrs_packet_ring2dma(rdrs_packet_ring2dma),
  .rdrs_packet_w2e_esto(strm_rdrs_packet_w2e_esto),
  .wr_packet_e2w_wsto(strm_wr_packet_e2w_wsto),
  .wr_packet_ring2bank(wr_packet_ring2bank),
  .wr_packet_w2e_esto(strm_wr_packet_w2e_esto)
);

glb_ring_switch_RD glb_pcfg_ring_switch (
  .cfg_ld_dma_on(glb_pcfg_ring_switch_cfg_ld_dma_on),
  .cfg_tile_connected_next(cfg_pcfg_tile_connected_next),
  .cfg_tile_connected_prev(cfg_pcfg_tile_connected_prev),
  .clk(gclk_pcfg_switch),
  .glb_tile_id(glb_tile_id),
  .rdrq_packet_dma2ring(rdrq_packet_pcfgdma2ring),
  .rdrq_packet_e2w_esti(pcfg_rdrq_packet_e2w_esti),
  .rdrq_packet_w2e_wsti(pcfg_rdrq_packet_w2e_wsti),
  .rdrs_packet_bank2ring(rdrs_packet_bank2pcfgring),
  .rdrs_packet_e2w_esti(pcfg_rdrs_packet_e2w_esti),
  .rdrs_packet_w2e_wsti(pcfg_rdrs_packet_w2e_wsti),
  .reset(reset),
  .clk_en_ring2bank(clk_en_pcfgring2bank),
  .rdrq_packet_e2w_wsto(pcfg_rdrq_packet_e2w_wsto),
  .rdrq_packet_ring2bank(rdrq_packet_pcfgring2bank),
  .rdrq_packet_w2e_esto(pcfg_rdrq_packet_w2e_esto),
  .rdrs_packet_e2w_wsto(pcfg_rdrs_packet_e2w_wsto),
  .rdrs_packet_ring2dma(rdrs_packet_pcfgring2dma),
  .rdrs_packet_w2e_esto(pcfg_rdrs_packet_w2e_esto)
);

glb_bank glb_bank_0 (
  .clk(gclk_bank),
  .rdrq_packet(rdrq_packet_sw2bankarr[0]),
  .reset(reset),
  .wr_packet(wr_packet_sw2bankarr[0]),
  .rdrs_packet(glb_bank_0_rdrs_packet)
);

glb_bank glb_bank_1 (
  .clk(gclk_bank),
  .rdrq_packet(rdrq_packet_sw2bankarr[1]),
  .reset(reset),
  .wr_packet(wr_packet_sw2bankarr[1]),
  .rdrs_packet(glb_bank_1_rdrs_packet)
);

endmodule   // glb_tile

module global_buffer (
  input logic [31:0] cgra_cfg_jtag_gc2glb_addr,
  input logic [31:0] cgra_cfg_jtag_gc2glb_data,
  input logic cgra_cfg_jtag_gc2glb_rd_en,
  input logic cgra_cfg_jtag_gc2glb_wr_en,
  input logic [3:0] cgra_stall_in,
  input logic clk,
  input logic flush_crossbar_sel,
  input logic [1:0] glb_clk_en_bank_master,
  input logic [1:0] glb_clk_en_master,
  input logic [11:0] if_cfg_rd_addr,
  input logic if_cfg_rd_clk_en,
  input logic if_cfg_rd_en,
  input logic [11:0] if_cfg_wr_addr,
  input logic if_cfg_wr_clk_en,
  input logic [31:0] if_cfg_wr_data,
  input logic if_cfg_wr_en,
  input logic [18:0] if_sram_cfg_rd_addr,
  input logic if_sram_cfg_rd_en,
  input logic [18:0] if_sram_cfg_wr_addr,
  input logic [31:0] if_sram_cfg_wr_data,
  input logic if_sram_cfg_wr_en,
  input logic [1:0] pcfg_broadcast_stall,
  input logic [1:0] pcfg_start_pulse,
  input logic [18:0] proc_rd_addr,
  input logic proc_rd_en,
  input logic [18:0] proc_wr_addr,
  input logic [63:0] proc_wr_data,
  input logic proc_wr_en,
  input logic [7:0] proc_wr_strb,
  input logic reset,
  input logic [1:0][1:0] strm_ctrl_f2g,
  input logic [1:0][1:0] [15:0] strm_data_f2g,
  input logic [1:0][1:0] strm_data_f2g_vld,
  input logic [1:0][1:0] strm_data_g2f_rdy,
  input logic [1:0] strm_f2g_start_pulse,
  input logic [1:0] strm_g2f_start_pulse,
  output logic [1:0][1:0] [31:0] cgra_cfg_g2f_cfg_addr,
  output logic [1:0][1:0] [31:0] cgra_cfg_g2f_cfg_data,
  output logic [1:0][1:0] cgra_cfg_g2f_cfg_rd_en,
  output logic [1:0][1:0] cgra_cfg_g2f_cfg_wr_en,
  output logic [3:0] cgra_stall,
  output logic [31:0] if_cfg_rd_data,
  output logic if_cfg_rd_data_valid,
  output logic [31:0] if_sram_cfg_rd_data,
  output logic if_sram_cfg_rd_data_valid,
  output logic [1:0] pcfg_g2f_interrupt_pulse,
  output logic [63:0] proc_rd_data,
  output logic proc_rd_data_valid,
  output logic [1:0][1:0] strm_ctrl_g2f,
  output logic [1:0][1:0] strm_data_f2g_rdy,
  output logic strm_data_flush_g2f,
  output logic [1:0][1:0] [15:0] strm_data_g2f,
  output logic [1:0][1:0] strm_data_g2f_vld,
  output logic [1:0] strm_f2g_interrupt_pulse,
  output logic [1:0] strm_g2f_interrupt_pulse
);

typedef enum logic {
  axi = 1'h0,
  jtag = 1'h1
} proc_rd_type_e;
logic [2:0] cfg_pcfg_tile_connected;
logic [2:0] cfg_tile_connected;
logic [1:0][31:0] cgra_cfg_jtag_addr_bypass_esto;
logic [1:0][31:0] cgra_cfg_jtag_addr_bypass_wsti;
logic [1:0][31:0] cgra_cfg_jtag_addr_esto;
logic [1:0][31:0] cgra_cfg_jtag_addr_wsti;
logic [1:0][31:0] cgra_cfg_jtag_data_esto;
logic [1:0][31:0] cgra_cfg_jtag_data_wsti;
logic [31:0] cgra_cfg_jtag_gc2glb_addr_d;
logic [31:0] cgra_cfg_jtag_gc2glb_data_d;
logic cgra_cfg_jtag_gc2glb_rd_en_d;
logic cgra_cfg_jtag_gc2glb_wr_en_d;
logic [1:0] cgra_cfg_jtag_rd_en_bypass_esto;
logic [1:0] cgra_cfg_jtag_rd_en_bypass_wsti;
logic [1:0] cgra_cfg_jtag_rd_en_esto;
logic [1:0] cgra_cfg_jtag_rd_en_wsti;
logic [1:0] cgra_cfg_jtag_wr_en_esto;
logic [1:0] cgra_cfg_jtag_wr_en_wsti;
logic [1:0][31:0] cgra_cfg_pcfg_addr_esti;
logic [1:0][31:0] cgra_cfg_pcfg_addr_esto;
logic [1:0][31:0] cgra_cfg_pcfg_addr_wsti;
logic [1:0][31:0] cgra_cfg_pcfg_addr_wsto;
logic [1:0][31:0] cgra_cfg_pcfg_data_esti;
logic [1:0][31:0] cgra_cfg_pcfg_data_esto;
logic [1:0][31:0] cgra_cfg_pcfg_data_wsti;
logic [1:0][31:0] cgra_cfg_pcfg_data_wsto;
logic [1:0] cgra_cfg_pcfg_rd_en_esti;
logic [1:0] cgra_cfg_pcfg_rd_en_esto;
logic [1:0] cgra_cfg_pcfg_rd_en_wsti;
logic [1:0] cgra_cfg_pcfg_rd_en_wsto;
logic [1:0] cgra_cfg_pcfg_wr_en_esti;
logic [1:0] cgra_cfg_pcfg_wr_en_esto;
logic [1:0] cgra_cfg_pcfg_wr_en_wsti;
logic [1:0] cgra_cfg_pcfg_wr_en_wsto;
logic [1:0] data_flush;
logic [1:0] data_flush_d;
logic [1:0] flush_crossbar_in;
logic flush_crossbar_sel_w;
logic glb_tile_gen_0_cfg_pcfg_tile_connected_esto;
logic glb_tile_gen_0_cfg_tile_connected_esto;
logic [1:0][31:0] glb_tile_gen_0_cgra_cfg_g2f_cfg_addr;
logic [1:0][31:0] glb_tile_gen_0_cgra_cfg_g2f_cfg_data;
logic [1:0] glb_tile_gen_0_cgra_cfg_g2f_cfg_rd_en;
logic [1:0] glb_tile_gen_0_cgra_cfg_g2f_cfg_wr_en;
logic [31:0] glb_tile_gen_0_cgra_cfg_jtag_addr_bypass_esto;
logic [31:0] glb_tile_gen_0_cgra_cfg_jtag_addr_esto;
logic [31:0] glb_tile_gen_0_cgra_cfg_jtag_data_esto;
logic glb_tile_gen_0_cgra_cfg_jtag_rd_en_bypass_esto;
logic glb_tile_gen_0_cgra_cfg_jtag_rd_en_esto;
logic glb_tile_gen_0_cgra_cfg_jtag_wr_en_esto;
logic [31:0] glb_tile_gen_0_cgra_cfg_pcfg_addr_e2w_wsto;
logic [31:0] glb_tile_gen_0_cgra_cfg_pcfg_addr_w2e_esto;
logic [31:0] glb_tile_gen_0_cgra_cfg_pcfg_data_e2w_wsto;
logic [31:0] glb_tile_gen_0_cgra_cfg_pcfg_data_w2e_esto;
logic glb_tile_gen_0_cgra_cfg_pcfg_rd_en_e2w_wsto;
logic glb_tile_gen_0_cgra_cfg_pcfg_rd_en_w2e_esto;
logic glb_tile_gen_0_cgra_cfg_pcfg_wr_en_e2w_wsto;
logic glb_tile_gen_0_cgra_cfg_pcfg_wr_en_w2e_esto;
logic glb_tile_gen_0_clk_en_bank_master;
logic glb_tile_gen_0_clk_en_master;
logic glb_tile_gen_0_clk_en_pcfg_broadcast;
logic glb_tile_gen_0_data_flush;
logic glb_tile_gen_0_pcfg_g2f_interrupt_pulse;
logic [18:0] glb_tile_gen_0_pcfg_rd_addr_e2w_wsto;
logic [18:0] glb_tile_gen_0_pcfg_rd_addr_w2e_esto;
logic [63:0] glb_tile_gen_0_pcfg_rd_data_e2w_wsto;
logic glb_tile_gen_0_pcfg_rd_data_valid_e2w_wsto;
logic glb_tile_gen_0_pcfg_rd_data_valid_w2e_esto;
logic [63:0] glb_tile_gen_0_pcfg_rd_data_w2e_esto;
logic glb_tile_gen_0_pcfg_rd_en_e2w_wsto;
logic glb_tile_gen_0_pcfg_rd_en_w2e_esto;
logic [1:0] glb_tile_gen_0_strm_ctrl_g2f;
logic [1:0] glb_tile_gen_0_strm_data_f2g_rdy;
logic [1:0][15:0] glb_tile_gen_0_strm_data_g2f;
logic [1:0] glb_tile_gen_0_strm_data_g2f_vld;
logic glb_tile_gen_0_strm_f2g_interrupt_pulse;
logic glb_tile_gen_0_strm_g2f_interrupt_pulse;
logic [18:0] glb_tile_gen_0_strm_rd_addr_e2w_wsto;
logic [18:0] glb_tile_gen_0_strm_rd_addr_w2e_esto;
logic [63:0] glb_tile_gen_0_strm_rd_data_e2w_wsto;
logic glb_tile_gen_0_strm_rd_data_valid_e2w_wsto;
logic glb_tile_gen_0_strm_rd_data_valid_w2e_esto;
logic [63:0] glb_tile_gen_0_strm_rd_data_w2e_esto;
logic glb_tile_gen_0_strm_rd_en_e2w_wsto;
logic glb_tile_gen_0_strm_rd_en_w2e_esto;
logic [18:0] glb_tile_gen_0_strm_wr_addr_e2w_wsto;
logic [18:0] glb_tile_gen_0_strm_wr_addr_w2e_esto;
logic [63:0] glb_tile_gen_0_strm_wr_data_e2w_wsto;
logic [63:0] glb_tile_gen_0_strm_wr_data_w2e_esto;
logic glb_tile_gen_0_strm_wr_en_e2w_wsto;
logic glb_tile_gen_0_strm_wr_en_w2e_esto;
logic [7:0] glb_tile_gen_0_strm_wr_strb_e2w_wsto;
logic [7:0] glb_tile_gen_0_strm_wr_strb_w2e_esto;
logic glb_tile_gen_1_cfg_pcfg_tile_connected_esto;
logic glb_tile_gen_1_cfg_tile_connected_esto;
logic [1:0][31:0] glb_tile_gen_1_cgra_cfg_g2f_cfg_addr;
logic [1:0][31:0] glb_tile_gen_1_cgra_cfg_g2f_cfg_data;
logic [1:0] glb_tile_gen_1_cgra_cfg_g2f_cfg_rd_en;
logic [1:0] glb_tile_gen_1_cgra_cfg_g2f_cfg_wr_en;
logic [31:0] glb_tile_gen_1_cgra_cfg_jtag_addr_bypass_esto;
logic [31:0] glb_tile_gen_1_cgra_cfg_jtag_addr_esto;
logic [31:0] glb_tile_gen_1_cgra_cfg_jtag_data_esto;
logic glb_tile_gen_1_cgra_cfg_jtag_rd_en_bypass_esto;
logic glb_tile_gen_1_cgra_cfg_jtag_rd_en_esto;
logic glb_tile_gen_1_cgra_cfg_jtag_wr_en_esto;
logic [31:0] glb_tile_gen_1_cgra_cfg_pcfg_addr_e2w_wsto;
logic [31:0] glb_tile_gen_1_cgra_cfg_pcfg_addr_w2e_esto;
logic [31:0] glb_tile_gen_1_cgra_cfg_pcfg_data_e2w_wsto;
logic [31:0] glb_tile_gen_1_cgra_cfg_pcfg_data_w2e_esto;
logic glb_tile_gen_1_cgra_cfg_pcfg_rd_en_e2w_wsto;
logic glb_tile_gen_1_cgra_cfg_pcfg_rd_en_w2e_esto;
logic glb_tile_gen_1_cgra_cfg_pcfg_wr_en_e2w_wsto;
logic glb_tile_gen_1_cgra_cfg_pcfg_wr_en_w2e_esto;
logic glb_tile_gen_1_clk_en_bank_master;
logic glb_tile_gen_1_clk_en_master;
logic glb_tile_gen_1_clk_en_pcfg_broadcast;
logic glb_tile_gen_1_data_flush;
logic glb_tile_gen_1_pcfg_g2f_interrupt_pulse;
logic [18:0] glb_tile_gen_1_pcfg_rd_addr_e2w_wsto;
logic [18:0] glb_tile_gen_1_pcfg_rd_addr_w2e_esto;
logic [63:0] glb_tile_gen_1_pcfg_rd_data_e2w_wsto;
logic glb_tile_gen_1_pcfg_rd_data_valid_e2w_wsto;
logic glb_tile_gen_1_pcfg_rd_data_valid_w2e_esto;
logic [63:0] glb_tile_gen_1_pcfg_rd_data_w2e_esto;
logic glb_tile_gen_1_pcfg_rd_en_e2w_wsto;
logic glb_tile_gen_1_pcfg_rd_en_w2e_esto;
logic [1:0] glb_tile_gen_1_strm_ctrl_g2f;
logic [1:0] glb_tile_gen_1_strm_data_f2g_rdy;
logic [1:0][15:0] glb_tile_gen_1_strm_data_g2f;
logic [1:0] glb_tile_gen_1_strm_data_g2f_vld;
logic glb_tile_gen_1_strm_f2g_interrupt_pulse;
logic glb_tile_gen_1_strm_g2f_interrupt_pulse;
logic [18:0] glb_tile_gen_1_strm_rd_addr_e2w_wsto;
logic [18:0] glb_tile_gen_1_strm_rd_addr_w2e_esto;
logic [63:0] glb_tile_gen_1_strm_rd_data_e2w_wsto;
logic glb_tile_gen_1_strm_rd_data_valid_e2w_wsto;
logic glb_tile_gen_1_strm_rd_data_valid_w2e_esto;
logic [63:0] glb_tile_gen_1_strm_rd_data_w2e_esto;
logic glb_tile_gen_1_strm_rd_en_e2w_wsto;
logic glb_tile_gen_1_strm_rd_en_w2e_esto;
logic [18:0] glb_tile_gen_1_strm_wr_addr_e2w_wsto;
logic [18:0] glb_tile_gen_1_strm_wr_addr_w2e_esto;
logic [63:0] glb_tile_gen_1_strm_wr_data_e2w_wsto;
logic [63:0] glb_tile_gen_1_strm_wr_data_w2e_esto;
logic glb_tile_gen_1_strm_wr_en_e2w_wsto;
logic glb_tile_gen_1_strm_wr_en_w2e_esto;
logic [7:0] glb_tile_gen_1_strm_wr_strb_e2w_wsto;
logic [7:0] glb_tile_gen_1_strm_wr_strb_w2e_esto;
logic if_sram_cfg_rd_data_valid_w;
logic [31:0] if_sram_cfg_rd_data_w;
logic [1:0] pcfg_g2f_interrupt_pulse_d;
logic [1:0] pcfg_g2f_interrupt_pulse_w;
rd_packet_t [1:0] pcfg_packet_e2w_esti;
rd_packet_t [1:0] pcfg_packet_e2w_wsto;
rd_packet_t [1:0] pcfg_packet_w2e_esto;
rd_packet_t [1:0] pcfg_packet_w2e_wsti;
logic [18:0] proc_rd_addr_d;
logic proc_rd_addr_sel;
logic proc_rd_clk_en;
logic proc_rd_clk_en_gen_enable;
logic proc_rd_data_valid_w;
logic [63:0] proc_rd_data_w;
logic proc_rd_en_d;
proc_rd_type_e proc_rd_type;
logic [18:0] proc_wr_addr_d;
logic proc_wr_clk_en;
logic proc_wr_clk_en_gen_enable;
logic [63:0] proc_wr_data_d;
logic proc_wr_en_d;
logic [7:0] proc_wr_strb_d;
logic [18:0] sram_cfg_rd_addr_d;
logic sram_cfg_rd_en_d;
logic [18:0] sram_cfg_wr_addr_d;
logic [63:0] sram_cfg_wr_data_d;
logic sram_cfg_wr_en_d;
logic [7:0] sram_cfg_wr_strb_d;
logic [1:0] strm_f2g_interrupt_pulse_d;
logic [1:0] strm_f2g_interrupt_pulse_w;
logic [1:0] strm_g2f_interrupt_pulse_d;
logic [1:0] strm_g2f_interrupt_pulse_w;
packet_t [1:0] strm_packet_e2w_esti;
packet_t [1:0] strm_packet_e2w_wsto;
packet_t [1:0] strm_packet_w2e_esto;
packet_t [1:0] strm_packet_w2e_wsti;
glb_tile_ifc_A_12_D_32 if_cfg_tile2tile_0();
glb_tile_ifc_A_12_D_32 if_cfg_tile2tile_1();
glb_tile_ifc_A_12_D_32 if_cfg_tile2tile_2();
glb_tile_ifc_A_19_D_64 if_proc_tile2tile_0();
glb_tile_ifc_A_19_D_64 if_proc_tile2tile_1();
glb_tile_ifc_A_19_D_64 if_proc_tile2tile_2();
glb_tile_ifc_A_19_D_32 if_sram_cfg_tile2tile_0();
glb_tile_ifc_A_19_D_32 if_sram_cfg_tile2tile_1();
glb_tile_ifc_A_19_D_32 if_sram_cfg_tile2tile_2();
assign cfg_tile_connected[0] = 1'h0;
assign cfg_pcfg_tile_connected[0] = 1'h0;
assign strm_f2g_interrupt_pulse = strm_f2g_interrupt_pulse_d;
assign strm_g2f_interrupt_pulse = strm_g2f_interrupt_pulse_d;
assign pcfg_g2f_interrupt_pulse = pcfg_g2f_interrupt_pulse_d;
assign cgra_stall = cgra_stall_in;
assign if_sram_cfg_tile2tile_2.rd_data = 32'h0;
assign if_sram_cfg_tile2tile_2.rd_data_valid = 1'h0;
assign glb_tile_gen_0_clk_en_pcfg_broadcast = ~pcfg_broadcast_stall[0];
assign glb_tile_gen_0_clk_en_master = glb_clk_en_master[0];
assign glb_tile_gen_0_clk_en_bank_master = glb_clk_en_bank_master[0];
assign strm_packet_w2e_esto[0].wr.wr_en = glb_tile_gen_0_strm_wr_en_w2e_esto;
assign strm_packet_w2e_esto[0].wr.wr_strb = glb_tile_gen_0_strm_wr_strb_w2e_esto;
assign strm_packet_w2e_esto[0].wr.wr_addr = glb_tile_gen_0_strm_wr_addr_w2e_esto;
assign strm_packet_w2e_esto[0].wr.wr_data = glb_tile_gen_0_strm_wr_data_w2e_esto;
assign strm_packet_w2e_esto[0].rdrq.rd_en = glb_tile_gen_0_strm_rd_en_w2e_esto;
assign strm_packet_w2e_esto[0].rdrq.rd_addr = glb_tile_gen_0_strm_rd_addr_w2e_esto;
assign strm_packet_w2e_esto[0].rdrs.rd_data = glb_tile_gen_0_strm_rd_data_w2e_esto;
assign strm_packet_w2e_esto[0].rdrs.rd_data_valid = glb_tile_gen_0_strm_rd_data_valid_w2e_esto;
assign strm_packet_e2w_wsto[0].wr.wr_en = glb_tile_gen_0_strm_wr_en_e2w_wsto;
assign strm_packet_e2w_wsto[0].wr.wr_strb = glb_tile_gen_0_strm_wr_strb_e2w_wsto;
assign strm_packet_e2w_wsto[0].wr.wr_addr = glb_tile_gen_0_strm_wr_addr_e2w_wsto;
assign strm_packet_e2w_wsto[0].wr.wr_data = glb_tile_gen_0_strm_wr_data_e2w_wsto;
assign strm_packet_e2w_wsto[0].rdrq.rd_en = glb_tile_gen_0_strm_rd_en_e2w_wsto;
assign strm_packet_e2w_wsto[0].rdrq.rd_addr = glb_tile_gen_0_strm_rd_addr_e2w_wsto;
assign strm_packet_e2w_wsto[0].rdrs.rd_data = glb_tile_gen_0_strm_rd_data_e2w_wsto;
assign strm_packet_e2w_wsto[0].rdrs.rd_data_valid = glb_tile_gen_0_strm_rd_data_valid_e2w_wsto;
assign pcfg_packet_w2e_esto[0].rdrq.rd_en = glb_tile_gen_0_pcfg_rd_en_w2e_esto;
assign pcfg_packet_w2e_esto[0].rdrq.rd_addr = glb_tile_gen_0_pcfg_rd_addr_w2e_esto;
assign pcfg_packet_w2e_esto[0].rdrs.rd_data = glb_tile_gen_0_pcfg_rd_data_w2e_esto;
assign pcfg_packet_w2e_esto[0].rdrs.rd_data_valid = glb_tile_gen_0_pcfg_rd_data_valid_w2e_esto;
assign pcfg_packet_e2w_wsto[0].rdrq.rd_en = glb_tile_gen_0_pcfg_rd_en_e2w_wsto;
assign pcfg_packet_e2w_wsto[0].rdrq.rd_addr = glb_tile_gen_0_pcfg_rd_addr_e2w_wsto;
assign pcfg_packet_e2w_wsto[0].rdrs.rd_data = glb_tile_gen_0_pcfg_rd_data_e2w_wsto;
assign pcfg_packet_e2w_wsto[0].rdrs.rd_data_valid = glb_tile_gen_0_pcfg_rd_data_valid_e2w_wsto;
assign cfg_tile_connected[1] = glb_tile_gen_0_cfg_tile_connected_esto;
assign cfg_pcfg_tile_connected[1] = glb_tile_gen_0_cfg_pcfg_tile_connected_esto;
assign strm_data_f2g_rdy[0] = glb_tile_gen_0_strm_data_f2g_rdy;
assign strm_data_g2f[0] = glb_tile_gen_0_strm_data_g2f;
assign strm_data_g2f_vld[0] = glb_tile_gen_0_strm_data_g2f_vld;
assign strm_ctrl_g2f[0] = glb_tile_gen_0_strm_ctrl_g2f;
assign data_flush[0] = glb_tile_gen_0_data_flush;
assign cgra_cfg_g2f_cfg_wr_en[0] = glb_tile_gen_0_cgra_cfg_g2f_cfg_wr_en;
assign cgra_cfg_g2f_cfg_rd_en[0] = glb_tile_gen_0_cgra_cfg_g2f_cfg_rd_en;
assign cgra_cfg_g2f_cfg_addr[0] = glb_tile_gen_0_cgra_cfg_g2f_cfg_addr;
assign cgra_cfg_g2f_cfg_data[0] = glb_tile_gen_0_cgra_cfg_g2f_cfg_data;
assign cgra_cfg_pcfg_wr_en_esto[0] = glb_tile_gen_0_cgra_cfg_pcfg_wr_en_w2e_esto;
assign cgra_cfg_pcfg_rd_en_esto[0] = glb_tile_gen_0_cgra_cfg_pcfg_rd_en_w2e_esto;
assign cgra_cfg_pcfg_addr_esto[0] = glb_tile_gen_0_cgra_cfg_pcfg_addr_w2e_esto;
assign cgra_cfg_pcfg_data_esto[0] = glb_tile_gen_0_cgra_cfg_pcfg_data_w2e_esto;
assign cgra_cfg_pcfg_wr_en_wsto[0] = glb_tile_gen_0_cgra_cfg_pcfg_wr_en_e2w_wsto;
assign cgra_cfg_pcfg_rd_en_wsto[0] = glb_tile_gen_0_cgra_cfg_pcfg_rd_en_e2w_wsto;
assign cgra_cfg_pcfg_addr_wsto[0] = glb_tile_gen_0_cgra_cfg_pcfg_addr_e2w_wsto;
assign cgra_cfg_pcfg_data_wsto[0] = glb_tile_gen_0_cgra_cfg_pcfg_data_e2w_wsto;
assign cgra_cfg_jtag_wr_en_esto[0] = glb_tile_gen_0_cgra_cfg_jtag_wr_en_esto;
assign cgra_cfg_jtag_rd_en_esto[0] = glb_tile_gen_0_cgra_cfg_jtag_rd_en_esto;
assign cgra_cfg_jtag_addr_esto[0] = glb_tile_gen_0_cgra_cfg_jtag_addr_esto;
assign cgra_cfg_jtag_data_esto[0] = glb_tile_gen_0_cgra_cfg_jtag_data_esto;
assign cgra_cfg_jtag_rd_en_bypass_esto[0] = glb_tile_gen_0_cgra_cfg_jtag_rd_en_bypass_esto;
assign cgra_cfg_jtag_addr_bypass_esto[0] = glb_tile_gen_0_cgra_cfg_jtag_addr_bypass_esto;
assign strm_f2g_interrupt_pulse_w[0] = glb_tile_gen_0_strm_f2g_interrupt_pulse;
assign strm_g2f_interrupt_pulse_w[0] = glb_tile_gen_0_strm_g2f_interrupt_pulse;
assign pcfg_g2f_interrupt_pulse_w[0] = glb_tile_gen_0_pcfg_g2f_interrupt_pulse;
assign glb_tile_gen_1_clk_en_pcfg_broadcast = ~pcfg_broadcast_stall[1];
assign glb_tile_gen_1_clk_en_master = glb_clk_en_master[1];
assign glb_tile_gen_1_clk_en_bank_master = glb_clk_en_bank_master[1];
assign strm_packet_w2e_esto[1].wr.wr_en = glb_tile_gen_1_strm_wr_en_w2e_esto;
assign strm_packet_w2e_esto[1].wr.wr_strb = glb_tile_gen_1_strm_wr_strb_w2e_esto;
assign strm_packet_w2e_esto[1].wr.wr_addr = glb_tile_gen_1_strm_wr_addr_w2e_esto;
assign strm_packet_w2e_esto[1].wr.wr_data = glb_tile_gen_1_strm_wr_data_w2e_esto;
assign strm_packet_w2e_esto[1].rdrq.rd_en = glb_tile_gen_1_strm_rd_en_w2e_esto;
assign strm_packet_w2e_esto[1].rdrq.rd_addr = glb_tile_gen_1_strm_rd_addr_w2e_esto;
assign strm_packet_w2e_esto[1].rdrs.rd_data = glb_tile_gen_1_strm_rd_data_w2e_esto;
assign strm_packet_w2e_esto[1].rdrs.rd_data_valid = glb_tile_gen_1_strm_rd_data_valid_w2e_esto;
assign strm_packet_e2w_wsto[1].wr.wr_en = glb_tile_gen_1_strm_wr_en_e2w_wsto;
assign strm_packet_e2w_wsto[1].wr.wr_strb = glb_tile_gen_1_strm_wr_strb_e2w_wsto;
assign strm_packet_e2w_wsto[1].wr.wr_addr = glb_tile_gen_1_strm_wr_addr_e2w_wsto;
assign strm_packet_e2w_wsto[1].wr.wr_data = glb_tile_gen_1_strm_wr_data_e2w_wsto;
assign strm_packet_e2w_wsto[1].rdrq.rd_en = glb_tile_gen_1_strm_rd_en_e2w_wsto;
assign strm_packet_e2w_wsto[1].rdrq.rd_addr = glb_tile_gen_1_strm_rd_addr_e2w_wsto;
assign strm_packet_e2w_wsto[1].rdrs.rd_data = glb_tile_gen_1_strm_rd_data_e2w_wsto;
assign strm_packet_e2w_wsto[1].rdrs.rd_data_valid = glb_tile_gen_1_strm_rd_data_valid_e2w_wsto;
assign pcfg_packet_w2e_esto[1].rdrq.rd_en = glb_tile_gen_1_pcfg_rd_en_w2e_esto;
assign pcfg_packet_w2e_esto[1].rdrq.rd_addr = glb_tile_gen_1_pcfg_rd_addr_w2e_esto;
assign pcfg_packet_w2e_esto[1].rdrs.rd_data = glb_tile_gen_1_pcfg_rd_data_w2e_esto;
assign pcfg_packet_w2e_esto[1].rdrs.rd_data_valid = glb_tile_gen_1_pcfg_rd_data_valid_w2e_esto;
assign pcfg_packet_e2w_wsto[1].rdrq.rd_en = glb_tile_gen_1_pcfg_rd_en_e2w_wsto;
assign pcfg_packet_e2w_wsto[1].rdrq.rd_addr = glb_tile_gen_1_pcfg_rd_addr_e2w_wsto;
assign pcfg_packet_e2w_wsto[1].rdrs.rd_data = glb_tile_gen_1_pcfg_rd_data_e2w_wsto;
assign pcfg_packet_e2w_wsto[1].rdrs.rd_data_valid = glb_tile_gen_1_pcfg_rd_data_valid_e2w_wsto;
assign cfg_tile_connected[2] = glb_tile_gen_1_cfg_tile_connected_esto;
assign cfg_pcfg_tile_connected[2] = glb_tile_gen_1_cfg_pcfg_tile_connected_esto;
assign strm_data_f2g_rdy[1] = glb_tile_gen_1_strm_data_f2g_rdy;
assign strm_data_g2f[1] = glb_tile_gen_1_strm_data_g2f;
assign strm_data_g2f_vld[1] = glb_tile_gen_1_strm_data_g2f_vld;
assign strm_ctrl_g2f[1] = glb_tile_gen_1_strm_ctrl_g2f;
assign data_flush[1] = glb_tile_gen_1_data_flush;
assign cgra_cfg_g2f_cfg_wr_en[1] = glb_tile_gen_1_cgra_cfg_g2f_cfg_wr_en;
assign cgra_cfg_g2f_cfg_rd_en[1] = glb_tile_gen_1_cgra_cfg_g2f_cfg_rd_en;
assign cgra_cfg_g2f_cfg_addr[1] = glb_tile_gen_1_cgra_cfg_g2f_cfg_addr;
assign cgra_cfg_g2f_cfg_data[1] = glb_tile_gen_1_cgra_cfg_g2f_cfg_data;
assign cgra_cfg_pcfg_wr_en_esto[1] = glb_tile_gen_1_cgra_cfg_pcfg_wr_en_w2e_esto;
assign cgra_cfg_pcfg_rd_en_esto[1] = glb_tile_gen_1_cgra_cfg_pcfg_rd_en_w2e_esto;
assign cgra_cfg_pcfg_addr_esto[1] = glb_tile_gen_1_cgra_cfg_pcfg_addr_w2e_esto;
assign cgra_cfg_pcfg_data_esto[1] = glb_tile_gen_1_cgra_cfg_pcfg_data_w2e_esto;
assign cgra_cfg_pcfg_wr_en_wsto[1] = glb_tile_gen_1_cgra_cfg_pcfg_wr_en_e2w_wsto;
assign cgra_cfg_pcfg_rd_en_wsto[1] = glb_tile_gen_1_cgra_cfg_pcfg_rd_en_e2w_wsto;
assign cgra_cfg_pcfg_addr_wsto[1] = glb_tile_gen_1_cgra_cfg_pcfg_addr_e2w_wsto;
assign cgra_cfg_pcfg_data_wsto[1] = glb_tile_gen_1_cgra_cfg_pcfg_data_e2w_wsto;
assign cgra_cfg_jtag_wr_en_esto[1] = glb_tile_gen_1_cgra_cfg_jtag_wr_en_esto;
assign cgra_cfg_jtag_rd_en_esto[1] = glb_tile_gen_1_cgra_cfg_jtag_rd_en_esto;
assign cgra_cfg_jtag_addr_esto[1] = glb_tile_gen_1_cgra_cfg_jtag_addr_esto;
assign cgra_cfg_jtag_data_esto[1] = glb_tile_gen_1_cgra_cfg_jtag_data_esto;
assign cgra_cfg_jtag_rd_en_bypass_esto[1] = glb_tile_gen_1_cgra_cfg_jtag_rd_en_bypass_esto;
assign cgra_cfg_jtag_addr_bypass_esto[1] = glb_tile_gen_1_cgra_cfg_jtag_addr_bypass_esto;
assign strm_f2g_interrupt_pulse_w[1] = glb_tile_gen_1_strm_f2g_interrupt_pulse;
assign strm_g2f_interrupt_pulse_w[1] = glb_tile_gen_1_strm_g2f_interrupt_pulse;
assign pcfg_g2f_interrupt_pulse_w[1] = glb_tile_gen_1_pcfg_g2f_interrupt_pulse;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    proc_wr_en_d <= 1'h0;
    proc_wr_strb_d <= 8'h0;
    proc_wr_addr_d <= 19'h0;
    proc_wr_data_d <= 64'h0;
    proc_rd_en_d <= 1'h0;
    proc_rd_addr_d <= 19'h0;
  end
  else begin
    proc_wr_en_d <= proc_wr_en;
    proc_wr_strb_d <= proc_wr_strb;
    proc_wr_addr_d <= proc_wr_addr;
    proc_wr_data_d <= proc_wr_data;
    proc_rd_en_d <= proc_rd_en;
    proc_rd_addr_d <= proc_rd_addr;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    sram_cfg_wr_en_d <= 1'h0;
    sram_cfg_wr_strb_d <= 8'h0;
    sram_cfg_wr_addr_d <= 19'h0;
    sram_cfg_wr_data_d <= 64'h0;
    sram_cfg_rd_en_d <= 1'h0;
    sram_cfg_rd_addr_d <= 19'h0;
  end
  else begin
    sram_cfg_wr_en_d <= if_sram_cfg_wr_en;
    sram_cfg_wr_addr_d <= if_sram_cfg_wr_addr;
    if (if_sram_cfg_wr_addr[2] == 1'h0) begin
      sram_cfg_wr_data_d <= {32'h0, if_sram_cfg_wr_data};
      sram_cfg_wr_strb_d <= {4'h0, 4'hF};
    end
    else begin
      sram_cfg_wr_data_d <= {if_sram_cfg_wr_data[31:0], 32'h0};
      sram_cfg_wr_strb_d <= {4'hF, 4'h0};
    end
    sram_cfg_rd_en_d <= if_sram_cfg_rd_en;
    sram_cfg_rd_addr_d <= if_sram_cfg_rd_addr;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    if_proc_tile2tile_0.wr_en <= 1'h0;
    if_proc_tile2tile_0.wr_strb <= 8'h0;
    if_proc_tile2tile_0.wr_addr <= 19'h0;
    if_proc_tile2tile_0.wr_data <= 64'h0;
  end
  else if (proc_wr_en_d) begin
    if_proc_tile2tile_0.wr_en <= proc_wr_en_d;
    if_proc_tile2tile_0.wr_strb <= proc_wr_strb_d;
    if_proc_tile2tile_0.wr_addr <= proc_wr_addr_d;
    if_proc_tile2tile_0.wr_data <= proc_wr_data_d;
  end
  else if (sram_cfg_wr_en_d) begin
    if_proc_tile2tile_0.wr_en <= sram_cfg_wr_en_d;
    if_proc_tile2tile_0.wr_strb <= sram_cfg_wr_strb_d;
    if_proc_tile2tile_0.wr_addr <= sram_cfg_wr_addr_d;
    if_proc_tile2tile_0.wr_data <= sram_cfg_wr_data_d;
  end
  else begin
    if_proc_tile2tile_0.wr_en <= proc_wr_en_d;
    if_proc_tile2tile_0.wr_strb <= proc_wr_strb_d;
    if_proc_tile2tile_0.wr_addr <= proc_wr_addr_d;
    if_proc_tile2tile_0.wr_data <= proc_wr_data_d;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    if_proc_tile2tile_0.rd_en <= 1'h0;
    if_proc_tile2tile_0.rd_addr <= 19'h0;
    proc_rd_type <= axi;
    proc_rd_addr_sel <= 1'h0;
  end
  else if (proc_rd_en_d) begin
    if_proc_tile2tile_0.rd_en <= proc_rd_en_d;
    if_proc_tile2tile_0.rd_addr <= proc_rd_addr_d;
    proc_rd_type <= axi;
    proc_rd_addr_sel <= 1'h0;
  end
  else if (sram_cfg_rd_en_d) begin
    if_proc_tile2tile_0.rd_en <= sram_cfg_rd_en_d;
    if_proc_tile2tile_0.rd_addr <= sram_cfg_rd_addr_d;
    proc_rd_addr_sel <= sram_cfg_rd_addr_d[2];
    proc_rd_type <= jtag;
  end
  else begin
    if_proc_tile2tile_0.rd_en <= proc_rd_en_d;
    if_proc_tile2tile_0.rd_addr <= proc_rd_addr_d;
    proc_rd_type <= proc_rd_type;
    proc_rd_addr_sel <= proc_rd_addr_sel;
  end
end
always_comb begin
  if (proc_rd_type == axi) begin
    proc_rd_data_w = if_proc_tile2tile_0.rd_data;
    proc_rd_data_valid_w = if_proc_tile2tile_0.rd_data_valid;
    if_sram_cfg_rd_data_w = 32'h0;
    if_sram_cfg_rd_data_valid_w = 1'h0;
  end
  else if (proc_rd_type == jtag) begin
    proc_rd_data_w = 64'h0;
    proc_rd_data_valid_w = 1'h0;
    if (proc_rd_addr_sel == 1'h0) begin
      if_sram_cfg_rd_data_w = if_proc_tile2tile_0.rd_data[31:0];
    end
    else if_sram_cfg_rd_data_w = if_proc_tile2tile_0.rd_data[63:32];
    if_sram_cfg_rd_data_valid_w = if_proc_tile2tile_0.rd_data_valid;
  end
  else begin
    proc_rd_data_w = if_proc_tile2tile_0.rd_data;
    proc_rd_data_valid_w = if_proc_tile2tile_0.rd_data_valid;
    if_sram_cfg_rd_data_w = 32'h0;
    if_sram_cfg_rd_data_valid_w = 1'h0;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    proc_rd_data <= 64'h0;
    proc_rd_data_valid <= 1'h0;
    if_sram_cfg_rd_data <= 32'h0;
    if_sram_cfg_rd_data_valid <= 1'h0;
  end
  else begin
    proc_rd_data <= proc_rd_data_w;
    proc_rd_data_valid <= proc_rd_data_valid_w;
    if_sram_cfg_rd_data <= if_sram_cfg_rd_data_w;
    if_sram_cfg_rd_data_valid <= if_sram_cfg_rd_data_valid_w;
  end
end
assign proc_wr_clk_en_gen_enable = proc_wr_en_d | sram_cfg_wr_en_d;
assign if_proc_tile2tile_0.wr_clk_en = proc_wr_clk_en;
assign proc_rd_clk_en_gen_enable = proc_rd_en_d | sram_cfg_rd_en_d;
assign if_proc_tile2tile_0.rd_clk_en = proc_rd_clk_en;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    if_cfg_tile2tile_0.wr_en <= 1'h0;
    if_cfg_tile2tile_0.wr_clk_en <= 1'h0;
    if_cfg_tile2tile_0.wr_addr <= 12'h0;
    if_cfg_tile2tile_0.wr_data <= 32'h0;
    if_cfg_tile2tile_0.rd_en <= 1'h0;
    if_cfg_tile2tile_0.rd_clk_en <= 1'h0;
    if_cfg_tile2tile_0.rd_addr <= 12'h0;
  end
  else begin
    if_cfg_tile2tile_0.wr_en <= if_cfg_wr_en;
    if_cfg_tile2tile_0.wr_clk_en <= if_cfg_wr_clk_en;
    if_cfg_tile2tile_0.wr_addr <= if_cfg_wr_addr;
    if_cfg_tile2tile_0.wr_data <= if_cfg_wr_data;
    if_cfg_tile2tile_0.rd_en <= if_cfg_rd_en;
    if_cfg_tile2tile_0.rd_clk_en <= if_cfg_rd_clk_en;
    if_cfg_tile2tile_0.rd_addr <= if_cfg_rd_addr;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    cgra_cfg_jtag_gc2glb_wr_en_d <= 1'h0;
    cgra_cfg_jtag_gc2glb_rd_en_d <= 1'h0;
    cgra_cfg_jtag_gc2glb_addr_d <= 32'h0;
    cgra_cfg_jtag_gc2glb_data_d <= 32'h0;
  end
  else begin
    cgra_cfg_jtag_gc2glb_wr_en_d <= cgra_cfg_jtag_gc2glb_wr_en;
    cgra_cfg_jtag_gc2glb_rd_en_d <= cgra_cfg_jtag_gc2glb_rd_en;
    cgra_cfg_jtag_gc2glb_addr_d <= cgra_cfg_jtag_gc2glb_addr;
    cgra_cfg_jtag_gc2glb_data_d <= cgra_cfg_jtag_gc2glb_data;
  end
end
assign strm_packet_e2w_esti[1] = 177'h0;
assign pcfg_packet_e2w_esti[1] = 85'h0;
assign strm_packet_e2w_esti[0] = strm_packet_e2w_wsto[1];
assign pcfg_packet_e2w_esti[0] = pcfg_packet_e2w_wsto[1];
assign strm_packet_w2e_wsti[0] = 177'h0;
assign pcfg_packet_w2e_wsti[0] = 85'h0;
assign strm_packet_w2e_wsti[1] = strm_packet_w2e_esto[0];
assign pcfg_packet_w2e_wsti[1] = pcfg_packet_w2e_esto[0];
always_comb begin
  cgra_cfg_jtag_rd_en_wsti[0] = 1'h0;
  cgra_cfg_jtag_wr_en_wsti[0] = cgra_cfg_jtag_gc2glb_wr_en_d;
  cgra_cfg_jtag_addr_wsti[0] = cgra_cfg_jtag_gc2glb_addr_d;
  cgra_cfg_jtag_data_wsti[0] = cgra_cfg_jtag_gc2glb_data_d;
  cgra_cfg_jtag_rd_en_bypass_wsti[0] = cgra_cfg_jtag_gc2glb_rd_en_d;
  cgra_cfg_jtag_addr_bypass_wsti[0] = cgra_cfg_jtag_gc2glb_addr_d;
  cgra_cfg_pcfg_rd_en_wsti[0] = 1'h0;
  cgra_cfg_pcfg_wr_en_wsti[0] = 1'h0;
  cgra_cfg_pcfg_addr_wsti[0] = 32'h0;
  cgra_cfg_pcfg_data_wsti[0] = 32'h0;
  cgra_cfg_jtag_rd_en_wsti[1] = cgra_cfg_jtag_rd_en_esto[0];
  cgra_cfg_jtag_wr_en_wsti[1] = cgra_cfg_jtag_wr_en_esto[0];
  cgra_cfg_jtag_addr_wsti[1] = cgra_cfg_jtag_addr_esto[0];
  cgra_cfg_jtag_data_wsti[1] = cgra_cfg_jtag_data_esto[0];
  cgra_cfg_jtag_rd_en_bypass_wsti[1] = cgra_cfg_jtag_rd_en_bypass_esto[0];
  cgra_cfg_jtag_addr_bypass_wsti[1] = cgra_cfg_jtag_addr_bypass_esto[0];
  cgra_cfg_pcfg_rd_en_wsti[1] = cgra_cfg_pcfg_rd_en_esto[0];
  cgra_cfg_pcfg_wr_en_wsti[1] = cgra_cfg_pcfg_wr_en_esto[0];
  cgra_cfg_pcfg_addr_wsti[1] = cgra_cfg_pcfg_addr_esto[0];
  cgra_cfg_pcfg_data_wsti[1] = cgra_cfg_pcfg_data_esto[0];
end
always_comb begin
  cgra_cfg_pcfg_rd_en_esti[0] = cgra_cfg_pcfg_rd_en_wsto[1];
  cgra_cfg_pcfg_wr_en_esti[0] = cgra_cfg_pcfg_wr_en_wsto[1];
  cgra_cfg_pcfg_addr_esti[0] = cgra_cfg_pcfg_addr_wsto[1];
  cgra_cfg_pcfg_data_esti[0] = cgra_cfg_pcfg_data_wsto[1];
  cgra_cfg_pcfg_rd_en_esti[1] = 1'h0;
  cgra_cfg_pcfg_wr_en_esti[1] = 1'h0;
  cgra_cfg_pcfg_addr_esti[1] = 32'h0;
  cgra_cfg_pcfg_data_esti[1] = 32'h0;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    for (int unsigned i = 0; i < 2; i += 1) begin
        strm_f2g_interrupt_pulse_d[1'(i)] <= 1'h0;
        strm_g2f_interrupt_pulse_d[1'(i)] <= 1'h0;
        pcfg_g2f_interrupt_pulse_d[1'(i)] <= 1'h0;
      end
  end
  else begin
    for (int unsigned i = 0; i < 2; i += 1) begin
        strm_f2g_interrupt_pulse_d[1'(i)] <= strm_f2g_interrupt_pulse_w[1'(i)];
        strm_g2f_interrupt_pulse_d[1'(i)] <= strm_g2f_interrupt_pulse_w[1'(i)];
        pcfg_g2f_interrupt_pulse_d[1'(i)] <= pcfg_g2f_interrupt_pulse_w[1'(i)];
      end
  end
end
assign if_cfg_rd_data = if_cfg_tile2tile_0.rd_data;
assign if_cfg_rd_data_valid = if_cfg_tile2tile_0.rd_data_valid;
assign flush_crossbar_in[0] = data_flush_d[0];
assign flush_crossbar_in[1] = data_flush_d[1];
assign flush_crossbar_sel_w = flush_crossbar_sel;
glb_tile glb_tile_gen_0 (
  .cfg_pcfg_tile_connected_wsti(cfg_pcfg_tile_connected[0]),
  .cfg_tile_connected_wsti(cfg_tile_connected[0]),
  .cgra_cfg_jtag_addr_bypass_wsti(cgra_cfg_jtag_addr_bypass_wsti[0]),
  .cgra_cfg_jtag_addr_wsti(cgra_cfg_jtag_addr_wsti[0]),
  .cgra_cfg_jtag_data_wsti(cgra_cfg_jtag_data_wsti[0]),
  .cgra_cfg_jtag_rd_en_bypass_wsti(cgra_cfg_jtag_rd_en_bypass_wsti[0]),
  .cgra_cfg_jtag_rd_en_wsti(cgra_cfg_jtag_rd_en_wsti[0]),
  .cgra_cfg_jtag_wr_en_wsti(cgra_cfg_jtag_wr_en_wsti[0]),
  .cgra_cfg_pcfg_addr_e2w_esti(cgra_cfg_pcfg_addr_esti[0]),
  .cgra_cfg_pcfg_addr_w2e_wsti(cgra_cfg_pcfg_addr_wsti[0]),
  .cgra_cfg_pcfg_data_e2w_esti(cgra_cfg_pcfg_data_esti[0]),
  .cgra_cfg_pcfg_data_w2e_wsti(cgra_cfg_pcfg_data_wsti[0]),
  .cgra_cfg_pcfg_rd_en_e2w_esti(cgra_cfg_pcfg_rd_en_esti[0]),
  .cgra_cfg_pcfg_rd_en_w2e_wsti(cgra_cfg_pcfg_rd_en_wsti[0]),
  .cgra_cfg_pcfg_wr_en_e2w_esti(cgra_cfg_pcfg_wr_en_esti[0]),
  .cgra_cfg_pcfg_wr_en_w2e_wsti(cgra_cfg_pcfg_wr_en_wsti[0]),
  .clk(clk),
  .clk_en_bank_master(glb_tile_gen_0_clk_en_bank_master),
  .clk_en_master(glb_tile_gen_0_clk_en_master),
  .clk_en_pcfg_broadcast(glb_tile_gen_0_clk_en_pcfg_broadcast),
  .glb_tile_id(1'h0),
  .if_cfg_est_m_rd_data(if_cfg_tile2tile_1.rd_data),
  .if_cfg_est_m_rd_data_valid(if_cfg_tile2tile_1.rd_data_valid),
  .if_cfg_wst_s_rd_addr(if_cfg_tile2tile_0.rd_addr),
  .if_cfg_wst_s_rd_clk_en(if_cfg_tile2tile_0.rd_clk_en),
  .if_cfg_wst_s_rd_en(if_cfg_tile2tile_0.rd_en),
  .if_cfg_wst_s_wr_addr(if_cfg_tile2tile_0.wr_addr),
  .if_cfg_wst_s_wr_clk_en(if_cfg_tile2tile_0.wr_clk_en),
  .if_cfg_wst_s_wr_data(if_cfg_tile2tile_0.wr_data),
  .if_cfg_wst_s_wr_en(if_cfg_tile2tile_0.wr_en),
  .if_proc_est_m_rd_data(if_proc_tile2tile_1.rd_data),
  .if_proc_est_m_rd_data_valid(if_proc_tile2tile_1.rd_data_valid),
  .if_proc_wst_s_rd_addr(if_proc_tile2tile_0.rd_addr),
  .if_proc_wst_s_rd_clk_en(if_proc_tile2tile_0.rd_clk_en),
  .if_proc_wst_s_rd_en(if_proc_tile2tile_0.rd_en),
  .if_proc_wst_s_wr_addr(if_proc_tile2tile_0.wr_addr),
  .if_proc_wst_s_wr_clk_en(if_proc_tile2tile_0.wr_clk_en),
  .if_proc_wst_s_wr_data(if_proc_tile2tile_0.wr_data),
  .if_proc_wst_s_wr_en(if_proc_tile2tile_0.wr_en),
  .if_proc_wst_s_wr_strb(if_proc_tile2tile_0.wr_strb),
  .pcfg_rd_addr_e2w_esti(pcfg_packet_e2w_esti[0].rdrq.rd_addr),
  .pcfg_rd_addr_w2e_wsti(pcfg_packet_w2e_wsti[0].rdrq.rd_addr),
  .pcfg_rd_data_e2w_esti(pcfg_packet_e2w_esti[0].rdrs.rd_data),
  .pcfg_rd_data_valid_e2w_esti(pcfg_packet_e2w_esti[0].rdrs.rd_data_valid),
  .pcfg_rd_data_valid_w2e_wsti(pcfg_packet_w2e_wsti[0].rdrs.rd_data_valid),
  .pcfg_rd_data_w2e_wsti(pcfg_packet_w2e_wsti[0].rdrs.rd_data),
  .pcfg_rd_en_e2w_esti(pcfg_packet_e2w_esti[0].rdrq.rd_en),
  .pcfg_rd_en_w2e_wsti(pcfg_packet_w2e_wsti[0].rdrq.rd_en),
  .pcfg_start_pulse(pcfg_start_pulse[0]),
  .reset(reset),
  .strm_ctrl_f2g(strm_ctrl_f2g[0]),
  .strm_data_f2g(strm_data_f2g[0]),
  .strm_data_f2g_vld(strm_data_f2g_vld[0]),
  .strm_data_g2f_rdy(strm_data_g2f_rdy[0]),
  .strm_f2g_start_pulse(strm_f2g_start_pulse[0]),
  .strm_g2f_start_pulse(strm_g2f_start_pulse[0]),
  .strm_rd_addr_e2w_esti(strm_packet_e2w_esti[0].rdrq.rd_addr),
  .strm_rd_addr_w2e_wsti(strm_packet_w2e_wsti[0].rdrq.rd_addr),
  .strm_rd_data_e2w_esti(strm_packet_e2w_esti[0].rdrs.rd_data),
  .strm_rd_data_valid_e2w_esti(strm_packet_e2w_esti[0].rdrs.rd_data_valid),
  .strm_rd_data_valid_w2e_wsti(strm_packet_w2e_wsti[0].rdrs.rd_data_valid),
  .strm_rd_data_w2e_wsti(strm_packet_w2e_wsti[0].rdrs.rd_data),
  .strm_rd_en_e2w_esti(strm_packet_e2w_esti[0].rdrq.rd_en),
  .strm_rd_en_w2e_wsti(strm_packet_w2e_wsti[0].rdrq.rd_en),
  .strm_wr_addr_e2w_esti(strm_packet_e2w_esti[0].wr.wr_addr),
  .strm_wr_addr_w2e_wsti(strm_packet_w2e_wsti[0].wr.wr_addr),
  .strm_wr_data_e2w_esti(strm_packet_e2w_esti[0].wr.wr_data),
  .strm_wr_data_w2e_wsti(strm_packet_w2e_wsti[0].wr.wr_data),
  .strm_wr_en_e2w_esti(strm_packet_e2w_esti[0].wr.wr_en),
  .strm_wr_en_w2e_wsti(strm_packet_w2e_wsti[0].wr.wr_en),
  .strm_wr_strb_e2w_esti(strm_packet_e2w_esti[0].wr.wr_strb),
  .strm_wr_strb_w2e_wsti(strm_packet_w2e_wsti[0].wr.wr_strb),
  .cfg_pcfg_tile_connected_esto(glb_tile_gen_0_cfg_pcfg_tile_connected_esto),
  .cfg_tile_connected_esto(glb_tile_gen_0_cfg_tile_connected_esto),
  .cgra_cfg_g2f_cfg_addr(glb_tile_gen_0_cgra_cfg_g2f_cfg_addr),
  .cgra_cfg_g2f_cfg_data(glb_tile_gen_0_cgra_cfg_g2f_cfg_data),
  .cgra_cfg_g2f_cfg_rd_en(glb_tile_gen_0_cgra_cfg_g2f_cfg_rd_en),
  .cgra_cfg_g2f_cfg_wr_en(glb_tile_gen_0_cgra_cfg_g2f_cfg_wr_en),
  .cgra_cfg_jtag_addr_bypass_esto(glb_tile_gen_0_cgra_cfg_jtag_addr_bypass_esto),
  .cgra_cfg_jtag_addr_esto(glb_tile_gen_0_cgra_cfg_jtag_addr_esto),
  .cgra_cfg_jtag_data_esto(glb_tile_gen_0_cgra_cfg_jtag_data_esto),
  .cgra_cfg_jtag_rd_en_bypass_esto(glb_tile_gen_0_cgra_cfg_jtag_rd_en_bypass_esto),
  .cgra_cfg_jtag_rd_en_esto(glb_tile_gen_0_cgra_cfg_jtag_rd_en_esto),
  .cgra_cfg_jtag_wr_en_esto(glb_tile_gen_0_cgra_cfg_jtag_wr_en_esto),
  .cgra_cfg_pcfg_addr_e2w_wsto(glb_tile_gen_0_cgra_cfg_pcfg_addr_e2w_wsto),
  .cgra_cfg_pcfg_addr_w2e_esto(glb_tile_gen_0_cgra_cfg_pcfg_addr_w2e_esto),
  .cgra_cfg_pcfg_data_e2w_wsto(glb_tile_gen_0_cgra_cfg_pcfg_data_e2w_wsto),
  .cgra_cfg_pcfg_data_w2e_esto(glb_tile_gen_0_cgra_cfg_pcfg_data_w2e_esto),
  .cgra_cfg_pcfg_rd_en_e2w_wsto(glb_tile_gen_0_cgra_cfg_pcfg_rd_en_e2w_wsto),
  .cgra_cfg_pcfg_rd_en_w2e_esto(glb_tile_gen_0_cgra_cfg_pcfg_rd_en_w2e_esto),
  .cgra_cfg_pcfg_wr_en_e2w_wsto(glb_tile_gen_0_cgra_cfg_pcfg_wr_en_e2w_wsto),
  .cgra_cfg_pcfg_wr_en_w2e_esto(glb_tile_gen_0_cgra_cfg_pcfg_wr_en_w2e_esto),
  .data_flush(glb_tile_gen_0_data_flush),
  .if_cfg_est_m_rd_addr(if_cfg_tile2tile_1.rd_addr),
  .if_cfg_est_m_rd_clk_en(if_cfg_tile2tile_1.rd_clk_en),
  .if_cfg_est_m_rd_en(if_cfg_tile2tile_1.rd_en),
  .if_cfg_est_m_wr_addr(if_cfg_tile2tile_1.wr_addr),
  .if_cfg_est_m_wr_clk_en(if_cfg_tile2tile_1.wr_clk_en),
  .if_cfg_est_m_wr_data(if_cfg_tile2tile_1.wr_data),
  .if_cfg_est_m_wr_en(if_cfg_tile2tile_1.wr_en),
  .if_cfg_wst_s_rd_data(if_cfg_tile2tile_0.rd_data),
  .if_cfg_wst_s_rd_data_valid(if_cfg_tile2tile_0.rd_data_valid),
  .if_proc_est_m_rd_addr(if_proc_tile2tile_1.rd_addr),
  .if_proc_est_m_rd_clk_en(if_proc_tile2tile_1.rd_clk_en),
  .if_proc_est_m_rd_en(if_proc_tile2tile_1.rd_en),
  .if_proc_est_m_wr_addr(if_proc_tile2tile_1.wr_addr),
  .if_proc_est_m_wr_clk_en(if_proc_tile2tile_1.wr_clk_en),
  .if_proc_est_m_wr_data(if_proc_tile2tile_1.wr_data),
  .if_proc_est_m_wr_en(if_proc_tile2tile_1.wr_en),
  .if_proc_est_m_wr_strb(if_proc_tile2tile_1.wr_strb),
  .if_proc_wst_s_rd_data(if_proc_tile2tile_0.rd_data),
  .if_proc_wst_s_rd_data_valid(if_proc_tile2tile_0.rd_data_valid),
  .pcfg_g2f_interrupt_pulse(glb_tile_gen_0_pcfg_g2f_interrupt_pulse),
  .pcfg_rd_addr_e2w_wsto(glb_tile_gen_0_pcfg_rd_addr_e2w_wsto),
  .pcfg_rd_addr_w2e_esto(glb_tile_gen_0_pcfg_rd_addr_w2e_esto),
  .pcfg_rd_data_e2w_wsto(glb_tile_gen_0_pcfg_rd_data_e2w_wsto),
  .pcfg_rd_data_valid_e2w_wsto(glb_tile_gen_0_pcfg_rd_data_valid_e2w_wsto),
  .pcfg_rd_data_valid_w2e_esto(glb_tile_gen_0_pcfg_rd_data_valid_w2e_esto),
  .pcfg_rd_data_w2e_esto(glb_tile_gen_0_pcfg_rd_data_w2e_esto),
  .pcfg_rd_en_e2w_wsto(glb_tile_gen_0_pcfg_rd_en_e2w_wsto),
  .pcfg_rd_en_w2e_esto(glb_tile_gen_0_pcfg_rd_en_w2e_esto),
  .strm_ctrl_g2f(glb_tile_gen_0_strm_ctrl_g2f),
  .strm_data_f2g_rdy(glb_tile_gen_0_strm_data_f2g_rdy),
  .strm_data_g2f(glb_tile_gen_0_strm_data_g2f),
  .strm_data_g2f_vld(glb_tile_gen_0_strm_data_g2f_vld),
  .strm_f2g_interrupt_pulse(glb_tile_gen_0_strm_f2g_interrupt_pulse),
  .strm_g2f_interrupt_pulse(glb_tile_gen_0_strm_g2f_interrupt_pulse),
  .strm_rd_addr_e2w_wsto(glb_tile_gen_0_strm_rd_addr_e2w_wsto),
  .strm_rd_addr_w2e_esto(glb_tile_gen_0_strm_rd_addr_w2e_esto),
  .strm_rd_data_e2w_wsto(glb_tile_gen_0_strm_rd_data_e2w_wsto),
  .strm_rd_data_valid_e2w_wsto(glb_tile_gen_0_strm_rd_data_valid_e2w_wsto),
  .strm_rd_data_valid_w2e_esto(glb_tile_gen_0_strm_rd_data_valid_w2e_esto),
  .strm_rd_data_w2e_esto(glb_tile_gen_0_strm_rd_data_w2e_esto),
  .strm_rd_en_e2w_wsto(glb_tile_gen_0_strm_rd_en_e2w_wsto),
  .strm_rd_en_w2e_esto(glb_tile_gen_0_strm_rd_en_w2e_esto),
  .strm_wr_addr_e2w_wsto(glb_tile_gen_0_strm_wr_addr_e2w_wsto),
  .strm_wr_addr_w2e_esto(glb_tile_gen_0_strm_wr_addr_w2e_esto),
  .strm_wr_data_e2w_wsto(glb_tile_gen_0_strm_wr_data_e2w_wsto),
  .strm_wr_data_w2e_esto(glb_tile_gen_0_strm_wr_data_w2e_esto),
  .strm_wr_en_e2w_wsto(glb_tile_gen_0_strm_wr_en_e2w_wsto),
  .strm_wr_en_w2e_esto(glb_tile_gen_0_strm_wr_en_w2e_esto),
  .strm_wr_strb_e2w_wsto(glb_tile_gen_0_strm_wr_strb_e2w_wsto),
  .strm_wr_strb_w2e_esto(glb_tile_gen_0_strm_wr_strb_w2e_esto)
);

glb_tile glb_tile_gen_1 (
  .cfg_pcfg_tile_connected_wsti(cfg_pcfg_tile_connected[1]),
  .cfg_tile_connected_wsti(cfg_tile_connected[1]),
  .cgra_cfg_jtag_addr_bypass_wsti(cgra_cfg_jtag_addr_bypass_wsti[1]),
  .cgra_cfg_jtag_addr_wsti(cgra_cfg_jtag_addr_wsti[1]),
  .cgra_cfg_jtag_data_wsti(cgra_cfg_jtag_data_wsti[1]),
  .cgra_cfg_jtag_rd_en_bypass_wsti(cgra_cfg_jtag_rd_en_bypass_wsti[1]),
  .cgra_cfg_jtag_rd_en_wsti(cgra_cfg_jtag_rd_en_wsti[1]),
  .cgra_cfg_jtag_wr_en_wsti(cgra_cfg_jtag_wr_en_wsti[1]),
  .cgra_cfg_pcfg_addr_e2w_esti(cgra_cfg_pcfg_addr_esti[1]),
  .cgra_cfg_pcfg_addr_w2e_wsti(cgra_cfg_pcfg_addr_wsti[1]),
  .cgra_cfg_pcfg_data_e2w_esti(cgra_cfg_pcfg_data_esti[1]),
  .cgra_cfg_pcfg_data_w2e_wsti(cgra_cfg_pcfg_data_wsti[1]),
  .cgra_cfg_pcfg_rd_en_e2w_esti(cgra_cfg_pcfg_rd_en_esti[1]),
  .cgra_cfg_pcfg_rd_en_w2e_wsti(cgra_cfg_pcfg_rd_en_wsti[1]),
  .cgra_cfg_pcfg_wr_en_e2w_esti(cgra_cfg_pcfg_wr_en_esti[1]),
  .cgra_cfg_pcfg_wr_en_w2e_wsti(cgra_cfg_pcfg_wr_en_wsti[1]),
  .clk(clk),
  .clk_en_bank_master(glb_tile_gen_1_clk_en_bank_master),
  .clk_en_master(glb_tile_gen_1_clk_en_master),
  .clk_en_pcfg_broadcast(glb_tile_gen_1_clk_en_pcfg_broadcast),
  .glb_tile_id(1'h1),
  .if_cfg_est_m_rd_data(32'h0),
  .if_cfg_est_m_rd_data_valid(1'h0),
  .if_cfg_wst_s_rd_addr(if_cfg_tile2tile_1.rd_addr),
  .if_cfg_wst_s_rd_clk_en(if_cfg_tile2tile_1.rd_clk_en),
  .if_cfg_wst_s_rd_en(if_cfg_tile2tile_1.rd_en),
  .if_cfg_wst_s_wr_addr(if_cfg_tile2tile_1.wr_addr),
  .if_cfg_wst_s_wr_clk_en(if_cfg_tile2tile_1.wr_clk_en),
  .if_cfg_wst_s_wr_data(if_cfg_tile2tile_1.wr_data),
  .if_cfg_wst_s_wr_en(if_cfg_tile2tile_1.wr_en),
  .if_proc_est_m_rd_data(64'h0),
  .if_proc_est_m_rd_data_valid(1'h0),
  .if_proc_wst_s_rd_addr(if_proc_tile2tile_1.rd_addr),
  .if_proc_wst_s_rd_clk_en(if_proc_tile2tile_1.rd_clk_en),
  .if_proc_wst_s_rd_en(if_proc_tile2tile_1.rd_en),
  .if_proc_wst_s_wr_addr(if_proc_tile2tile_1.wr_addr),
  .if_proc_wst_s_wr_clk_en(if_proc_tile2tile_1.wr_clk_en),
  .if_proc_wst_s_wr_data(if_proc_tile2tile_1.wr_data),
  .if_proc_wst_s_wr_en(if_proc_tile2tile_1.wr_en),
  .if_proc_wst_s_wr_strb(if_proc_tile2tile_1.wr_strb),
  .pcfg_rd_addr_e2w_esti(pcfg_packet_e2w_esti[1].rdrq.rd_addr),
  .pcfg_rd_addr_w2e_wsti(pcfg_packet_w2e_wsti[1].rdrq.rd_addr),
  .pcfg_rd_data_e2w_esti(pcfg_packet_e2w_esti[1].rdrs.rd_data),
  .pcfg_rd_data_valid_e2w_esti(pcfg_packet_e2w_esti[1].rdrs.rd_data_valid),
  .pcfg_rd_data_valid_w2e_wsti(pcfg_packet_w2e_wsti[1].rdrs.rd_data_valid),
  .pcfg_rd_data_w2e_wsti(pcfg_packet_w2e_wsti[1].rdrs.rd_data),
  .pcfg_rd_en_e2w_esti(pcfg_packet_e2w_esti[1].rdrq.rd_en),
  .pcfg_rd_en_w2e_wsti(pcfg_packet_w2e_wsti[1].rdrq.rd_en),
  .pcfg_start_pulse(pcfg_start_pulse[1]),
  .reset(reset),
  .strm_ctrl_f2g(strm_ctrl_f2g[1]),
  .strm_data_f2g(strm_data_f2g[1]),
  .strm_data_f2g_vld(strm_data_f2g_vld[1]),
  .strm_data_g2f_rdy(strm_data_g2f_rdy[1]),
  .strm_f2g_start_pulse(strm_f2g_start_pulse[1]),
  .strm_g2f_start_pulse(strm_g2f_start_pulse[1]),
  .strm_rd_addr_e2w_esti(strm_packet_e2w_esti[1].rdrq.rd_addr),
  .strm_rd_addr_w2e_wsti(strm_packet_w2e_wsti[1].rdrq.rd_addr),
  .strm_rd_data_e2w_esti(strm_packet_e2w_esti[1].rdrs.rd_data),
  .strm_rd_data_valid_e2w_esti(strm_packet_e2w_esti[1].rdrs.rd_data_valid),
  .strm_rd_data_valid_w2e_wsti(strm_packet_w2e_wsti[1].rdrs.rd_data_valid),
  .strm_rd_data_w2e_wsti(strm_packet_w2e_wsti[1].rdrs.rd_data),
  .strm_rd_en_e2w_esti(strm_packet_e2w_esti[1].rdrq.rd_en),
  .strm_rd_en_w2e_wsti(strm_packet_w2e_wsti[1].rdrq.rd_en),
  .strm_wr_addr_e2w_esti(strm_packet_e2w_esti[1].wr.wr_addr),
  .strm_wr_addr_w2e_wsti(strm_packet_w2e_wsti[1].wr.wr_addr),
  .strm_wr_data_e2w_esti(strm_packet_e2w_esti[1].wr.wr_data),
  .strm_wr_data_w2e_wsti(strm_packet_w2e_wsti[1].wr.wr_data),
  .strm_wr_en_e2w_esti(strm_packet_e2w_esti[1].wr.wr_en),
  .strm_wr_en_w2e_wsti(strm_packet_w2e_wsti[1].wr.wr_en),
  .strm_wr_strb_e2w_esti(strm_packet_e2w_esti[1].wr.wr_strb),
  .strm_wr_strb_w2e_wsti(strm_packet_w2e_wsti[1].wr.wr_strb),
  .cfg_pcfg_tile_connected_esto(glb_tile_gen_1_cfg_pcfg_tile_connected_esto),
  .cfg_tile_connected_esto(glb_tile_gen_1_cfg_tile_connected_esto),
  .cgra_cfg_g2f_cfg_addr(glb_tile_gen_1_cgra_cfg_g2f_cfg_addr),
  .cgra_cfg_g2f_cfg_data(glb_tile_gen_1_cgra_cfg_g2f_cfg_data),
  .cgra_cfg_g2f_cfg_rd_en(glb_tile_gen_1_cgra_cfg_g2f_cfg_rd_en),
  .cgra_cfg_g2f_cfg_wr_en(glb_tile_gen_1_cgra_cfg_g2f_cfg_wr_en),
  .cgra_cfg_jtag_addr_bypass_esto(glb_tile_gen_1_cgra_cfg_jtag_addr_bypass_esto),
  .cgra_cfg_jtag_addr_esto(glb_tile_gen_1_cgra_cfg_jtag_addr_esto),
  .cgra_cfg_jtag_data_esto(glb_tile_gen_1_cgra_cfg_jtag_data_esto),
  .cgra_cfg_jtag_rd_en_bypass_esto(glb_tile_gen_1_cgra_cfg_jtag_rd_en_bypass_esto),
  .cgra_cfg_jtag_rd_en_esto(glb_tile_gen_1_cgra_cfg_jtag_rd_en_esto),
  .cgra_cfg_jtag_wr_en_esto(glb_tile_gen_1_cgra_cfg_jtag_wr_en_esto),
  .cgra_cfg_pcfg_addr_e2w_wsto(glb_tile_gen_1_cgra_cfg_pcfg_addr_e2w_wsto),
  .cgra_cfg_pcfg_addr_w2e_esto(glb_tile_gen_1_cgra_cfg_pcfg_addr_w2e_esto),
  .cgra_cfg_pcfg_data_e2w_wsto(glb_tile_gen_1_cgra_cfg_pcfg_data_e2w_wsto),
  .cgra_cfg_pcfg_data_w2e_esto(glb_tile_gen_1_cgra_cfg_pcfg_data_w2e_esto),
  .cgra_cfg_pcfg_rd_en_e2w_wsto(glb_tile_gen_1_cgra_cfg_pcfg_rd_en_e2w_wsto),
  .cgra_cfg_pcfg_rd_en_w2e_esto(glb_tile_gen_1_cgra_cfg_pcfg_rd_en_w2e_esto),
  .cgra_cfg_pcfg_wr_en_e2w_wsto(glb_tile_gen_1_cgra_cfg_pcfg_wr_en_e2w_wsto),
  .cgra_cfg_pcfg_wr_en_w2e_esto(glb_tile_gen_1_cgra_cfg_pcfg_wr_en_w2e_esto),
  .data_flush(glb_tile_gen_1_data_flush),
  .if_cfg_est_m_rd_addr(if_cfg_tile2tile_2.rd_addr),
  .if_cfg_est_m_rd_clk_en(if_cfg_tile2tile_2.rd_clk_en),
  .if_cfg_est_m_rd_en(if_cfg_tile2tile_2.rd_en),
  .if_cfg_est_m_wr_addr(if_cfg_tile2tile_2.wr_addr),
  .if_cfg_est_m_wr_clk_en(if_cfg_tile2tile_2.wr_clk_en),
  .if_cfg_est_m_wr_data(if_cfg_tile2tile_2.wr_data),
  .if_cfg_est_m_wr_en(if_cfg_tile2tile_2.wr_en),
  .if_cfg_wst_s_rd_data(if_cfg_tile2tile_1.rd_data),
  .if_cfg_wst_s_rd_data_valid(if_cfg_tile2tile_1.rd_data_valid),
  .if_proc_est_m_rd_addr(if_proc_tile2tile_2.rd_addr),
  .if_proc_est_m_rd_clk_en(if_proc_tile2tile_2.rd_clk_en),
  .if_proc_est_m_rd_en(if_proc_tile2tile_2.rd_en),
  .if_proc_est_m_wr_addr(if_proc_tile2tile_2.wr_addr),
  .if_proc_est_m_wr_clk_en(if_proc_tile2tile_2.wr_clk_en),
  .if_proc_est_m_wr_data(if_proc_tile2tile_2.wr_data),
  .if_proc_est_m_wr_en(if_proc_tile2tile_2.wr_en),
  .if_proc_est_m_wr_strb(if_proc_tile2tile_2.wr_strb),
  .if_proc_wst_s_rd_data(if_proc_tile2tile_1.rd_data),
  .if_proc_wst_s_rd_data_valid(if_proc_tile2tile_1.rd_data_valid),
  .pcfg_g2f_interrupt_pulse(glb_tile_gen_1_pcfg_g2f_interrupt_pulse),
  .pcfg_rd_addr_e2w_wsto(glb_tile_gen_1_pcfg_rd_addr_e2w_wsto),
  .pcfg_rd_addr_w2e_esto(glb_tile_gen_1_pcfg_rd_addr_w2e_esto),
  .pcfg_rd_data_e2w_wsto(glb_tile_gen_1_pcfg_rd_data_e2w_wsto),
  .pcfg_rd_data_valid_e2w_wsto(glb_tile_gen_1_pcfg_rd_data_valid_e2w_wsto),
  .pcfg_rd_data_valid_w2e_esto(glb_tile_gen_1_pcfg_rd_data_valid_w2e_esto),
  .pcfg_rd_data_w2e_esto(glb_tile_gen_1_pcfg_rd_data_w2e_esto),
  .pcfg_rd_en_e2w_wsto(glb_tile_gen_1_pcfg_rd_en_e2w_wsto),
  .pcfg_rd_en_w2e_esto(glb_tile_gen_1_pcfg_rd_en_w2e_esto),
  .strm_ctrl_g2f(glb_tile_gen_1_strm_ctrl_g2f),
  .strm_data_f2g_rdy(glb_tile_gen_1_strm_data_f2g_rdy),
  .strm_data_g2f(glb_tile_gen_1_strm_data_g2f),
  .strm_data_g2f_vld(glb_tile_gen_1_strm_data_g2f_vld),
  .strm_f2g_interrupt_pulse(glb_tile_gen_1_strm_f2g_interrupt_pulse),
  .strm_g2f_interrupt_pulse(glb_tile_gen_1_strm_g2f_interrupt_pulse),
  .strm_rd_addr_e2w_wsto(glb_tile_gen_1_strm_rd_addr_e2w_wsto),
  .strm_rd_addr_w2e_esto(glb_tile_gen_1_strm_rd_addr_w2e_esto),
  .strm_rd_data_e2w_wsto(glb_tile_gen_1_strm_rd_data_e2w_wsto),
  .strm_rd_data_valid_e2w_wsto(glb_tile_gen_1_strm_rd_data_valid_e2w_wsto),
  .strm_rd_data_valid_w2e_esto(glb_tile_gen_1_strm_rd_data_valid_w2e_esto),
  .strm_rd_data_w2e_esto(glb_tile_gen_1_strm_rd_data_w2e_esto),
  .strm_rd_en_e2w_wsto(glb_tile_gen_1_strm_rd_en_e2w_wsto),
  .strm_rd_en_w2e_esto(glb_tile_gen_1_strm_rd_en_w2e_esto),
  .strm_wr_addr_e2w_wsto(glb_tile_gen_1_strm_wr_addr_e2w_wsto),
  .strm_wr_addr_w2e_esto(glb_tile_gen_1_strm_wr_addr_w2e_esto),
  .strm_wr_data_e2w_wsto(glb_tile_gen_1_strm_wr_data_e2w_wsto),
  .strm_wr_data_w2e_esto(glb_tile_gen_1_strm_wr_data_w2e_esto),
  .strm_wr_en_e2w_wsto(glb_tile_gen_1_strm_wr_en_e2w_wsto),
  .strm_wr_en_w2e_esto(glb_tile_gen_1_strm_wr_en_w2e_esto),
  .strm_wr_strb_e2w_wsto(glb_tile_gen_1_strm_wr_strb_e2w_wsto),
  .strm_wr_strb_w2e_esto(glb_tile_gen_1_strm_wr_strb_w2e_esto)
);

glb_clk_en_gen_5 #(
  .cnt(32'h5))
proc_wr_clk_en_gen (
  .clk(clk),
  .enable(proc_wr_clk_en_gen_enable),
  .reset(reset),
  .clk_en(proc_wr_clk_en)
);

glb_clk_en_gen_11 #(
  .cnt(32'hB))
proc_rd_clk_en_gen (
  .clk(clk),
  .enable(proc_rd_clk_en_gen_enable),
  .reset(reset),
  .clk_en(proc_rd_clk_en)
);

pipeline_w_2_d_1 flush_pipeline (
  .clk(clk),
  .clk_en(1'h1),
  .in_(data_flush),
  .reset(reset),
  .out_(data_flush_d)
);

glb_crossbar_I_2_O_1_W_1 flush_crossbar (
  .in_(flush_crossbar_in),
  .sel_(flush_crossbar_sel_w),
  .out_(strm_data_flush_g2f)
);

endmodule   // global_buffer

module global_buffer_W (
  input logic [31:0] cgra_cfg_jtag_gc2glb_addr,
  input logic [31:0] cgra_cfg_jtag_gc2glb_data,
  input logic cgra_cfg_jtag_gc2glb_rd_en,
  input logic cgra_cfg_jtag_gc2glb_wr_en,
  input logic [3:0] cgra_stall_in,
  input logic clk,
  input logic flush_crossbar_sel,
  input logic [1:0] glb_clk_en_bank_master,
  input logic [1:0] glb_clk_en_master,
  input logic [11:0] if_cfg_rd_addr,
  input logic if_cfg_rd_clk_en,
  input logic if_cfg_rd_en,
  input logic [11:0] if_cfg_wr_addr,
  input logic if_cfg_wr_clk_en,
  input logic [31:0] if_cfg_wr_data,
  input logic if_cfg_wr_en,
  input logic [18:0] if_sram_cfg_rd_addr,
  input logic if_sram_cfg_rd_en,
  input logic [18:0] if_sram_cfg_wr_addr,
  input logic [31:0] if_sram_cfg_wr_data,
  input logic if_sram_cfg_wr_en,
  input logic [1:0] pcfg_broadcast_stall,
  input logic [1:0] pcfg_start_pulse,
  input logic [18:0] proc_rd_addr,
  input logic proc_rd_en,
  input logic [18:0] proc_wr_addr,
  input logic [63:0] proc_wr_data,
  input logic proc_wr_en,
  input logic [7:0] proc_wr_strb,
  input logic reset,
  input logic strm_ctrl_f2g_0_0,
  input logic strm_ctrl_f2g_0_1,
  input logic strm_ctrl_f2g_1_0,
  input logic strm_ctrl_f2g_1_1,
  input logic [15:0] strm_data_f2g_0_0,
  input logic [15:0] strm_data_f2g_0_1,
  input logic [15:0] strm_data_f2g_1_0,
  input logic [15:0] strm_data_f2g_1_1,
  input logic strm_data_f2g_vld_0_0,
  input logic strm_data_f2g_vld_0_1,
  input logic strm_data_f2g_vld_1_0,
  input logic strm_data_f2g_vld_1_1,
  input logic strm_data_g2f_rdy_0_0,
  input logic strm_data_g2f_rdy_0_1,
  input logic strm_data_g2f_rdy_1_0,
  input logic strm_data_g2f_rdy_1_1,
  input logic [1:0] strm_f2g_start_pulse,
  input logic [1:0] strm_g2f_start_pulse,
  output logic [31:0] cgra_cfg_g2f_cfg_addr_0_0,
  output logic [31:0] cgra_cfg_g2f_cfg_addr_0_1,
  output logic [31:0] cgra_cfg_g2f_cfg_addr_1_0,
  output logic [31:0] cgra_cfg_g2f_cfg_addr_1_1,
  output logic [31:0] cgra_cfg_g2f_cfg_data_0_0,
  output logic [31:0] cgra_cfg_g2f_cfg_data_0_1,
  output logic [31:0] cgra_cfg_g2f_cfg_data_1_0,
  output logic [31:0] cgra_cfg_g2f_cfg_data_1_1,
  output logic cgra_cfg_g2f_cfg_rd_en_0_0,
  output logic cgra_cfg_g2f_cfg_rd_en_0_1,
  output logic cgra_cfg_g2f_cfg_rd_en_1_0,
  output logic cgra_cfg_g2f_cfg_rd_en_1_1,
  output logic cgra_cfg_g2f_cfg_wr_en_0_0,
  output logic cgra_cfg_g2f_cfg_wr_en_0_1,
  output logic cgra_cfg_g2f_cfg_wr_en_1_0,
  output logic cgra_cfg_g2f_cfg_wr_en_1_1,
  output logic [3:0] cgra_stall,
  output logic [31:0] if_cfg_rd_data,
  output logic if_cfg_rd_data_valid,
  output logic [31:0] if_sram_cfg_rd_data,
  output logic if_sram_cfg_rd_data_valid,
  output logic [1:0] pcfg_g2f_interrupt_pulse,
  output logic [63:0] proc_rd_data,
  output logic proc_rd_data_valid,
  output logic strm_ctrl_g2f_0_0,
  output logic strm_ctrl_g2f_0_1,
  output logic strm_ctrl_g2f_1_0,
  output logic strm_ctrl_g2f_1_1,
  output logic strm_data_f2g_rdy_0_0,
  output logic strm_data_f2g_rdy_0_1,
  output logic strm_data_f2g_rdy_1_0,
  output logic strm_data_f2g_rdy_1_1,
  output logic strm_data_flush_g2f,
  output logic [15:0] strm_data_g2f_0_0,
  output logic [15:0] strm_data_g2f_0_1,
  output logic [15:0] strm_data_g2f_1_0,
  output logic [15:0] strm_data_g2f_1_1,
  output logic strm_data_g2f_vld_0_0,
  output logic strm_data_g2f_vld_0_1,
  output logic strm_data_g2f_vld_1_0,
  output logic strm_data_g2f_vld_1_1,
  output logic [1:0] strm_f2g_interrupt_pulse,
  output logic [1:0] strm_g2f_interrupt_pulse
);

logic [1:0][1:0][31:0] global_buffer_cgra_cfg_g2f_cfg_addr;
logic [1:0][1:0][31:0] global_buffer_cgra_cfg_g2f_cfg_data;
logic [1:0][1:0] global_buffer_cgra_cfg_g2f_cfg_rd_en;
logic [1:0][1:0] global_buffer_cgra_cfg_g2f_cfg_wr_en;
logic [1:0][1:0] global_buffer_strm_ctrl_f2g;
logic [1:0][1:0] global_buffer_strm_ctrl_g2f;
logic [1:0][1:0][15:0] global_buffer_strm_data_f2g;
logic [1:0][1:0] global_buffer_strm_data_f2g_rdy;
logic [1:0][1:0] global_buffer_strm_data_f2g_vld;
logic [1:0][1:0][15:0] global_buffer_strm_data_g2f;
logic [1:0][1:0] global_buffer_strm_data_g2f_rdy;
logic [1:0][1:0] global_buffer_strm_data_g2f_vld;
assign cgra_cfg_g2f_cfg_addr_0_0 = global_buffer_cgra_cfg_g2f_cfg_addr[0][0];
assign cgra_cfg_g2f_cfg_addr_0_1 = global_buffer_cgra_cfg_g2f_cfg_addr[0][1];
assign cgra_cfg_g2f_cfg_addr_1_0 = global_buffer_cgra_cfg_g2f_cfg_addr[1][0];
assign cgra_cfg_g2f_cfg_addr_1_1 = global_buffer_cgra_cfg_g2f_cfg_addr[1][1];
assign cgra_cfg_g2f_cfg_data_0_0 = global_buffer_cgra_cfg_g2f_cfg_data[0][0];
assign cgra_cfg_g2f_cfg_data_0_1 = global_buffer_cgra_cfg_g2f_cfg_data[0][1];
assign cgra_cfg_g2f_cfg_data_1_0 = global_buffer_cgra_cfg_g2f_cfg_data[1][0];
assign cgra_cfg_g2f_cfg_data_1_1 = global_buffer_cgra_cfg_g2f_cfg_data[1][1];
assign cgra_cfg_g2f_cfg_rd_en_0_0 = global_buffer_cgra_cfg_g2f_cfg_rd_en[0][0];
assign cgra_cfg_g2f_cfg_rd_en_0_1 = global_buffer_cgra_cfg_g2f_cfg_rd_en[0][1];
assign cgra_cfg_g2f_cfg_rd_en_1_0 = global_buffer_cgra_cfg_g2f_cfg_rd_en[1][0];
assign cgra_cfg_g2f_cfg_rd_en_1_1 = global_buffer_cgra_cfg_g2f_cfg_rd_en[1][1];
assign cgra_cfg_g2f_cfg_wr_en_0_0 = global_buffer_cgra_cfg_g2f_cfg_wr_en[0][0];
assign cgra_cfg_g2f_cfg_wr_en_0_1 = global_buffer_cgra_cfg_g2f_cfg_wr_en[0][1];
assign cgra_cfg_g2f_cfg_wr_en_1_0 = global_buffer_cgra_cfg_g2f_cfg_wr_en[1][0];
assign cgra_cfg_g2f_cfg_wr_en_1_1 = global_buffer_cgra_cfg_g2f_cfg_wr_en[1][1];
assign global_buffer_strm_ctrl_f2g[0][0] = strm_ctrl_f2g_0_0;
assign global_buffer_strm_ctrl_f2g[0][1] = strm_ctrl_f2g_0_1;
assign global_buffer_strm_ctrl_f2g[1][0] = strm_ctrl_f2g_1_0;
assign global_buffer_strm_ctrl_f2g[1][1] = strm_ctrl_f2g_1_1;
assign strm_ctrl_g2f_0_0 = global_buffer_strm_ctrl_g2f[0][0];
assign strm_ctrl_g2f_0_1 = global_buffer_strm_ctrl_g2f[0][1];
assign strm_ctrl_g2f_1_0 = global_buffer_strm_ctrl_g2f[1][0];
assign strm_ctrl_g2f_1_1 = global_buffer_strm_ctrl_g2f[1][1];
assign global_buffer_strm_data_f2g[0][0] = strm_data_f2g_0_0;
assign global_buffer_strm_data_f2g[0][1] = strm_data_f2g_0_1;
assign global_buffer_strm_data_f2g[1][0] = strm_data_f2g_1_0;
assign global_buffer_strm_data_f2g[1][1] = strm_data_f2g_1_1;
assign strm_data_f2g_rdy_0_0 = global_buffer_strm_data_f2g_rdy[0][0];
assign strm_data_f2g_rdy_0_1 = global_buffer_strm_data_f2g_rdy[0][1];
assign strm_data_f2g_rdy_1_0 = global_buffer_strm_data_f2g_rdy[1][0];
assign strm_data_f2g_rdy_1_1 = global_buffer_strm_data_f2g_rdy[1][1];
assign global_buffer_strm_data_f2g_vld[0][0] = strm_data_f2g_vld_0_0;
assign global_buffer_strm_data_f2g_vld[0][1] = strm_data_f2g_vld_0_1;
assign global_buffer_strm_data_f2g_vld[1][0] = strm_data_f2g_vld_1_0;
assign global_buffer_strm_data_f2g_vld[1][1] = strm_data_f2g_vld_1_1;
assign strm_data_g2f_0_0 = global_buffer_strm_data_g2f[0][0];
assign strm_data_g2f_0_1 = global_buffer_strm_data_g2f[0][1];
assign strm_data_g2f_1_0 = global_buffer_strm_data_g2f[1][0];
assign strm_data_g2f_1_1 = global_buffer_strm_data_g2f[1][1];
assign global_buffer_strm_data_g2f_rdy[0][0] = strm_data_g2f_rdy_0_0;
assign global_buffer_strm_data_g2f_rdy[0][1] = strm_data_g2f_rdy_0_1;
assign global_buffer_strm_data_g2f_rdy[1][0] = strm_data_g2f_rdy_1_0;
assign global_buffer_strm_data_g2f_rdy[1][1] = strm_data_g2f_rdy_1_1;
assign strm_data_g2f_vld_0_0 = global_buffer_strm_data_g2f_vld[0][0];
assign strm_data_g2f_vld_0_1 = global_buffer_strm_data_g2f_vld[0][1];
assign strm_data_g2f_vld_1_0 = global_buffer_strm_data_g2f_vld[1][0];
assign strm_data_g2f_vld_1_1 = global_buffer_strm_data_g2f_vld[1][1];
global_buffer global_buffer (
  .cgra_cfg_jtag_gc2glb_addr(cgra_cfg_jtag_gc2glb_addr),
  .cgra_cfg_jtag_gc2glb_data(cgra_cfg_jtag_gc2glb_data),
  .cgra_cfg_jtag_gc2glb_rd_en(cgra_cfg_jtag_gc2glb_rd_en),
  .cgra_cfg_jtag_gc2glb_wr_en(cgra_cfg_jtag_gc2glb_wr_en),
  .cgra_stall_in(cgra_stall_in),
  .clk(clk),
  .flush_crossbar_sel(flush_crossbar_sel),
  .glb_clk_en_bank_master(glb_clk_en_bank_master),
  .glb_clk_en_master(glb_clk_en_master),
  .if_cfg_rd_addr(if_cfg_rd_addr),
  .if_cfg_rd_clk_en(if_cfg_rd_clk_en),
  .if_cfg_rd_en(if_cfg_rd_en),
  .if_cfg_wr_addr(if_cfg_wr_addr),
  .if_cfg_wr_clk_en(if_cfg_wr_clk_en),
  .if_cfg_wr_data(if_cfg_wr_data),
  .if_cfg_wr_en(if_cfg_wr_en),
  .if_sram_cfg_rd_addr(if_sram_cfg_rd_addr),
  .if_sram_cfg_rd_en(if_sram_cfg_rd_en),
  .if_sram_cfg_wr_addr(if_sram_cfg_wr_addr),
  .if_sram_cfg_wr_data(if_sram_cfg_wr_data),
  .if_sram_cfg_wr_en(if_sram_cfg_wr_en),
  .pcfg_broadcast_stall(pcfg_broadcast_stall),
  .pcfg_start_pulse(pcfg_start_pulse),
  .proc_rd_addr(proc_rd_addr),
  .proc_rd_en(proc_rd_en),
  .proc_wr_addr(proc_wr_addr),
  .proc_wr_data(proc_wr_data),
  .proc_wr_en(proc_wr_en),
  .proc_wr_strb(proc_wr_strb),
  .reset(reset),
  .strm_ctrl_f2g(global_buffer_strm_ctrl_f2g),
  .strm_data_f2g(global_buffer_strm_data_f2g),
  .strm_data_f2g_vld(global_buffer_strm_data_f2g_vld),
  .strm_data_g2f_rdy(global_buffer_strm_data_g2f_rdy),
  .strm_f2g_start_pulse(strm_f2g_start_pulse),
  .strm_g2f_start_pulse(strm_g2f_start_pulse),
  .cgra_cfg_g2f_cfg_addr(global_buffer_cgra_cfg_g2f_cfg_addr),
  .cgra_cfg_g2f_cfg_data(global_buffer_cgra_cfg_g2f_cfg_data),
  .cgra_cfg_g2f_cfg_rd_en(global_buffer_cgra_cfg_g2f_cfg_rd_en),
  .cgra_cfg_g2f_cfg_wr_en(global_buffer_cgra_cfg_g2f_cfg_wr_en),
  .cgra_stall(cgra_stall),
  .if_cfg_rd_data(if_cfg_rd_data),
  .if_cfg_rd_data_valid(if_cfg_rd_data_valid),
  .if_sram_cfg_rd_data(if_sram_cfg_rd_data),
  .if_sram_cfg_rd_data_valid(if_sram_cfg_rd_data_valid),
  .pcfg_g2f_interrupt_pulse(pcfg_g2f_interrupt_pulse),
  .proc_rd_data(proc_rd_data),
  .proc_rd_data_valid(proc_rd_data_valid),
  .strm_ctrl_g2f(global_buffer_strm_ctrl_g2f),
  .strm_data_f2g_rdy(global_buffer_strm_data_f2g_rdy),
  .strm_data_flush_g2f(strm_data_flush_g2f),
  .strm_data_g2f(global_buffer_strm_data_g2f),
  .strm_data_g2f_vld(global_buffer_strm_data_g2f_vld),
  .strm_f2g_interrupt_pulse(strm_f2g_interrupt_pulse),
  .strm_g2f_interrupt_pulse(strm_g2f_interrupt_pulse)
);

endmodule   // global_buffer_W

module pipeline_w_144_d_0 (
  input logic clk,
  input logic clk_en,
  input logic [143:0] in_,
  input logic reset,
  output logic [143:0] out_
);

assign out_ = in_;
endmodule   // pipeline_w_144_d_0

module pipeline_w_18_d_0 (
  input logic clk,
  input logic clk_en,
  input logic [17:0] in_,
  input logic reset,
  output logic [17:0] out_
);

assign out_ = in_;
endmodule   // pipeline_w_18_d_0

module pipeline_w_1_d_0 (
  input logic clk,
  input logic clk_en,
  input logic in_,
  input logic reset,
  output logic out_
);

assign out_ = in_;
endmodule   // pipeline_w_1_d_0

module pipeline_w_1_d_1 (
  input logic clk,
  input logic clk_en,
  input logic in_,
  input logic reset,
  output logic out_
);

logic pipeline_r;
assign out_ = pipeline_r;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    pipeline_r <= 1'h0;
  end
  else if (clk_en) begin
    pipeline_r <= in_;
  end
end
endmodule   // pipeline_w_1_d_1

module pipeline_w_1_d_12_array (
  input logic clk,
  input logic clk_en,
  input logic in_,
  input logic reset,
  output logic out_ [11:0]
);

logic pipeline_r [11:0];
assign out_ = pipeline_r;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    pipeline_r[0] <= 1'h0;
    pipeline_r[1] <= 1'h0;
    pipeline_r[2] <= 1'h0;
    pipeline_r[3] <= 1'h0;
    pipeline_r[4] <= 1'h0;
    pipeline_r[5] <= 1'h0;
    pipeline_r[6] <= 1'h0;
    pipeline_r[7] <= 1'h0;
    pipeline_r[8] <= 1'h0;
    pipeline_r[9] <= 1'h0;
    pipeline_r[10] <= 1'h0;
    pipeline_r[11] <= 1'h0;
  end
  else if (clk_en) begin
    pipeline_r[0] <= in_;
    pipeline_r[1] <= pipeline_r[4'h0];
    pipeline_r[2] <= pipeline_r[4'h1];
    pipeline_r[3] <= pipeline_r[4'h2];
    pipeline_r[4] <= pipeline_r[4'h3];
    pipeline_r[5] <= pipeline_r[4'h4];
    pipeline_r[6] <= pipeline_r[4'h5];
    pipeline_r[7] <= pipeline_r[4'h6];
    pipeline_r[8] <= pipeline_r[4'h7];
    pipeline_r[9] <= pipeline_r[4'h8];
    pipeline_r[10] <= pipeline_r[4'h9];
    pipeline_r[11] <= pipeline_r[4'hA];
  end
end
endmodule   // pipeline_w_1_d_12_array

module pipeline_w_1_d_20_array (
  input logic clk,
  input logic clk_en,
  input logic in_,
  input logic reset,
  output logic out_ [19:0]
);

logic pipeline_r [19:0];
assign out_ = pipeline_r;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    pipeline_r[0] <= 1'h0;
    pipeline_r[1] <= 1'h0;
    pipeline_r[2] <= 1'h0;
    pipeline_r[3] <= 1'h0;
    pipeline_r[4] <= 1'h0;
    pipeline_r[5] <= 1'h0;
    pipeline_r[6] <= 1'h0;
    pipeline_r[7] <= 1'h0;
    pipeline_r[8] <= 1'h0;
    pipeline_r[9] <= 1'h0;
    pipeline_r[10] <= 1'h0;
    pipeline_r[11] <= 1'h0;
    pipeline_r[12] <= 1'h0;
    pipeline_r[13] <= 1'h0;
    pipeline_r[14] <= 1'h0;
    pipeline_r[15] <= 1'h0;
    pipeline_r[16] <= 1'h0;
    pipeline_r[17] <= 1'h0;
    pipeline_r[18] <= 1'h0;
    pipeline_r[19] <= 1'h0;
  end
  else if (clk_en) begin
    pipeline_r[0] <= in_;
    pipeline_r[1] <= pipeline_r[5'h0];
    pipeline_r[2] <= pipeline_r[5'h1];
    pipeline_r[3] <= pipeline_r[5'h2];
    pipeline_r[4] <= pipeline_r[5'h3];
    pipeline_r[5] <= pipeline_r[5'h4];
    pipeline_r[6] <= pipeline_r[5'h5];
    pipeline_r[7] <= pipeline_r[5'h6];
    pipeline_r[8] <= pipeline_r[5'h7];
    pipeline_r[9] <= pipeline_r[5'h8];
    pipeline_r[10] <= pipeline_r[5'h9];
    pipeline_r[11] <= pipeline_r[5'hA];
    pipeline_r[12] <= pipeline_r[5'hB];
    pipeline_r[13] <= pipeline_r[5'hC];
    pipeline_r[14] <= pipeline_r[5'hD];
    pipeline_r[15] <= pipeline_r[5'hE];
    pipeline_r[16] <= pipeline_r[5'hF];
    pipeline_r[17] <= pipeline_r[5'h10];
    pipeline_r[18] <= pipeline_r[5'h11];
    pipeline_r[19] <= pipeline_r[5'h12];
  end
end
endmodule   // pipeline_w_1_d_20_array

module pipeline_w_1_d_22_array (
  input logic clk,
  input logic clk_en,
  input logic in_,
  input logic reset,
  output logic out_ [21:0]
);

logic pipeline_r [21:0];
assign out_ = pipeline_r;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    pipeline_r[0] <= 1'h0;
    pipeline_r[1] <= 1'h0;
    pipeline_r[2] <= 1'h0;
    pipeline_r[3] <= 1'h0;
    pipeline_r[4] <= 1'h0;
    pipeline_r[5] <= 1'h0;
    pipeline_r[6] <= 1'h0;
    pipeline_r[7] <= 1'h0;
    pipeline_r[8] <= 1'h0;
    pipeline_r[9] <= 1'h0;
    pipeline_r[10] <= 1'h0;
    pipeline_r[11] <= 1'h0;
    pipeline_r[12] <= 1'h0;
    pipeline_r[13] <= 1'h0;
    pipeline_r[14] <= 1'h0;
    pipeline_r[15] <= 1'h0;
    pipeline_r[16] <= 1'h0;
    pipeline_r[17] <= 1'h0;
    pipeline_r[18] <= 1'h0;
    pipeline_r[19] <= 1'h0;
    pipeline_r[20] <= 1'h0;
    pipeline_r[21] <= 1'h0;
  end
  else if (clk_en) begin
    pipeline_r[0] <= in_;
    pipeline_r[1] <= pipeline_r[5'h0];
    pipeline_r[2] <= pipeline_r[5'h1];
    pipeline_r[3] <= pipeline_r[5'h2];
    pipeline_r[4] <= pipeline_r[5'h3];
    pipeline_r[5] <= pipeline_r[5'h4];
    pipeline_r[6] <= pipeline_r[5'h5];
    pipeline_r[7] <= pipeline_r[5'h6];
    pipeline_r[8] <= pipeline_r[5'h7];
    pipeline_r[9] <= pipeline_r[5'h8];
    pipeline_r[10] <= pipeline_r[5'h9];
    pipeline_r[11] <= pipeline_r[5'hA];
    pipeline_r[12] <= pipeline_r[5'hB];
    pipeline_r[13] <= pipeline_r[5'hC];
    pipeline_r[14] <= pipeline_r[5'hD];
    pipeline_r[15] <= pipeline_r[5'hE];
    pipeline_r[16] <= pipeline_r[5'hF];
    pipeline_r[17] <= pipeline_r[5'h10];
    pipeline_r[18] <= pipeline_r[5'h11];
    pipeline_r[19] <= pipeline_r[5'h12];
    pipeline_r[20] <= pipeline_r[5'h13];
    pipeline_r[21] <= pipeline_r[5'h14];
  end
end
endmodule   // pipeline_w_1_d_22_array

module pipeline_w_1_d_24_array (
  input logic clk,
  input logic clk_en,
  input logic in_,
  input logic reset,
  output logic out_ [23:0]
);

logic pipeline_r [23:0];
assign out_ = pipeline_r;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    pipeline_r[0] <= 1'h0;
    pipeline_r[1] <= 1'h0;
    pipeline_r[2] <= 1'h0;
    pipeline_r[3] <= 1'h0;
    pipeline_r[4] <= 1'h0;
    pipeline_r[5] <= 1'h0;
    pipeline_r[6] <= 1'h0;
    pipeline_r[7] <= 1'h0;
    pipeline_r[8] <= 1'h0;
    pipeline_r[9] <= 1'h0;
    pipeline_r[10] <= 1'h0;
    pipeline_r[11] <= 1'h0;
    pipeline_r[12] <= 1'h0;
    pipeline_r[13] <= 1'h0;
    pipeline_r[14] <= 1'h0;
    pipeline_r[15] <= 1'h0;
    pipeline_r[16] <= 1'h0;
    pipeline_r[17] <= 1'h0;
    pipeline_r[18] <= 1'h0;
    pipeline_r[19] <= 1'h0;
    pipeline_r[20] <= 1'h0;
    pipeline_r[21] <= 1'h0;
    pipeline_r[22] <= 1'h0;
    pipeline_r[23] <= 1'h0;
  end
  else if (clk_en) begin
    pipeline_r[0] <= in_;
    pipeline_r[1] <= pipeline_r[5'h0];
    pipeline_r[2] <= pipeline_r[5'h1];
    pipeline_r[3] <= pipeline_r[5'h2];
    pipeline_r[4] <= pipeline_r[5'h3];
    pipeline_r[5] <= pipeline_r[5'h4];
    pipeline_r[6] <= pipeline_r[5'h5];
    pipeline_r[7] <= pipeline_r[5'h6];
    pipeline_r[8] <= pipeline_r[5'h7];
    pipeline_r[9] <= pipeline_r[5'h8];
    pipeline_r[10] <= pipeline_r[5'h9];
    pipeline_r[11] <= pipeline_r[5'hA];
    pipeline_r[12] <= pipeline_r[5'hB];
    pipeline_r[13] <= pipeline_r[5'hC];
    pipeline_r[14] <= pipeline_r[5'hD];
    pipeline_r[15] <= pipeline_r[5'hE];
    pipeline_r[16] <= pipeline_r[5'hF];
    pipeline_r[17] <= pipeline_r[5'h10];
    pipeline_r[18] <= pipeline_r[5'h11];
    pipeline_r[19] <= pipeline_r[5'h12];
    pipeline_r[20] <= pipeline_r[5'h13];
    pipeline_r[21] <= pipeline_r[5'h14];
    pipeline_r[22] <= pipeline_r[5'h15];
    pipeline_r[23] <= pipeline_r[5'h16];
  end
end
endmodule   // pipeline_w_1_d_24_array

module pipeline_w_1_d_5 (
  input logic clk,
  input logic clk_en,
  input logic in_,
  input logic reset,
  output logic out_
);

logic pipeline_r [4:0];
assign out_ = pipeline_r[4];

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    pipeline_r[0] <= 1'h0;
    pipeline_r[1] <= 1'h0;
    pipeline_r[2] <= 1'h0;
    pipeline_r[3] <= 1'h0;
    pipeline_r[4] <= 1'h0;
  end
  else if (clk_en) begin
    pipeline_r[0] <= in_;
    pipeline_r[1] <= pipeline_r[3'h0];
    pipeline_r[2] <= pipeline_r[3'h1];
    pipeline_r[3] <= pipeline_r[3'h2];
    pipeline_r[4] <= pipeline_r[3'h3];
  end
end
endmodule   // pipeline_w_1_d_5

module pipeline_w_2_d_1 (
  input logic clk,
  input logic clk_en,
  input logic [1:0] in_,
  input logic reset,
  output logic [1:0] out_
);

logic [1:0] pipeline_r [0:0];
assign out_ = pipeline_r[0];

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    for (int unsigned i = 0; i < 1; i += 1) begin
        pipeline_r[1'(i)] <= 2'h0;
      end
  end
  else if (clk_en) begin
    for (int unsigned i = 0; i < 1; i += 1) begin
        if (i == 32'h0) begin
          pipeline_r[1'(i)] <= in_;
        end
        else pipeline_r[1'(i)] <= pipeline_r[1'(i - 32'h1)];
      end
  end
end
endmodule   // pipeline_w_2_d_1

module pipeline_w_2_d_2 (
  input logic clk,
  input logic clk_en,
  input logic [1:0] in_,
  input logic reset,
  output logic [1:0] out_
);

logic [1:0] pipeline_r [1:0];
assign out_ = pipeline_r[1];

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    for (int unsigned i = 0; i < 2; i += 1) begin
        pipeline_r[1'(i)] <= 2'h0;
      end
  end
  else if (clk_en) begin
    for (int unsigned i = 0; i < 2; i += 1) begin
        if (i == 32'h0) begin
          pipeline_r[1'(i)] <= in_;
        end
        else pipeline_r[1'(i)] <= pipeline_r[1'(i - 32'h1)];
      end
  end
end
endmodule   // pipeline_w_2_d_2

module pipeline_w_2_d_22_array (
  input logic clk,
  input logic clk_en,
  input logic [1:0] in_,
  input logic reset,
  output logic [1:0] out_ [21:0]
);

logic [1:0] pipeline_r [21:0];
assign out_ = pipeline_r;

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    for (int unsigned i = 0; i < 22; i += 1) begin
        pipeline_r[5'(i)] <= 2'h0;
      end
  end
  else if (clk_en) begin
    for (int unsigned i = 0; i < 22; i += 1) begin
        if (i == 32'h0) begin
          pipeline_r[5'(i)] <= in_;
        end
        else pipeline_r[5'(i)] <= pipeline_r[5'(i - 32'h1)];
      end
  end
end
endmodule   // pipeline_w_2_d_22_array

module pipeline_w_4_d_2 (
  input logic clk,
  input logic clk_en,
  input logic [3:0] in_,
  input logic reset,
  output logic [3:0] out_
);

logic [3:0] pipeline_r [1:0];
assign out_ = pipeline_r[1];

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    for (int unsigned i = 0; i < 2; i += 1) begin
        pipeline_r[1'(i)] <= 4'h0;
      end
  end
  else if (clk_en) begin
    for (int unsigned i = 0; i < 2; i += 1) begin
        if (i == 32'h0) begin
          pipeline_r[1'(i)] <= in_;
        end
        else pipeline_r[1'(i)] <= pipeline_r[1'(i - 32'h1)];
      end
  end
end
endmodule   // pipeline_w_4_d_2

module pipeline_w_64_d_0 (
  input logic clk,
  input logic clk_en,
  input logic [63:0] in_,
  input logic reset,
  output logic [63:0] out_
);

assign out_ = in_;
endmodule   // pipeline_w_64_d_0

module pipeline_w_65_d_1 (
  input logic clk,
  input logic clk_en,
  input logic [64:0] in_,
  input logic reset,
  output logic [64:0] out_
);

logic [64:0] pipeline_r [0:0];
assign out_ = pipeline_r[0];

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    for (int unsigned i = 0; i < 1; i += 1) begin
        pipeline_r[1'(i)] <= 65'h0;
      end
  end
  else if (clk_en) begin
    for (int unsigned i = 0; i < 1; i += 1) begin
        if (i == 32'h0) begin
          pipeline_r[1'(i)] <= in_;
        end
        else pipeline_r[1'(i)] <= pipeline_r[1'(i - 32'h1)];
      end
  end
end
endmodule   // pipeline_w_65_d_1

module pipeline_w_74_d_0_reset_high (
  input logic clk,
  input logic clk_en,
  input logic [73:0] in_,
  input logic reset,
  output logic [73:0] out_
);

assign out_ = in_;
endmodule   // pipeline_w_74_d_0_reset_high

module pipeline_w_78_d_0 (
  input logic clk,
  input logic clk_en,
  input logic [77:0] in_,
  input logic reset,
  output logic [77:0] out_
);

assign out_ = in_;
endmodule   // pipeline_w_78_d_0

module pipeline_w_90_d_0 (
  input logic clk,
  input logic clk_en,
  input logic [89:0] in_,
  input logic reset,
  output logic [89:0] out_
);

assign out_ = in_;
endmodule   // pipeline_w_90_d_0

module reg_fifo_d_19_w_16 #(
  parameter data_width = 16'h10
)
(
  input logic [4:0] almost_empty_diff,
  input logic [4:0] almost_full_diff,
  input logic clk,
  input logic clk_en,
  input logic [data_width-1:0] data_in,
  input logic flush,
  input logic pop,
  input logic push,
  input logic reset,
  output logic almost_empty,
  output logic almost_full,
  output logic [data_width-1:0] data_out,
  output logic empty,
  output logic full
);

logic [5:0] num_items;
logic [4:0] rd_ptr;
logic read;
logic [18:0][data_width-1:0] reg_array;
logic [4:0] wr_ptr;
logic write;
assign full = num_items == 6'h13;
assign empty = num_items == 6'h0;
assign read = pop & (~empty);
assign write = push & (~full);
always_comb begin
  almost_full = (6'h13 - 6'(almost_full_diff)) <= num_items;
  almost_empty = 6'(almost_empty_diff) >= num_items;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    num_items <= 6'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      num_items <= 6'h0;
    end
    else if (write & (~read)) begin
      num_items <= num_items + 6'h1;
    end
    else if ((~write) & read) begin
      num_items <= num_items - 6'h1;
    end
    else num_items <= num_items;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    reg_array <= 304'h0;
  end
  else if (clk_en) begin
    if (write) begin
      reg_array[wr_ptr] <= data_in;
    end
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    wr_ptr <= 5'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      wr_ptr <= 5'h0;
    end
    else if (write) begin
      if (wr_ptr == 5'h12) begin
        wr_ptr <= 5'h0;
      end
      else wr_ptr <= wr_ptr + 5'h1;
    end
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    rd_ptr <= 5'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      rd_ptr <= 5'h0;
    end
    else if (read) begin
      if (rd_ptr == 5'h12) begin
        rd_ptr <= 5'h0;
      end
      else rd_ptr <= rd_ptr + 5'h1;
    end
  end
end
always_comb begin
  data_out = reg_array[rd_ptr];
end
endmodule   // reg_fifo_d_19_w_16

module reg_fifo_d_2_w_16 #(
  parameter data_width = 16'h10
)
(
  input logic almost_empty_diff,
  input logic almost_full_diff,
  input logic clk,
  input logic clk_en,
  input logic [data_width-1:0] data_in,
  input logic flush,
  input logic pop,
  input logic push,
  input logic reset,
  output logic almost_empty,
  output logic almost_full,
  output logic [data_width-1:0] data_out,
  output logic empty,
  output logic full
);

logic [1:0] num_items;
logic rd_ptr;
logic read;
logic [1:0][data_width-1:0] reg_array;
logic wr_ptr;
logic write;
assign full = num_items == 2'h2;
assign empty = num_items == 2'h0;
assign read = pop & (~empty);
assign write = push & (~full);
always_comb begin
  almost_full = (2'h2 - 2'(almost_full_diff)) <= num_items;
  almost_empty = 2'(almost_empty_diff) >= num_items;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    num_items <= 2'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      num_items <= 2'h0;
    end
    else if (write & (~read)) begin
      num_items <= num_items + 2'h1;
    end
    else if ((~write) & read) begin
      num_items <= num_items - 2'h1;
    end
    else num_items <= num_items;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    reg_array <= 32'h0;
  end
  else if (clk_en) begin
    if (write) begin
      reg_array[wr_ptr] <= data_in;
    end
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    wr_ptr <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      wr_ptr <= 1'h0;
    end
    else if (write) begin
      if (wr_ptr == 1'h1) begin
        wr_ptr <= 1'h0;
      end
      else wr_ptr <= wr_ptr + 1'h1;
    end
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    rd_ptr <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      rd_ptr <= 1'h0;
    end
    else if (read) begin
      if (rd_ptr == 1'h1) begin
        rd_ptr <= 1'h0;
      end
      else rd_ptr <= rd_ptr + 1'h1;
    end
  end
end
always_comb begin
  data_out = reg_array[rd_ptr];
end
endmodule   // reg_fifo_d_2_w_16

module reg_fifo_d_4_w_16 #(
  parameter data_width = 16'h10
)
(
  input logic [1:0] almost_empty_diff,
  input logic [1:0] almost_full_diff,
  input logic clk,
  input logic clk_en,
  input logic [data_width-1:0] data_in,
  input logic flush,
  input logic pop,
  input logic push,
  input logic reset,
  output logic almost_empty,
  output logic almost_full,
  output logic [data_width-1:0] data_out,
  output logic empty,
  output logic full
);

logic [2:0] num_items;
logic [1:0] rd_ptr;
logic read;
logic [3:0][data_width-1:0] reg_array;
logic [1:0] wr_ptr;
logic write;
assign full = num_items == 3'h4;
assign empty = num_items == 3'h0;
assign read = pop & (~empty);
assign write = push & (~full);
always_comb begin
  almost_full = (3'h4 - 3'(almost_full_diff)) <= num_items;
  almost_empty = 3'(almost_empty_diff) >= num_items;
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    num_items <= 3'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      num_items <= 3'h0;
    end
    else if (write & (~read)) begin
      num_items <= num_items + 3'h1;
    end
    else if ((~write) & read) begin
      num_items <= num_items - 3'h1;
    end
    else num_items <= num_items;
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    reg_array <= 64'h0;
  end
  else if (clk_en) begin
    if (write) begin
      reg_array[wr_ptr] <= data_in;
    end
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    wr_ptr <= 2'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      wr_ptr <= 2'h0;
    end
    else if (write) begin
      if (wr_ptr == 2'h3) begin
        wr_ptr <= 2'h0;
      end
      else wr_ptr <= wr_ptr + 2'h1;
    end
  end
end

always_ff @(posedge clk, posedge reset) begin
  if (reset) begin
    rd_ptr <= 2'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      rd_ptr <= 2'h0;
    end
    else if (read) begin
      if (rd_ptr == 2'h3) begin
        rd_ptr <= 2'h0;
      end
      else rd_ptr <= rd_ptr + 2'h1;
    end
  end
end
always_comb begin
  data_out = reg_array[rd_ptr];
end
endmodule   // reg_fifo_d_4_w_16


module coreir_wrap (
    input in,
    output out
);
  assign out = in;
endmodule

module coreir_ult #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = in0 < in1;
endmodule

module coreir_reg #(
    parameter width = 1,
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input [width-1:0] in,
    output [width-1:0] out
);
  reg [width-1:0] outReg=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module coreir_orr #(
    parameter width = 1
) (
    input [width-1:0] in,
    output out
);
  assign out = |in;
endmodule

module coreir_or #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 | in1;
endmodule

module coreir_not #(
    parameter width = 1
) (
    input [width-1:0] in,
    output [width-1:0] out
);
  assign out = ~in;
endmodule

module coreir_mux #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    input sel,
    output [width-1:0] out
);
  assign out = sel ? in1 : in0;
endmodule

module coreir_eq #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = in0 == in1;
endmodule

module coreir_const #(
    parameter width = 1,
    parameter value = 1
) (
    output [width-1:0] out
);
  assign out = value;
endmodule

module coreir_andr #(
    parameter width = 1
) (
    input [width-1:0] in,
    output out
);
  assign out = &in;
endmodule

module coreir_and #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 & in1;
endmodule

module corebit_const #(
    parameter value = 1
) (
    output out
);
  assign out = value;
endmodule

module corebit_and (
    input in0,
    input in1,
    output out
);
  assign out = in0 & in1;
endmodule

module and_cell(input A, input B, output Z);
AN_CELL inst(.A1(A), .A2(B), .Z(Z));
endmodule
module SplitFifo_17 (
  input logic clk,
  input logic clk_en,
  input logic [16:0] data_in,
  input logic end_fifo,
  input logic fifo_en,
  input logic ready1,
  input logic rst,
  input logic start_fifo,
  input logic valid0,
  output logic [16:0] data_out,
  output logic ready0,
  output logic valid1
);

logic empty;
logic empty_n;
logic ready_in;
logic valid_in;
logic [16:0] value;
assign empty = ~empty_n;
assign ready_in = ready1 && (~start_fifo);
assign ready0 = fifo_en ? empty || ready_in: clk_en;
assign valid_in = valid0 && (~end_fifo);
assign valid1 = fifo_en ? (~empty) || valid_in: clk_en;
assign data_out = (empty && fifo_en) ? data_in: value;

always_ff @(posedge clk, posedge rst) begin
  if (rst) begin
    value <= 17'h0;
  end
  else if (clk_en) begin
    if ((~fifo_en) || (valid0 && ready0 && (~(empty && ready1 && valid1)))) begin
      value <= data_in;
    end
  end
end

always_ff @(posedge clk, posedge rst) begin
  if (rst) begin
    empty_n <= 1'h0;
  end
  else if (clk_en) begin
    if (fifo_en) begin
      if (valid1 && ready1) begin
        if (~(valid0 && ready0)) begin
          empty_n <= 1'h0;
        end
      end
      else if (valid0 && ready0) begin
        empty_n <= 1'h1;
      end
    end
  end
end
endmodule   // SplitFifo_17


module SplitFifo_1 (
  input logic clk,
  input logic clk_en,
  input logic data_in,
  input logic end_fifo,
  input logic fifo_en,
  input logic ready1,
  input logic rst,
  input logic start_fifo,
  input logic valid0,
  output logic data_out,
  output logic ready0,
  output logic valid1
);

logic empty;
logic empty_n;
logic ready_in;
logic valid_in;
logic value;
assign empty = ~empty_n;
assign ready_in = ready1 && (~start_fifo);
assign ready0 = fifo_en ? empty || ready_in: clk_en;
assign valid_in = valid0 && (~end_fifo);
assign valid1 = fifo_en ? (~empty) || valid_in: clk_en;
assign data_out = (empty && fifo_en) ? data_in: value;

always_ff @(posedge clk, posedge rst) begin
  if (rst) begin
    value <= 1'h0;
  end
  else if (clk_en) begin
    if ((~fifo_en) || (valid0 && ready0 && (~(empty && ready1 && valid1)))) begin
      value <= data_in;
    end
  end
end

always_ff @(posedge clk, posedge rst) begin
  if (rst) begin
    empty_n <= 1'h0;
  end
  else if (clk_en) begin
    if (fifo_en) begin
      if (valid1 && ready1) begin
        if (~(valid0 && ready0)) begin
          empty_n <= 1'h0;
        end
      end
      else if (valid0 && ready0) begin
        empty_n <= 1'h1;
      end
    end
  end
end
endmodule   // SplitFifo_1


module SliceWrapper_6_1_6 (
    input [5:0] I,
    output [4:0] O
);
assign O = I[5:1];
endmodule

module SliceWrapper_6_0_1 (
    input [5:0] I,
    output [0:0] O
);
assign O = I[0:0];
endmodule

module SliceWrapper_32_9_10 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[9:9];
endmodule

module SliceWrapper_32_8_9 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[8:8];
endmodule

module SliceWrapper_32_7_8 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[7:7];
endmodule

module SliceWrapper_32_6_7 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[6:6];
endmodule

module SliceWrapper_32_5_6 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[5:5];
endmodule

module SliceWrapper_32_4_5 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[4:4];
endmodule

module SliceWrapper_32_3_4 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[3:3];
endmodule

module SliceWrapper_32_31_32 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[31:31];
endmodule

module SliceWrapper_32_30_31 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[30:30];
endmodule

module SliceWrapper_32_2_3 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[2:2];
endmodule

module SliceWrapper_32_29_30 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[29:29];
endmodule

module SliceWrapper_32_28_31 (
    input [31:0] I,
    output [2:0] O
);
assign O = I[30:28];
endmodule

module SliceWrapper_32_28_29 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[28:28];
endmodule

module SliceWrapper_32_27_28 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[27:27];
endmodule

module SliceWrapper_32_26_27 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[26:26];
endmodule

module SliceWrapper_32_25_26 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[25:25];
endmodule

module SliceWrapper_32_24_25 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[24:24];
endmodule

module SliceWrapper_32_23_26 (
    input [31:0] I,
    output [2:0] O
);
assign O = I[25:23];
endmodule

module SliceWrapper_32_23_24 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[23:23];
endmodule

module SliceWrapper_32_22_23 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[22:22];
endmodule

module SliceWrapper_32_21_22 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[21:21];
endmodule

module SliceWrapper_32_20_21 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[20:20];
endmodule

module SliceWrapper_32_1_2 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[1:1];
endmodule

module SliceWrapper_32_19_20 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[19:19];
endmodule

module SliceWrapper_32_18_21 (
    input [31:0] I,
    output [2:0] O
);
assign O = I[20:18];
endmodule

module SliceWrapper_32_18_19 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[18:18];
endmodule

module SliceWrapper_32_17_18 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[17:17];
endmodule

module SliceWrapper_32_16_17 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[16:16];
endmodule

module SliceWrapper_32_15_16 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[15:15];
endmodule

module SliceWrapper_32_14_15 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[14:14];
endmodule

module SliceWrapper_32_13_14 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[13:13];
endmodule

module SliceWrapper_32_12_13 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[12:12];
endmodule

module SliceWrapper_32_11_12 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[11:11];
endmodule

module SliceWrapper_32_10_11 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[10:10];
endmodule

module SliceWrapper_32_0_32 (
    input [31:0] I,
    output [31:0] O
);
assign O = I;
endmodule

module SliceWrapper_32_0_22 (
    input [31:0] I,
    output [21:0] O
);
assign O = I[21:0];
endmodule

module SliceWrapper_32_0_1 (
    input [31:0] I,
    output [0:0] O
);
assign O = I[0:0];
endmodule

module SliceWrapper_31_9_10 (
    input [30:0] I,
    output [0:0] O
);
assign O = I[9:9];
endmodule

module SliceWrapper_31_6_9 (
    input [30:0] I,
    output [2:0] O
);
assign O = I[8:6];
endmodule

module SliceWrapper_31_5_6 (
    input [30:0] I,
    output [0:0] O
);
assign O = I[5:5];
endmodule

module SliceWrapper_31_4_5 (
    input [30:0] I,
    output [0:0] O
);
assign O = I[4:4];
endmodule

module SliceWrapper_31_30_31 (
    input [30:0] I,
    output [0:0] O
);
assign O = I[30:30];
endmodule

module SliceWrapper_31_29_30 (
    input [30:0] I,
    output [0:0] O
);
assign O = I[29:29];
endmodule

module SliceWrapper_31_26_29 (
    input [30:0] I,
    output [2:0] O
);
assign O = I[28:26];
endmodule

module SliceWrapper_31_25_26 (
    input [30:0] I,
    output [0:0] O
);
assign O = I[25:25];
endmodule

module SliceWrapper_31_24_25 (
    input [30:0] I,
    output [0:0] O
);
assign O = I[24:24];
endmodule

module SliceWrapper_31_21_24 (
    input [30:0] I,
    output [2:0] O
);
assign O = I[23:21];
endmodule

module SliceWrapper_31_20_21 (
    input [30:0] I,
    output [0:0] O
);
assign O = I[20:20];
endmodule

module SliceWrapper_31_1_4 (
    input [30:0] I,
    output [2:0] O
);
assign O = I[3:1];
endmodule

module SliceWrapper_31_19_20 (
    input [30:0] I,
    output [0:0] O
);
assign O = I[19:19];
endmodule

module SliceWrapper_31_16_19 (
    input [30:0] I,
    output [2:0] O
);
assign O = I[18:16];
endmodule

module SliceWrapper_31_15_16 (
    input [30:0] I,
    output [0:0] O
);
assign O = I[15:15];
endmodule

module SliceWrapper_31_14_15 (
    input [30:0] I,
    output [0:0] O
);
assign O = I[14:14];
endmodule

module SliceWrapper_31_11_14 (
    input [30:0] I,
    output [2:0] O
);
assign O = I[13:11];
endmodule

module SliceWrapper_31_10_11 (
    input [30:0] I,
    output [0:0] O
);
assign O = I[10:10];
endmodule

module SliceWrapper_31_0_1 (
    input [30:0] I,
    output [0:0] O
);
assign O = I[0:0];
endmodule

module SliceWrapper_30_9_10 (
    input [29:0] I,
    output [0:0] O
);
assign O = I[9:9];
endmodule

module SliceWrapper_30_8_9 (
    input [29:0] I,
    output [0:0] O
);
assign O = I[8:8];
endmodule

module SliceWrapper_30_5_8 (
    input [29:0] I,
    output [2:0] O
);
assign O = I[7:5];
endmodule

module SliceWrapper_30_4_5 (
    input [29:0] I,
    output [0:0] O
);
assign O = I[4:4];
endmodule

module SliceWrapper_30_3_4 (
    input [29:0] I,
    output [0:0] O
);
assign O = I[3:3];
endmodule

module SliceWrapper_30_29_30 (
    input [29:0] I,
    output [0:0] O
);
assign O = I[29:29];
endmodule

module SliceWrapper_30_28_29 (
    input [29:0] I,
    output [0:0] O
);
assign O = I[28:28];
endmodule

module SliceWrapper_30_25_28 (
    input [29:0] I,
    output [2:0] O
);
assign O = I[27:25];
endmodule

module SliceWrapper_30_24_25 (
    input [29:0] I,
    output [0:0] O
);
assign O = I[24:24];
endmodule

module SliceWrapper_30_23_24 (
    input [29:0] I,
    output [0:0] O
);
assign O = I[23:23];
endmodule

module SliceWrapper_30_20_23 (
    input [29:0] I,
    output [2:0] O
);
assign O = I[22:20];
endmodule

module SliceWrapper_30_19_20 (
    input [29:0] I,
    output [0:0] O
);
assign O = I[19:19];
endmodule

module SliceWrapper_30_18_19 (
    input [29:0] I,
    output [0:0] O
);
assign O = I[18:18];
endmodule

module SliceWrapper_30_15_18 (
    input [29:0] I,
    output [2:0] O
);
assign O = I[17:15];
endmodule

module SliceWrapper_30_14_15 (
    input [29:0] I,
    output [0:0] O
);
assign O = I[14:14];
endmodule

module SliceWrapper_30_13_14 (
    input [29:0] I,
    output [0:0] O
);
assign O = I[13:13];
endmodule

module SliceWrapper_30_10_13 (
    input [29:0] I,
    output [2:0] O
);
assign O = I[12:10];
endmodule

module SliceWrapper_30_0_30 (
    input [29:0] I,
    output [29:0] O
);
assign O = I;
endmodule

module SliceWrapper_30_0_3 (
    input [29:0] I,
    output [2:0] O
);
assign O = I[2:0];
endmodule

module SliceWrapper_25_9_10 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[9:9];
endmodule

module SliceWrapper_25_8_9 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[8:8];
endmodule

module SliceWrapper_25_7_8 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[7:7];
endmodule

module SliceWrapper_25_6_7 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[6:6];
endmodule

module SliceWrapper_25_5_6 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[5:5];
endmodule

module SliceWrapper_25_4_5 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[4:4];
endmodule

module SliceWrapper_25_3_4 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[3:3];
endmodule

module SliceWrapper_25_2_3 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[2:2];
endmodule

module SliceWrapper_25_24_25 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[24:24];
endmodule

module SliceWrapper_25_23_24 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[23:23];
endmodule

module SliceWrapper_25_21_23 (
    input [24:0] I,
    output [1:0] O
);
assign O = I[22:21];
endmodule

module SliceWrapper_25_20_21 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[20:20];
endmodule

module SliceWrapper_25_1_2 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[1:1];
endmodule

module SliceWrapper_25_19_20 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[19:19];
endmodule

module SliceWrapper_25_18_19 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[18:18];
endmodule

module SliceWrapper_25_17_18 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[17:17];
endmodule

module SliceWrapper_25_16_17 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[16:16];
endmodule

module SliceWrapper_25_15_16 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[15:15];
endmodule

module SliceWrapper_25_14_15 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[14:14];
endmodule

module SliceWrapper_25_13_14 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[13:13];
endmodule

module SliceWrapper_25_12_13 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[12:12];
endmodule

module SliceWrapper_25_11_12 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[11:11];
endmodule

module SliceWrapper_25_10_11 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[10:10];
endmodule

module SliceWrapper_25_0_1 (
    input [24:0] I,
    output [0:0] O
);
assign O = I[0:0];
endmodule

module SliceWrapper_24_9_10 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[9:9];
endmodule

module SliceWrapper_24_8_9 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[8:8];
endmodule

module SliceWrapper_24_7_8 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[7:7];
endmodule

module SliceWrapper_24_6_7 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[6:6];
endmodule

module SliceWrapper_24_5_6 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[5:5];
endmodule

module SliceWrapper_24_4_5 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[4:4];
endmodule

module SliceWrapper_24_3_4 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[3:3];
endmodule

module SliceWrapper_24_2_3 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[2:2];
endmodule

module SliceWrapper_24_23_24 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[23:23];
endmodule

module SliceWrapper_24_22_23 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[22:22];
endmodule

module SliceWrapper_24_21_22 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[21:21];
endmodule

module SliceWrapper_24_20_21 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[20:20];
endmodule

module SliceWrapper_24_1_2 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[1:1];
endmodule

module SliceWrapper_24_19_20 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[19:19];
endmodule

module SliceWrapper_24_18_19 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[18:18];
endmodule

module SliceWrapper_24_17_18 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[17:17];
endmodule

module SliceWrapper_24_16_17 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[16:16];
endmodule

module SliceWrapper_24_15_16 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[15:15];
endmodule

module SliceWrapper_24_14_15 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[14:14];
endmodule

module SliceWrapper_24_13_14 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[13:13];
endmodule

module SliceWrapper_24_12_13 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[12:12];
endmodule

module SliceWrapper_24_11_12 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[11:11];
endmodule

module SliceWrapper_24_10_11 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[10:10];
endmodule

module SliceWrapper_24_0_1 (
    input [23:0] I,
    output [0:0] O
);
assign O = I[0:0];
endmodule

module SliceWrapper_23_9_10 (
    input [22:0] I,
    output [0:0] O
);
assign O = I[9:9];
endmodule

module SliceWrapper_23_8_9 (
    input [22:0] I,
    output [0:0] O
);
assign O = I[8:8];
endmodule

module SliceWrapper_23_5_8 (
    input [22:0] I,
    output [2:0] O
);
assign O = I[7:5];
endmodule

module SliceWrapper_23_4_5 (
    input [22:0] I,
    output [0:0] O
);
assign O = I[4:4];
endmodule

module SliceWrapper_23_3_4 (
    input [22:0] I,
    output [0:0] O
);
assign O = I[3:3];
endmodule

module SliceWrapper_23_20_23 (
    input [22:0] I,
    output [2:0] O
);
assign O = I[22:20];
endmodule

module SliceWrapper_23_19_20 (
    input [22:0] I,
    output [0:0] O
);
assign O = I[19:19];
endmodule

module SliceWrapper_23_18_19 (
    input [22:0] I,
    output [0:0] O
);
assign O = I[18:18];
endmodule

module SliceWrapper_23_15_18 (
    input [22:0] I,
    output [2:0] O
);
assign O = I[17:15];
endmodule

module SliceWrapper_23_14_15 (
    input [22:0] I,
    output [0:0] O
);
assign O = I[14:14];
endmodule

module SliceWrapper_23_13_14 (
    input [22:0] I,
    output [0:0] O
);
assign O = I[13:13];
endmodule

module SliceWrapper_23_10_13 (
    input [22:0] I,
    output [2:0] O
);
assign O = I[12:10];
endmodule

module SliceWrapper_23_0_3 (
    input [22:0] I,
    output [2:0] O
);
assign O = I[2:0];
endmodule

module SliceWrapper_20_9_10 (
    input [19:0] I,
    output [0:0] O
);
assign O = I[9:9];
endmodule

module SliceWrapper_20_8_9 (
    input [19:0] I,
    output [0:0] O
);
assign O = I[8:8];
endmodule

module SliceWrapper_20_7_8 (
    input [19:0] I,
    output [0:0] O
);
assign O = I[7:7];
endmodule

module SliceWrapper_20_6_7 (
    input [19:0] I,
    output [0:0] O
);
assign O = I[6:6];
endmodule

module SliceWrapper_20_5_6 (
    input [19:0] I,
    output [0:0] O
);
assign O = I[5:5];
endmodule

module SliceWrapper_20_4_5 (
    input [19:0] I,
    output [0:0] O
);
assign O = I[4:4];
endmodule

module SliceWrapper_20_3_4 (
    input [19:0] I,
    output [0:0] O
);
assign O = I[3:3];
endmodule

module SliceWrapper_20_2_3 (
    input [19:0] I,
    output [0:0] O
);
assign O = I[2:2];
endmodule

module SliceWrapper_20_1_2 (
    input [19:0] I,
    output [0:0] O
);
assign O = I[1:1];
endmodule

module SliceWrapper_20_19_20 (
    input [19:0] I,
    output [0:0] O
);
assign O = I[19:19];
endmodule

module SliceWrapper_20_16_19 (
    input [19:0] I,
    output [2:0] O
);
assign O = I[18:16];
endmodule

module SliceWrapper_20_15_16 (
    input [19:0] I,
    output [0:0] O
);
assign O = I[15:15];
endmodule

module SliceWrapper_20_14_15 (
    input [19:0] I,
    output [0:0] O
);
assign O = I[14:14];
endmodule

module SliceWrapper_20_13_14 (
    input [19:0] I,
    output [0:0] O
);
assign O = I[13:13];
endmodule

module SliceWrapper_20_12_13 (
    input [19:0] I,
    output [0:0] O
);
assign O = I[12:12];
endmodule

module SliceWrapper_20_11_12 (
    input [19:0] I,
    output [0:0] O
);
assign O = I[11:11];
endmodule

module SliceWrapper_20_10_11 (
    input [19:0] I,
    output [0:0] O
);
assign O = I[10:10];
endmodule

module SliceWrapper_20_0_1 (
    input [19:0] I,
    output [0:0] O
);
assign O = I[0:0];
endmodule

module SliceWrapper_1_0_1 (
    input [0:0] I,
    output [0:0] O
);
assign O = I;
endmodule

module SliceWrapper_19_0_19 (
    input [18:0] I,
    output [18:0] O
);
assign O = I;
endmodule

module SliceWrapper_16_0_16 (
    input [15:0] I,
    output [15:0] O
);
assign O = I;
endmodule

module Register_unq9 (
    input [23:0] I,
    output [23:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [23:0] reg_PR24_inst0__CE_out;
regCE_arst #(
    .init(24'h000000),
    .width(24)
) reg_PR24_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR24_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR24_inst0__CE_out;
endmodule

module Register_unq8 (
    input [24:0] I,
    output [24:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [24:0] reg_PR25_inst0__CE_out;
regCE_arst #(
    .init(25'h0000000),
    .width(25)
) reg_PR25_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR25_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR25_inst0__CE_out;
endmodule

module Register_unq7 (
    input [18:0] I,
    output [18:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [18:0] reg_PR19_inst0__CE_out;
regCE_arst #(
    .init(19'h00000),
    .width(19)
) reg_PR19_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR19_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR19_inst0__CE_out;
endmodule

module Register_unq6 (
    input [22:0] I,
    output [22:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [22:0] reg_PR23_inst0__CE_out;
regCE_arst #(
    .init(23'h000000),
    .width(23)
) reg_PR23_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR23_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR23_inst0__CE_out;
endmodule

module Register_unq5 (
    input [30:0] I,
    output [30:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [30:0] reg_PR31_inst0__CE_out;
regCE_arst #(
    .init(31'h00000000),
    .width(31)
) reg_PR31_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR31_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR31_inst0__CE_out;
endmodule

module Register_unq4 (
    input [0:0] I,
    output [0:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [0:0] reg_PR1_inst0__CE_out;
regCE_arst #(
    .init(1'h0),
    .width(1)
) reg_PR1_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR1_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR1_inst0__CE_out;
endmodule

module Register_unq3 (
    input [29:0] I,
    output [29:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [29:0] reg_PR30_inst0__CE_out;
regCE_arst #(
    .init(30'h00000000),
    .width(30)
) reg_PR30_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR30_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR30_inst0__CE_out;
endmodule

module Register_unq2 (
    input [5:0] I,
    output [5:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [5:0] reg_PR6_inst0__CE_out;
regCE_arst #(
    .init(6'h00),
    .width(6)
) reg_PR6_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR6_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR6_inst0__CE_out;
endmodule

module Register_unq1 (
    input [19:0] I,
    output [19:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [19:0] reg_PR20_inst0__CE_out;
regCE_arst #(
    .init(20'h00000),
    .width(20)
) reg_PR20_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR20_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR20_inst0__CE_out;
endmodule

module Register (
    input [31:0] I,
    output [31:0] O,
    input CE,
    input CLK,
    input ASYNCRESET
);
wire [31:0] reg_PR32_inst0__CE_out;
regCE_arst #(
    .init(32'h00000000),
    .width(32)
) reg_PR32_inst0__CE (
    .in(I),
    .ce(CE),
    .out(reg_PR32_inst0__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = reg_PR32_inst0__CE_out;
endmodule

module ReadyValidLoopBack (
  input logic ready_in,
  input logic valid_in,
  output logic valid_out
);

assign valid_out = ready_in & valid_in;
endmodule   // ReadyValidLoopBack


module PowerDomainOR (
    input [31:0] I0,
    input [31:0] I1,
    output [31:0] O,
    input [0:0] I_not
);
wire [0:0] Invert1_inst0_out;
wire [0:0] and1_inst0_out;
wire [0:0] and1_inst1_out;
wire [0:0] and1_inst10_out;
wire [0:0] and1_inst11_out;
wire [0:0] and1_inst12_out;
wire [0:0] and1_inst13_out;
wire [0:0] and1_inst14_out;
wire [0:0] and1_inst15_out;
wire [0:0] and1_inst16_out;
wire [0:0] and1_inst17_out;
wire [0:0] and1_inst18_out;
wire [0:0] and1_inst19_out;
wire [0:0] and1_inst2_out;
wire [0:0] and1_inst20_out;
wire [0:0] and1_inst21_out;
wire [0:0] and1_inst22_out;
wire [0:0] and1_inst23_out;
wire [0:0] and1_inst24_out;
wire [0:0] and1_inst25_out;
wire [0:0] and1_inst26_out;
wire [0:0] and1_inst27_out;
wire [0:0] and1_inst28_out;
wire [0:0] and1_inst29_out;
wire [0:0] and1_inst3_out;
wire [0:0] and1_inst30_out;
wire [0:0] and1_inst31_out;
wire [0:0] and1_inst4_out;
wire [0:0] and1_inst5_out;
wire [0:0] and1_inst6_out;
wire [0:0] and1_inst7_out;
wire [0:0] and1_inst8_out;
wire [0:0] and1_inst9_out;
wire [31:0] or32_inst0_out;
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(I_not),
    .out(Invert1_inst0_out)
);
coreir_and #(
    .width(1)
) and1_inst0 (
    .in0(I0[0]),
    .in1(Invert1_inst0_out),
    .out(and1_inst0_out)
);
coreir_and #(
    .width(1)
) and1_inst1 (
    .in0(I0[1]),
    .in1(Invert1_inst0_out),
    .out(and1_inst1_out)
);
coreir_and #(
    .width(1)
) and1_inst10 (
    .in0(I0[10]),
    .in1(Invert1_inst0_out),
    .out(and1_inst10_out)
);
coreir_and #(
    .width(1)
) and1_inst11 (
    .in0(I0[11]),
    .in1(Invert1_inst0_out),
    .out(and1_inst11_out)
);
coreir_and #(
    .width(1)
) and1_inst12 (
    .in0(I0[12]),
    .in1(Invert1_inst0_out),
    .out(and1_inst12_out)
);
coreir_and #(
    .width(1)
) and1_inst13 (
    .in0(I0[13]),
    .in1(Invert1_inst0_out),
    .out(and1_inst13_out)
);
coreir_and #(
    .width(1)
) and1_inst14 (
    .in0(I0[14]),
    .in1(Invert1_inst0_out),
    .out(and1_inst14_out)
);
coreir_and #(
    .width(1)
) and1_inst15 (
    .in0(I0[15]),
    .in1(Invert1_inst0_out),
    .out(and1_inst15_out)
);
coreir_and #(
    .width(1)
) and1_inst16 (
    .in0(I0[16]),
    .in1(Invert1_inst0_out),
    .out(and1_inst16_out)
);
coreir_and #(
    .width(1)
) and1_inst17 (
    .in0(I0[17]),
    .in1(Invert1_inst0_out),
    .out(and1_inst17_out)
);
coreir_and #(
    .width(1)
) and1_inst18 (
    .in0(I0[18]),
    .in1(Invert1_inst0_out),
    .out(and1_inst18_out)
);
coreir_and #(
    .width(1)
) and1_inst19 (
    .in0(I0[19]),
    .in1(Invert1_inst0_out),
    .out(and1_inst19_out)
);
coreir_and #(
    .width(1)
) and1_inst2 (
    .in0(I0[2]),
    .in1(Invert1_inst0_out),
    .out(and1_inst2_out)
);
coreir_and #(
    .width(1)
) and1_inst20 (
    .in0(I0[20]),
    .in1(Invert1_inst0_out),
    .out(and1_inst20_out)
);
coreir_and #(
    .width(1)
) and1_inst21 (
    .in0(I0[21]),
    .in1(Invert1_inst0_out),
    .out(and1_inst21_out)
);
coreir_and #(
    .width(1)
) and1_inst22 (
    .in0(I0[22]),
    .in1(Invert1_inst0_out),
    .out(and1_inst22_out)
);
coreir_and #(
    .width(1)
) and1_inst23 (
    .in0(I0[23]),
    .in1(Invert1_inst0_out),
    .out(and1_inst23_out)
);
coreir_and #(
    .width(1)
) and1_inst24 (
    .in0(I0[24]),
    .in1(Invert1_inst0_out),
    .out(and1_inst24_out)
);
coreir_and #(
    .width(1)
) and1_inst25 (
    .in0(I0[25]),
    .in1(Invert1_inst0_out),
    .out(and1_inst25_out)
);
coreir_and #(
    .width(1)
) and1_inst26 (
    .in0(I0[26]),
    .in1(Invert1_inst0_out),
    .out(and1_inst26_out)
);
coreir_and #(
    .width(1)
) and1_inst27 (
    .in0(I0[27]),
    .in1(Invert1_inst0_out),
    .out(and1_inst27_out)
);
coreir_and #(
    .width(1)
) and1_inst28 (
    .in0(I0[28]),
    .in1(Invert1_inst0_out),
    .out(and1_inst28_out)
);
coreir_and #(
    .width(1)
) and1_inst29 (
    .in0(I0[29]),
    .in1(Invert1_inst0_out),
    .out(and1_inst29_out)
);
coreir_and #(
    .width(1)
) and1_inst3 (
    .in0(I0[3]),
    .in1(Invert1_inst0_out),
    .out(and1_inst3_out)
);
coreir_and #(
    .width(1)
) and1_inst30 (
    .in0(I0[30]),
    .in1(Invert1_inst0_out),
    .out(and1_inst30_out)
);
coreir_and #(
    .width(1)
) and1_inst31 (
    .in0(I0[31]),
    .in1(Invert1_inst0_out),
    .out(and1_inst31_out)
);
coreir_and #(
    .width(1)
) and1_inst4 (
    .in0(I0[4]),
    .in1(Invert1_inst0_out),
    .out(and1_inst4_out)
);
coreir_and #(
    .width(1)
) and1_inst5 (
    .in0(I0[5]),
    .in1(Invert1_inst0_out),
    .out(and1_inst5_out)
);
coreir_and #(
    .width(1)
) and1_inst6 (
    .in0(I0[6]),
    .in1(Invert1_inst0_out),
    .out(and1_inst6_out)
);
coreir_and #(
    .width(1)
) and1_inst7 (
    .in0(I0[7]),
    .in1(Invert1_inst0_out),
    .out(and1_inst7_out)
);
coreir_and #(
    .width(1)
) and1_inst8 (
    .in0(I0[8]),
    .in1(Invert1_inst0_out),
    .out(and1_inst8_out)
);
coreir_and #(
    .width(1)
) and1_inst9 (
    .in0(I0[9]),
    .in1(Invert1_inst0_out),
    .out(and1_inst9_out)
);
wire [31:0] or32_inst0_in0;
assign or32_inst0_in0 = {and1_inst31_out[0],and1_inst30_out[0],and1_inst29_out[0],and1_inst28_out[0],and1_inst27_out[0],and1_inst26_out[0],and1_inst25_out[0],and1_inst24_out[0],and1_inst23_out[0],and1_inst22_out[0],and1_inst21_out[0],and1_inst20_out[0],and1_inst19_out[0],and1_inst18_out[0],and1_inst17_out[0],and1_inst16_out[0],and1_inst15_out[0],and1_inst14_out[0],and1_inst13_out[0],and1_inst12_out[0],and1_inst11_out[0],and1_inst10_out[0],and1_inst9_out[0],and1_inst8_out[0],and1_inst7_out[0],and1_inst6_out[0],and1_inst5_out[0],and1_inst4_out[0],and1_inst3_out[0],and1_inst2_out[0],and1_inst1_out[0],and1_inst0_out[0]};
coreir_or #(
    .width(32)
) or32_inst0 (
    .in0(or32_inst0_in0),
    .in1(I1),
    .out(or32_inst0_out)
);
assign O = or32_inst0_out;
endmodule

module PondTop (
  input logic [31:0] CONFIG_SPACE_0,
  input logic [31:0] CONFIG_SPACE_1,
  input logic [31:0] CONFIG_SPACE_10,
  input logic [31:0] CONFIG_SPACE_11,
  input logic [31:0] CONFIG_SPACE_12,
  input logic [31:0] CONFIG_SPACE_13,
  input logic [31:0] CONFIG_SPACE_14,
  input logic [31:0] CONFIG_SPACE_15,
  input logic [29:0] CONFIG_SPACE_16,
  input logic [31:0] CONFIG_SPACE_2,
  input logic [31:0] CONFIG_SPACE_3,
  input logic [31:0] CONFIG_SPACE_4,
  input logic [31:0] CONFIG_SPACE_5,
  input logic [31:0] CONFIG_SPACE_6,
  input logic [31:0] CONFIG_SPACE_7,
  input logic [31:0] CONFIG_SPACE_8,
  input logic [31:0] CONFIG_SPACE_9,
  input logic [0:0] [16:0] PondTop_input_width_17_num_0,
  input logic [0:0] [16:0] PondTop_input_width_17_num_1,
  input logic clk,
  input logic clk_en,
  input logic [7:0] config_addr_in,
  input logic [31:0] config_data_in,
  input logic config_en,
  input logic config_read,
  input logic config_write,
  input logic flush,
  input logic rst_n,
  input logic tile_en,
  output logic [0:0] [16:0] PondTop_output_width_17_num_0,
  output logic [0:0] [16:0] PondTop_output_width_17_num_1,
  output logic PondTop_output_width_1_num_0,
  output logic PondTop_output_width_1_num_1,
  output logic [0:0] [31:0] config_data_out
);

logic [541:0] CONFIG_SPACE;
logic [15:0] config_data_in_shrt;
logic [0:0][15:0] config_data_out_shrt;
logic [4:0] config_seq_addr_out;
logic config_seq_clk_en;
logic [0:0][0:0][15:0] config_seq_rd_data_stg;
logic config_seq_ren_out;
logic config_seq_wen_out;
logic [0:0][15:0] config_seq_wr_data;
logic gclk;
logic mem_ctrl_strg_ub_thin_flat_clk;
logic [0:0][16:0] mem_ctrl_strg_ub_thin_flat_data_out_f_0;
logic [0:0][16:0] mem_ctrl_strg_ub_thin_flat_data_out_f_1;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_data_from_strg_lifted;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_data_to_strg_lifted;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_starting_addr;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_starting_addr2;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_strides2_0;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_strides2_1;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_strides_0;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_strides_1;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_strides_2;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_strides_3;
logic [2:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_dimensionality;
logic [1:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_dimensionality2;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_ranges2_0;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_ranges2_1;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_ranges_0;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_ranges_1;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_ranges_2;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_ranges_3;
logic mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_enable;
logic mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_enable2;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr2;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_0;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_1;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_0;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_1;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_2;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_3;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_rd_addr_out_lifted;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_starting_addr;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_starting_addr2;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_strides2_0;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_strides2_1;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_strides_0;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_strides_1;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_strides_2;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_strides_3;
logic [2:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_dimensionality;
logic [1:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_dimensionality2;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_ranges2_0;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_ranges2_1;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_ranges_0;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_ranges_1;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_ranges_2;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_ranges_3;
logic mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_enable;
logic mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_enable2;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr2;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_0;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_1;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_0;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_1;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_2;
logic [15:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_3;
logic mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_ren_to_strg_lifted;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_tmp0_rdaddr_lifted;
logic mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_tmp0_rden_lifted;
logic mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_wen_to_strg_lifted;
logic [4:0] mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_wr_addr_out_lifted;
logic mem_ctrl_strg_ub_thin_flat_valid_out_f_b_0;
logic mem_ctrl_strg_ub_thin_flat_valid_out_f_b_1;
logic memory_0_clk_en;
logic [15:0] memory_0_data_in_p0;
logic [15:0] memory_0_data_out_p0;
logic [4:0] memory_0_read_addr_p0;
logic [4:0] memory_0_read_addr_p1;
logic memory_0_read_enable_p0;
logic memory_0_read_enable_p1;
logic [4:0] memory_0_write_addr_p0;
logic memory_0_write_enable_p0;
logic mode;
assign mode = 1'h0;
assign gclk = clk & tile_en;
assign mem_ctrl_strg_ub_thin_flat_clk = gclk;
always_comb begin
  PondTop_output_width_17_num_0 = 17'h0;
  if (1'h0 == mode) begin
    PondTop_output_width_17_num_0 = mem_ctrl_strg_ub_thin_flat_data_out_f_0;
  end
  else PondTop_output_width_17_num_0 = 17'h0;
end
always_comb begin
  PondTop_output_width_17_num_1 = 17'h0;
  if (1'h0 == mode) begin
    PondTop_output_width_17_num_1 = mem_ctrl_strg_ub_thin_flat_data_out_f_1;
  end
  else PondTop_output_width_17_num_1 = 17'h0;
end
always_comb begin
  PondTop_output_width_1_num_0 = 1'h0;
  if (1'h0 == mode) begin
    PondTop_output_width_1_num_0 = mem_ctrl_strg_ub_thin_flat_valid_out_f_b_0;
  end
  else PondTop_output_width_1_num_0 = 1'h0;
end
always_comb begin
  PondTop_output_width_1_num_1 = 1'h0;
  if (1'h0 == mode) begin
    PondTop_output_width_1_num_1 = mem_ctrl_strg_ub_thin_flat_valid_out_f_b_1;
  end
  else PondTop_output_width_1_num_1 = 1'h0;
end
always_comb begin
  memory_0_data_in_p0 = 16'h0;
  memory_0_write_addr_p0 = 5'h0;
  memory_0_write_enable_p0 = 1'h0;
  memory_0_read_addr_p0 = 5'h0;
  memory_0_read_enable_p0 = 1'h0;
  if (|config_en) begin
    memory_0_data_in_p0 = config_seq_wr_data;
    memory_0_write_addr_p0 = config_seq_addr_out;
    memory_0_write_enable_p0 = config_seq_wen_out;
    memory_0_read_addr_p0 = config_seq_addr_out;
    memory_0_read_enable_p0 = config_seq_ren_out;
  end
  else if (1'h0 == mode) begin
    memory_0_data_in_p0 = mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_data_to_strg_lifted;
    memory_0_write_addr_p0 = mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_wr_addr_out_lifted;
    memory_0_write_enable_p0 = mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_wen_to_strg_lifted;
    memory_0_read_addr_p0 = mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_rd_addr_out_lifted;
    memory_0_read_enable_p0 = mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_ren_to_strg_lifted;
  end
end
always_comb begin
  mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_data_from_strg_lifted = memory_0_data_out_p0;
  config_seq_rd_data_stg = memory_0_data_out_p0;
end
always_comb begin
  memory_0_read_addr_p1 = 5'h0;
  memory_0_read_enable_p1 = 1'h0;
  if (1'h0 == mode) begin
    memory_0_read_addr_p1 = mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_tmp0_rdaddr_lifted;
    memory_0_read_enable_p1 = mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_tmp0_rden_lifted;
  end
end
assign config_data_in_shrt = config_data_in[15:0];
assign config_data_out[0] = 32'(config_data_out_shrt[0]);
assign config_seq_clk_en = clk_en | (|config_en);
assign memory_0_clk_en = clk_en | (|config_en);
assign {mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_starting_addr, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_starting_addr2, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_strides2_0, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_strides2_1, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_strides_0, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_strides_1, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_strides_2, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_strides_3, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_dimensionality, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_dimensionality2, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_ranges2_0, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_ranges2_1, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_ranges_0, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_ranges_1, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_ranges_2, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_ranges_3, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_enable, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_enable2, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr2, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_0, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_1, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_0, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_1, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_2, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_3, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_starting_addr, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_starting_addr2, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_strides2_0, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_strides2_1, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_strides_0, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_strides_1, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_strides_2, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_strides_3, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_dimensionality, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_dimensionality2, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_ranges2_0, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_ranges2_1, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_ranges_0, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_ranges_1, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_ranges_2, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_ranges_3, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_enable, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_enable2, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr2, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_0, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_1, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_0, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_1, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_2, mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_3} = CONFIG_SPACE[541:0];
assign CONFIG_SPACE[31:0] = CONFIG_SPACE_0;
assign CONFIG_SPACE[63:32] = CONFIG_SPACE_1;
assign CONFIG_SPACE[95:64] = CONFIG_SPACE_2;
assign CONFIG_SPACE[127:96] = CONFIG_SPACE_3;
assign CONFIG_SPACE[159:128] = CONFIG_SPACE_4;
assign CONFIG_SPACE[191:160] = CONFIG_SPACE_5;
assign CONFIG_SPACE[223:192] = CONFIG_SPACE_6;
assign CONFIG_SPACE[255:224] = CONFIG_SPACE_7;
assign CONFIG_SPACE[287:256] = CONFIG_SPACE_8;
assign CONFIG_SPACE[319:288] = CONFIG_SPACE_9;
assign CONFIG_SPACE[351:320] = CONFIG_SPACE_10;
assign CONFIG_SPACE[383:352] = CONFIG_SPACE_11;
assign CONFIG_SPACE[415:384] = CONFIG_SPACE_12;
assign CONFIG_SPACE[447:416] = CONFIG_SPACE_13;
assign CONFIG_SPACE[479:448] = CONFIG_SPACE_14;
assign CONFIG_SPACE[511:480] = CONFIG_SPACE_15;
assign CONFIG_SPACE[541:512] = CONFIG_SPACE_16;
strg_ub_thin_flat mem_ctrl_strg_ub_thin_flat (
  .clk(mem_ctrl_strg_ub_thin_flat_clk),
  .clk_en(clk_en),
  .data_in_f_0(PondTop_input_width_17_num_0),
  .data_in_f_1(PondTop_input_width_17_num_1),
  .flush(flush),
  .rst_n(rst_n),
  .strg_ub_thin_inst_data_from_strg_lifted(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_data_from_strg_lifted),
  .strg_ub_thin_inst_in2regfile_0_addr_gen_starting_addr(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_starting_addr),
  .strg_ub_thin_inst_in2regfile_0_addr_gen_starting_addr2(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_starting_addr2),
  .strg_ub_thin_inst_in2regfile_0_addr_gen_strides2_0(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_strides2_0),
  .strg_ub_thin_inst_in2regfile_0_addr_gen_strides2_1(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_strides2_1),
  .strg_ub_thin_inst_in2regfile_0_addr_gen_strides_0(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_strides_0),
  .strg_ub_thin_inst_in2regfile_0_addr_gen_strides_1(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_strides_1),
  .strg_ub_thin_inst_in2regfile_0_addr_gen_strides_2(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_strides_2),
  .strg_ub_thin_inst_in2regfile_0_addr_gen_strides_3(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_addr_gen_strides_3),
  .strg_ub_thin_inst_in2regfile_0_for_loop_dimensionality(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_dimensionality),
  .strg_ub_thin_inst_in2regfile_0_for_loop_dimensionality2(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_dimensionality2),
  .strg_ub_thin_inst_in2regfile_0_for_loop_ranges2_0(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_ranges2_0),
  .strg_ub_thin_inst_in2regfile_0_for_loop_ranges2_1(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_ranges2_1),
  .strg_ub_thin_inst_in2regfile_0_for_loop_ranges_0(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_ranges_0),
  .strg_ub_thin_inst_in2regfile_0_for_loop_ranges_1(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_ranges_1),
  .strg_ub_thin_inst_in2regfile_0_for_loop_ranges_2(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_ranges_2),
  .strg_ub_thin_inst_in2regfile_0_for_loop_ranges_3(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_for_loop_ranges_3),
  .strg_ub_thin_inst_in2regfile_0_sched_gen_enable(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_enable),
  .strg_ub_thin_inst_in2regfile_0_sched_gen_enable2(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_enable2),
  .strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr),
  .strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr2(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr2),
  .strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_0(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_0),
  .strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_1(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_1),
  .strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_0(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_0),
  .strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_1(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_1),
  .strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_2(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_2),
  .strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_3(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_3),
  .strg_ub_thin_inst_regfile2out_0_addr_gen_starting_addr(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_starting_addr),
  .strg_ub_thin_inst_regfile2out_0_addr_gen_starting_addr2(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_starting_addr2),
  .strg_ub_thin_inst_regfile2out_0_addr_gen_strides2_0(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_strides2_0),
  .strg_ub_thin_inst_regfile2out_0_addr_gen_strides2_1(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_strides2_1),
  .strg_ub_thin_inst_regfile2out_0_addr_gen_strides_0(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_strides_0),
  .strg_ub_thin_inst_regfile2out_0_addr_gen_strides_1(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_strides_1),
  .strg_ub_thin_inst_regfile2out_0_addr_gen_strides_2(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_strides_2),
  .strg_ub_thin_inst_regfile2out_0_addr_gen_strides_3(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_addr_gen_strides_3),
  .strg_ub_thin_inst_regfile2out_0_for_loop_dimensionality(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_dimensionality),
  .strg_ub_thin_inst_regfile2out_0_for_loop_dimensionality2(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_dimensionality2),
  .strg_ub_thin_inst_regfile2out_0_for_loop_ranges2_0(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_ranges2_0),
  .strg_ub_thin_inst_regfile2out_0_for_loop_ranges2_1(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_ranges2_1),
  .strg_ub_thin_inst_regfile2out_0_for_loop_ranges_0(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_ranges_0),
  .strg_ub_thin_inst_regfile2out_0_for_loop_ranges_1(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_ranges_1),
  .strg_ub_thin_inst_regfile2out_0_for_loop_ranges_2(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_ranges_2),
  .strg_ub_thin_inst_regfile2out_0_for_loop_ranges_3(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_for_loop_ranges_3),
  .strg_ub_thin_inst_regfile2out_0_sched_gen_enable(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_enable),
  .strg_ub_thin_inst_regfile2out_0_sched_gen_enable2(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_enable2),
  .strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr),
  .strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr2(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr2),
  .strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_0(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_0),
  .strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_1(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_1),
  .strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_0(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_0),
  .strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_1(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_1),
  .strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_2(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_2),
  .strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_3(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_3),
  .data_out_f_0(mem_ctrl_strg_ub_thin_flat_data_out_f_0),
  .data_out_f_1(mem_ctrl_strg_ub_thin_flat_data_out_f_1),
  .strg_ub_thin_inst_data_to_strg_lifted(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_data_to_strg_lifted),
  .strg_ub_thin_inst_rd_addr_out_lifted(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_rd_addr_out_lifted),
  .strg_ub_thin_inst_ren_to_strg_lifted(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_ren_to_strg_lifted),
  .strg_ub_thin_inst_tmp0_rdaddr_lifted(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_tmp0_rdaddr_lifted),
  .strg_ub_thin_inst_tmp0_rden_lifted(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_tmp0_rden_lifted),
  .strg_ub_thin_inst_wen_to_strg_lifted(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_wen_to_strg_lifted),
  .strg_ub_thin_inst_wr_addr_out_lifted(mem_ctrl_strg_ub_thin_flat_strg_ub_thin_inst_wr_addr_out_lifted),
  .valid_out_f_b_0(mem_ctrl_strg_ub_thin_flat_valid_out_f_b_0),
  .valid_out_f_b_1(mem_ctrl_strg_ub_thin_flat_valid_out_f_b_1)
);

sram_dp__0 memory_0 (
  .clk(gclk),
  .clk_en(memory_0_clk_en),
  .data_in_p0(memory_0_data_in_p0),
  .flush(flush),
  .read_addr_p0(memory_0_read_addr_p0),
  .read_addr_p1(memory_0_read_addr_p1),
  .read_enable_p0(memory_0_read_enable_p0),
  .read_enable_p1(memory_0_read_enable_p1),
  .write_addr_p0(memory_0_write_addr_p0),
  .write_enable_p0(memory_0_write_enable_p0),
  .data_out_p0(memory_0_data_out_p0)
);

storage_config_seq_1_16_16 config_seq (
  .clk(gclk),
  .clk_en(config_seq_clk_en),
  .config_addr_in(config_addr_in),
  .config_data_in(config_data_in_shrt),
  .config_en(config_en),
  .config_rd(config_read),
  .config_wr(config_write),
  .flush(flush),
  .rd_data_stg(config_seq_rd_data_stg),
  .rst_n(rst_n),
  .addr_out(config_seq_addr_out),
  .rd_data_out(config_data_out_shrt),
  .ren_out(config_seq_ren_out),
  .wen_out(config_seq_wen_out),
  .wr_data(config_seq_wr_data)
);

endmodule   // PondTop

module PondTop_W (
  input logic [31:0] CONFIG_SPACE_0,
  input logic [31:0] CONFIG_SPACE_1,
  input logic [31:0] CONFIG_SPACE_10,
  input logic [31:0] CONFIG_SPACE_11,
  input logic [31:0] CONFIG_SPACE_12,
  input logic [31:0] CONFIG_SPACE_13,
  input logic [31:0] CONFIG_SPACE_14,
  input logic [31:0] CONFIG_SPACE_15,
  input logic [29:0] CONFIG_SPACE_16,
  input logic [31:0] CONFIG_SPACE_2,
  input logic [31:0] CONFIG_SPACE_3,
  input logic [31:0] CONFIG_SPACE_4,
  input logic [31:0] CONFIG_SPACE_5,
  input logic [31:0] CONFIG_SPACE_6,
  input logic [31:0] CONFIG_SPACE_7,
  input logic [31:0] CONFIG_SPACE_8,
  input logic [31:0] CONFIG_SPACE_9,
  input logic [0:0] [16:0] PondTop_input_width_17_num_0,
  input logic [0:0] [16:0] PondTop_input_width_17_num_1,
  input logic clk,
  input logic clk_en,
  input logic [7:0] config_addr_in,
  input logic [31:0] config_data_in,
  input logic config_en,
  input logic config_read,
  input logic config_write,
  input logic flush,
  input logic rst_n,
  input logic tile_en,
  output logic [0:0] [16:0] PondTop_output_width_17_num_0,
  output logic [0:0] [16:0] PondTop_output_width_17_num_1,
  output logic PondTop_output_width_1_num_0,
  output logic PondTop_output_width_1_num_1,
  output logic [0:0] [31:0] config_data_out
);

PondTop PondTop (
  .CONFIG_SPACE_0(CONFIG_SPACE_0),
  .CONFIG_SPACE_1(CONFIG_SPACE_1),
  .CONFIG_SPACE_10(CONFIG_SPACE_10),
  .CONFIG_SPACE_11(CONFIG_SPACE_11),
  .CONFIG_SPACE_12(CONFIG_SPACE_12),
  .CONFIG_SPACE_13(CONFIG_SPACE_13),
  .CONFIG_SPACE_14(CONFIG_SPACE_14),
  .CONFIG_SPACE_15(CONFIG_SPACE_15),
  .CONFIG_SPACE_16(CONFIG_SPACE_16),
  .CONFIG_SPACE_2(CONFIG_SPACE_2),
  .CONFIG_SPACE_3(CONFIG_SPACE_3),
  .CONFIG_SPACE_4(CONFIG_SPACE_4),
  .CONFIG_SPACE_5(CONFIG_SPACE_5),
  .CONFIG_SPACE_6(CONFIG_SPACE_6),
  .CONFIG_SPACE_7(CONFIG_SPACE_7),
  .CONFIG_SPACE_8(CONFIG_SPACE_8),
  .CONFIG_SPACE_9(CONFIG_SPACE_9),
  .PondTop_input_width_17_num_0(PondTop_input_width_17_num_0),
  .PondTop_input_width_17_num_1(PondTop_input_width_17_num_1),
  .clk(clk),
  .clk_en(clk_en),
  .config_addr_in(config_addr_in),
  .config_data_in(config_data_in),
  .config_en(config_en),
  .config_read(config_read),
  .config_write(config_write),
  .flush(flush),
  .rst_n(rst_n),
  .tile_en(tile_en),
  .PondTop_output_width_17_num_0(PondTop_output_width_17_num_0),
  .PondTop_output_width_17_num_1(PondTop_output_width_17_num_1),
  .PondTop_output_width_1_num_0(PondTop_output_width_1_num_0),
  .PondTop_output_width_1_num_1(PondTop_output_width_1_num_1),
  .config_data_out(config_data_out)
);

endmodule   // PondTop_W

module addr_gen_4_16_dual_config_2 (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [2:0] mux_sel,
  input logic mux_sel_msb_init,
  input logic restart,
  input logic rst_n,
  input logic [15:0] starting_addr,
  input logic [15:0] starting_addr2,
  input logic step,
  input logic [3:0] [15:0] strides,
  input logic [1:0] [15:0] strides2,
  output logic [15:0] addr_out,
  output logic starting_addr_comp
);

logic [15:0] calc_addr;
logic [15:0] cur_stride;
logic [15:0] current_addr;
logic [15:0] flush_addr;
logic [1:0] mux_sel_iter1;
logic mux_sel_iter2;
logic mux_sel_msb;
logic [15:0] restart_addr;
logic [15:0] strt_addr;
assign starting_addr_comp = starting_addr2 < starting_addr;
assign mux_sel_iter1 = mux_sel[1:0];
assign mux_sel_iter2 = mux_sel[0];
assign mux_sel_msb = mux_sel[2];
assign flush_addr = mux_sel_msb_init ? starting_addr2: starting_addr;
assign strt_addr = mux_sel_msb ? starting_addr2: starting_addr;
assign restart_addr = (~mux_sel_msb) ? starting_addr2: starting_addr;
assign cur_stride = mux_sel_msb ? strides2[mux_sel_iter2]: strides[mux_sel_iter1];
assign addr_out = calc_addr;
assign calc_addr = current_addr;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    current_addr <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      current_addr <= flush_addr;
    end
    else if (step) begin
      if (restart) begin
        current_addr <= restart_addr;
      end
      else current_addr <= current_addr + cur_stride;
    end
  end
end
endmodule   // addr_gen_4_16_dual_config_2

module addr_gen_4_5_dual_config_2 (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [2:0] mux_sel,
  input logic mux_sel_msb_init,
  input logic restart,
  input logic rst_n,
  input logic [4:0] starting_addr,
  input logic [4:0] starting_addr2,
  input logic step,
  input logic [3:0] [4:0] strides,
  input logic [1:0] [4:0] strides2,
  output logic [4:0] addr_out,
  output logic starting_addr_comp
);

logic [4:0] calc_addr;
logic [4:0] cur_stride;
logic [4:0] current_addr;
logic [4:0] flush_addr;
logic [1:0] mux_sel_iter1;
logic mux_sel_iter2;
logic mux_sel_msb;
logic [4:0] restart_addr;
logic [4:0] strt_addr;
assign starting_addr_comp = starting_addr2 < starting_addr;
assign mux_sel_iter1 = mux_sel[1:0];
assign mux_sel_iter2 = mux_sel[0];
assign mux_sel_msb = mux_sel[2];
assign flush_addr = mux_sel_msb_init ? starting_addr2: starting_addr;
assign strt_addr = mux_sel_msb ? starting_addr2: starting_addr;
assign restart_addr = (~mux_sel_msb) ? starting_addr2: starting_addr;
assign cur_stride = mux_sel_msb ? strides2[mux_sel_iter2]: strides[mux_sel_iter1];
assign addr_out = calc_addr;
assign calc_addr = current_addr;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    current_addr <= 5'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      current_addr <= flush_addr;
    end
    else if (step) begin
      if (restart) begin
        current_addr <= restart_addr;
      end
      else current_addr <= current_addr + cur_stride;
    end
  end
end
endmodule   // addr_gen_4_5_dual_config_2

module for_loop_dual_config_4_2_16 #(
  parameter CONFIG_WIDTH = 5'h10,
  parameter ITERATOR_SUPPORT = 3'h4,
  parameter ITERATOR_SUPPORT2 = 2'h2
)
(
  input logic clk,
  input logic clk_en,
  input logic [2:0] dimensionality,
  input logic [1:0] dimensionality2,
  input logic flush,
  input logic mux_sel_msb_init,
  input logic [3:0] [15:0] ranges,
  input logic [1:0] [15:0] ranges2,
  input logic rst_n,
  input logic step,
  output logic [2:0] mux_sel_out,
  output logic restart
);

logic [3:0] clear;
logic [2:0] cur_dimensionality;
logic [15:0] cur_range;
logic [3:0][15:0] dim_counter;
logic done;
logic [3:0] inc;
logic [15:0] inced_cnt;
logic [3:0] max_value;
logic maxed_value;
logic [1:0] mux_sel;
logic [1:0] mux_sel_iter1;
logic mux_sel_iter2;
logic mux_sel_msb;
logic mux_sel_msb_r;
assign mux_sel_msb = mux_sel_msb_r;
assign cur_dimensionality = mux_sel_msb ? 3'(dimensionality2): dimensionality;
assign mux_sel_iter1 = mux_sel[1:0];
assign mux_sel_iter2 = mux_sel[0];
assign mux_sel_out = {mux_sel_msb, mux_sel};
assign inced_cnt = dim_counter[mux_sel] + 16'h1;
assign cur_range = mux_sel_msb ? ranges2[mux_sel_iter2]: ranges[mux_sel_iter1];
assign maxed_value = (dim_counter[mux_sel] == cur_range) & inc[mux_sel];
always_comb begin
  mux_sel = 2'h0;
  done = 1'h0;
  if (~done) begin
    if ((~max_value[0]) & (cur_dimensionality > 3'h0)) begin
      mux_sel = 2'h0;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[1]) & (cur_dimensionality > 3'h1)) begin
      mux_sel = 2'h1;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[2]) & (cur_dimensionality > 3'h2)) begin
      mux_sel = 2'h2;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[3]) & (cur_dimensionality > 3'h3)) begin
      mux_sel = 2'h3;
      done = 1'h1;
    end
  end
end
always_comb begin
  clear[0] = 1'h0;
  if (((mux_sel > 2'h0) | (~done)) & step) begin
    clear[0] = 1'h1;
  end
end
always_comb begin
  inc[0] = 1'h0;
  if ((5'h0 == 5'h0) & step & (cur_dimensionality > 3'h0)) begin
    inc[0] = 1'h1;
  end
  else if ((mux_sel == 2'h0) & step & (cur_dimensionality > 3'h0)) begin
    inc[0] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[0] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[0] <= 16'h0;
    end
    else if (clear[0]) begin
      dim_counter[0] <= 16'h0;
    end
    else if (inc[0]) begin
      dim_counter[0] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[0] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[0] <= 1'h0;
    end
    else if (clear[0]) begin
      max_value[0] <= 1'h0;
    end
    else if (inc[0]) begin
      max_value[0] <= maxed_value;
    end
  end
end
always_comb begin
  clear[1] = 1'h0;
  if (((mux_sel > 2'h1) | (~done)) & step) begin
    clear[1] = 1'h1;
  end
end
always_comb begin
  inc[1] = 1'h0;
  if ((5'h1 == 5'h0) & step & (cur_dimensionality > 3'h1)) begin
    inc[1] = 1'h1;
  end
  else if ((mux_sel == 2'h1) & step & (cur_dimensionality > 3'h1)) begin
    inc[1] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[1] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[1] <= 16'h0;
    end
    else if (clear[1]) begin
      dim_counter[1] <= 16'h0;
    end
    else if (inc[1]) begin
      dim_counter[1] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[1] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[1] <= 1'h0;
    end
    else if (clear[1]) begin
      max_value[1] <= 1'h0;
    end
    else if (inc[1]) begin
      max_value[1] <= maxed_value;
    end
  end
end
always_comb begin
  clear[2] = 1'h0;
  if (((mux_sel > 2'h2) | (~done)) & step) begin
    clear[2] = 1'h1;
  end
end
always_comb begin
  inc[2] = 1'h0;
  if ((5'h2 == 5'h0) & step & (cur_dimensionality > 3'h2)) begin
    inc[2] = 1'h1;
  end
  else if ((mux_sel == 2'h2) & step & (cur_dimensionality > 3'h2)) begin
    inc[2] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[2] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[2] <= 16'h0;
    end
    else if (clear[2]) begin
      dim_counter[2] <= 16'h0;
    end
    else if (inc[2]) begin
      dim_counter[2] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[2] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[2] <= 1'h0;
    end
    else if (clear[2]) begin
      max_value[2] <= 1'h0;
    end
    else if (inc[2]) begin
      max_value[2] <= maxed_value;
    end
  end
end
always_comb begin
  clear[3] = 1'h0;
  if (((mux_sel > 2'h3) | (~done)) & step) begin
    clear[3] = 1'h1;
  end
end
always_comb begin
  inc[3] = 1'h0;
  if ((5'h3 == 5'h0) & step & (cur_dimensionality > 3'h3)) begin
    inc[3] = 1'h1;
  end
  else if ((mux_sel == 2'h3) & step & (cur_dimensionality > 3'h3)) begin
    inc[3] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[3] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[3] <= 16'h0;
    end
    else if (clear[3]) begin
      dim_counter[3] <= 16'h0;
    end
    else if (inc[3]) begin
      dim_counter[3] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[3] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[3] <= 1'h0;
    end
    else if (clear[3]) begin
      max_value[3] <= 1'h0;
    end
    else if (inc[3]) begin
      max_value[3] <= maxed_value;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    mux_sel_msb_r <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      mux_sel_msb_r <= mux_sel_msb_init;
    end
    else if (restart) begin
      mux_sel_msb_r <= ~mux_sel_msb_r;
    end
  end
end
assign restart = step & (~done);
endmodule   // for_loop_dual_config_4_2_16

module sched_gen_4_16_dual_config_2 (
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic enable,
  input logic enable2,
  input logic finished,
  input logic flush,
  input logic [2:0] mux_sel,
  input logic rst_n,
  input logic [15:0] sched_addr_gen_starting_addr,
  input logic [15:0] sched_addr_gen_starting_addr2,
  input logic [15:0] sched_addr_gen_strides2_0,
  input logic [15:0] sched_addr_gen_strides2_1,
  input logic [15:0] sched_addr_gen_strides_0,
  input logic [15:0] sched_addr_gen_strides_1,
  input logic [15:0] sched_addr_gen_strides_2,
  input logic [15:0] sched_addr_gen_strides_3,
  output logic mux_sel_msb_init,
  output logic valid_output
);

logic [15:0] addr_out;
logic cur_enable;
logic cur_valid_gate;
logic mux_sel_msb_init_w;
logic sched_addr_gen_starting_addr_comp;
logic [3:0][15:0] sched_addr_gen_strides;
logic [1:0][15:0] sched_addr_gen_strides2;
logic [1:0] valid_gate;
logic [1:0] valid_gate_inv;
logic valid_out;
assign cur_valid_gate = valid_gate[mux_sel[2]];
assign valid_gate = ~valid_gate_inv;
assign cur_enable = mux_sel[2] ? enable2: enable;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    valid_gate_inv <= 2'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      valid_gate_inv <= 2'h0;
    end
    else if (finished) begin
      valid_gate_inv[mux_sel[2]] <= 1'h1;
    end
  end
end
always_comb begin
  if (enable & enable2) begin
    mux_sel_msb_init_w = sched_addr_gen_starting_addr_comp;
  end
  else if (enable & (~enable2)) begin
    mux_sel_msb_init_w = 1'h0;
  end
  else if ((~enable) & enable2) begin
    mux_sel_msb_init_w = 1'h1;
  end
  else mux_sel_msb_init_w = 1'h0;
end
assign mux_sel_msb_init = mux_sel_msb_init_w;
always_comb begin
  valid_out = (cycle_count == addr_out) & cur_valid_gate & cur_enable;
end
always_comb begin
  valid_output = valid_out;
end
assign sched_addr_gen_strides2[0] = sched_addr_gen_strides2_0;
assign sched_addr_gen_strides2[1] = sched_addr_gen_strides2_1;
assign sched_addr_gen_strides[0] = sched_addr_gen_strides_0;
assign sched_addr_gen_strides[1] = sched_addr_gen_strides_1;
assign sched_addr_gen_strides[2] = sched_addr_gen_strides_2;
assign sched_addr_gen_strides[3] = sched_addr_gen_strides_3;
addr_gen_4_16_dual_config_2 sched_addr_gen (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(mux_sel),
  .mux_sel_msb_init(mux_sel_msb_init_w),
  .restart(finished),
  .rst_n(rst_n),
  .starting_addr(sched_addr_gen_starting_addr),
  .starting_addr2(sched_addr_gen_starting_addr2),
  .step(valid_out),
  .strides(sched_addr_gen_strides),
  .strides2(sched_addr_gen_strides2),
  .addr_out(addr_out),
  .starting_addr_comp(sched_addr_gen_starting_addr_comp)
);

endmodule   // sched_gen_4_16_dual_config_2

module sram_dp__0 (
  input logic clk,
  input logic clk_en,
  input logic [15:0] data_in_p0,
  input logic flush,
  input logic [4:0] read_addr_p0,
  input logic [4:0] read_addr_p1,
  input logic read_enable_p0,
  input logic read_enable_p1,
  input logic [4:0] write_addr_p0,
  input logic write_enable_p0,
  output logic [15:0] data_out_p0,
  output logic [15:0] data_out_p1
);

logic [15:0] data_array [31:0];

always_ff @(posedge clk) begin
  if (clk_en) begin
    if (write_enable_p0 == 1'h1) begin
      data_array[write_addr_p0] <= data_in_p0;
    end
  end
end
assign data_out_p0 = data_array[read_addr_p0];
always_comb begin
  data_out_p1 = data_array[read_addr_p1];
end
endmodule   // sram_dp__0

module storage_config_seq_1_16_16 (
  input logic clk,
  input logic clk_en,
  input logic [7:0] config_addr_in,
  input logic [15:0] config_data_in,
  input logic config_en,
  input logic config_rd,
  input logic config_wr,
  input logic flush,
  input logic [0:0][0:0] [15:0] rd_data_stg,
  input logic rst_n,
  output logic [4:0] addr_out,
  output logic [0:0] [15:0] rd_data_out,
  output logic ren_out,
  output logic wen_out,
  output logic [0:0] [15:0] wr_data
);

assign addr_out = config_addr_in[4:0];
assign wr_data[0] = config_data_in;
assign rd_data_out[0] = rd_data_stg[0];
assign wen_out = config_wr;
assign ren_out = config_rd;
endmodule   // storage_config_seq_1_16_16

module strg_ub_thin (
  input logic clk,
  input logic clk_en,
  input logic [15:0] data_from_strg,
  input logic [1:0] [16:0] data_in,
  input logic flush,
  input logic [4:0] in2regfile_0_addr_gen_starting_addr,
  input logic [4:0] in2regfile_0_addr_gen_starting_addr2,
  input logic [4:0] in2regfile_0_addr_gen_strides2_0,
  input logic [4:0] in2regfile_0_addr_gen_strides2_1,
  input logic [4:0] in2regfile_0_addr_gen_strides_0,
  input logic [4:0] in2regfile_0_addr_gen_strides_1,
  input logic [4:0] in2regfile_0_addr_gen_strides_2,
  input logic [4:0] in2regfile_0_addr_gen_strides_3,
  input logic [2:0] in2regfile_0_for_loop_dimensionality,
  input logic [1:0] in2regfile_0_for_loop_dimensionality2,
  input logic [15:0] in2regfile_0_for_loop_ranges2_0,
  input logic [15:0] in2regfile_0_for_loop_ranges2_1,
  input logic [15:0] in2regfile_0_for_loop_ranges_0,
  input logic [15:0] in2regfile_0_for_loop_ranges_1,
  input logic [15:0] in2regfile_0_for_loop_ranges_2,
  input logic [15:0] in2regfile_0_for_loop_ranges_3,
  input logic in2regfile_0_sched_gen_enable,
  input logic in2regfile_0_sched_gen_enable2,
  input logic [15:0] in2regfile_0_sched_gen_sched_addr_gen_starting_addr,
  input logic [15:0] in2regfile_0_sched_gen_sched_addr_gen_starting_addr2,
  input logic [15:0] in2regfile_0_sched_gen_sched_addr_gen_strides2_0,
  input logic [15:0] in2regfile_0_sched_gen_sched_addr_gen_strides2_1,
  input logic [15:0] in2regfile_0_sched_gen_sched_addr_gen_strides_0,
  input logic [15:0] in2regfile_0_sched_gen_sched_addr_gen_strides_1,
  input logic [15:0] in2regfile_0_sched_gen_sched_addr_gen_strides_2,
  input logic [15:0] in2regfile_0_sched_gen_sched_addr_gen_strides_3,
  input logic [4:0] regfile2out_0_addr_gen_starting_addr,
  input logic [4:0] regfile2out_0_addr_gen_starting_addr2,
  input logic [4:0] regfile2out_0_addr_gen_strides2_0,
  input logic [4:0] regfile2out_0_addr_gen_strides2_1,
  input logic [4:0] regfile2out_0_addr_gen_strides_0,
  input logic [4:0] regfile2out_0_addr_gen_strides_1,
  input logic [4:0] regfile2out_0_addr_gen_strides_2,
  input logic [4:0] regfile2out_0_addr_gen_strides_3,
  input logic [2:0] regfile2out_0_for_loop_dimensionality,
  input logic [1:0] regfile2out_0_for_loop_dimensionality2,
  input logic [15:0] regfile2out_0_for_loop_ranges2_0,
  input logic [15:0] regfile2out_0_for_loop_ranges2_1,
  input logic [15:0] regfile2out_0_for_loop_ranges_0,
  input logic [15:0] regfile2out_0_for_loop_ranges_1,
  input logic [15:0] regfile2out_0_for_loop_ranges_2,
  input logic [15:0] regfile2out_0_for_loop_ranges_3,
  input logic regfile2out_0_sched_gen_enable,
  input logic regfile2out_0_sched_gen_enable2,
  input logic [15:0] regfile2out_0_sched_gen_sched_addr_gen_starting_addr,
  input logic [15:0] regfile2out_0_sched_gen_sched_addr_gen_starting_addr2,
  input logic [15:0] regfile2out_0_sched_gen_sched_addr_gen_strides2_0,
  input logic [15:0] regfile2out_0_sched_gen_sched_addr_gen_strides2_1,
  input logic [15:0] regfile2out_0_sched_gen_sched_addr_gen_strides_0,
  input logic [15:0] regfile2out_0_sched_gen_sched_addr_gen_strides_1,
  input logic [15:0] regfile2out_0_sched_gen_sched_addr_gen_strides_2,
  input logic [15:0] regfile2out_0_sched_gen_sched_addr_gen_strides_3,
  input logic rst_n,
  output logic [1:0] [16:0] data_out,
  output logic [15:0] data_to_strg,
  output logic [4:0] rd_addr_out,
  output logic ren_to_strg,
  output logic [4:0] tmp0_rdaddr,
  output logic tmp0_rden,
  output logic [1:0] valid_out,
  output logic wen_to_strg,
  output logic [4:0] wr_addr_out
);

logic [15:0] cycle_count;
logic [1:0][15:0] data_in_thin;
logic [1:0][15:0] data_out_int;
logic [1:0][15:0] data_out_int_thin;
logic in2regfile_0_addr_gen_mux_sel_msb_init;
logic [3:0][4:0] in2regfile_0_addr_gen_strides;
logic [1:0][4:0] in2regfile_0_addr_gen_strides2;
logic in2regfile_0_for_loop_mux_sel_msb_init;
logic [2:0] in2regfile_0_for_loop_mux_sel_out;
logic [3:0][15:0] in2regfile_0_for_loop_ranges;
logic [1:0][15:0] in2regfile_0_for_loop_ranges2;
logic in2regfile_0_for_loop_restart;
logic in2regfile_0_sched_gen_mux_sel_msb_init;
logic in2regfile_0_sched_gen_valid_output;
logic read;
logic [4:0] read_addr;
logic read_mux_sel_msb;
logic regfile2out_0_addr_gen_mux_sel_msb_init;
logic [3:0][4:0] regfile2out_0_addr_gen_strides;
logic [1:0][4:0] regfile2out_0_addr_gen_strides2;
logic regfile2out_0_for_loop_mux_sel_msb_init;
logic [2:0] regfile2out_0_for_loop_mux_sel_out;
logic [3:0][15:0] regfile2out_0_for_loop_ranges;
logic [1:0][15:0] regfile2out_0_for_loop_ranges2;
logic regfile2out_0_for_loop_restart;
logic regfile2out_0_sched_gen_mux_sel_msb_init;
logic regfile2out_0_sched_gen_valid_output;
logic [1:0] valid_out_int;
logic write;
logic [4:0] write_addr;
logic write_mux_sel_msb;
assign data_in_thin[0] = data_in[0][15:0];
assign data_in_thin[1] = data_in[1][15:0];

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    cycle_count <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      cycle_count <= 16'h0;
    end
    else cycle_count <= cycle_count + 16'h1;
  end
end
assign valid_out_int[0] = read & (~read_mux_sel_msb);
assign valid_out_int[1] = read & read_mux_sel_msb;
assign data_out_int_thin = data_out_int;
assign data_out[0][15:0] = data_out_int_thin[0];
assign data_out[0][16] = 1'h0;
assign data_out[1][15:0] = data_out_int_thin[1];
assign data_out[1][16] = 1'h0;
assign valid_out = valid_out_int;
assign write = in2regfile_0_sched_gen_valid_output;
assign in2regfile_0_for_loop_mux_sel_msb_init = in2regfile_0_sched_gen_mux_sel_msb_init;
assign in2regfile_0_addr_gen_mux_sel_msb_init = in2regfile_0_sched_gen_mux_sel_msb_init;
assign write_mux_sel_msb = in2regfile_0_for_loop_mux_sel_out[2];
assign read = regfile2out_0_sched_gen_valid_output;
assign regfile2out_0_for_loop_mux_sel_msb_init = regfile2out_0_sched_gen_mux_sel_msb_init;
assign regfile2out_0_addr_gen_mux_sel_msb_init = regfile2out_0_sched_gen_mux_sel_msb_init;
assign read_mux_sel_msb = regfile2out_0_for_loop_mux_sel_out[2];
assign wen_to_strg = |write;
assign ren_to_strg = |read;
assign data_out_int[0] = data_from_strg;
assign data_out_int[1] = data_from_strg;
assign wr_addr_out = write_addr[4:0];
assign data_to_strg = data_in_thin[write_mux_sel_msb];
assign rd_addr_out = read_addr[4:0];
assign tmp0_rdaddr = 5'h0;
assign tmp0_rden = 1'h0;
assign in2regfile_0_for_loop_ranges[0] = in2regfile_0_for_loop_ranges_0;
assign in2regfile_0_for_loop_ranges[1] = in2regfile_0_for_loop_ranges_1;
assign in2regfile_0_for_loop_ranges[2] = in2regfile_0_for_loop_ranges_2;
assign in2regfile_0_for_loop_ranges[3] = in2regfile_0_for_loop_ranges_3;
assign in2regfile_0_for_loop_ranges2[0] = in2regfile_0_for_loop_ranges2_0;
assign in2regfile_0_for_loop_ranges2[1] = in2regfile_0_for_loop_ranges2_1;
assign in2regfile_0_addr_gen_strides2[0] = in2regfile_0_addr_gen_strides2_0;
assign in2regfile_0_addr_gen_strides2[1] = in2regfile_0_addr_gen_strides2_1;
assign in2regfile_0_addr_gen_strides[0] = in2regfile_0_addr_gen_strides_0;
assign in2regfile_0_addr_gen_strides[1] = in2regfile_0_addr_gen_strides_1;
assign in2regfile_0_addr_gen_strides[2] = in2regfile_0_addr_gen_strides_2;
assign in2regfile_0_addr_gen_strides[3] = in2regfile_0_addr_gen_strides_3;
assign regfile2out_0_for_loop_ranges[0] = regfile2out_0_for_loop_ranges_0;
assign regfile2out_0_for_loop_ranges[1] = regfile2out_0_for_loop_ranges_1;
assign regfile2out_0_for_loop_ranges[2] = regfile2out_0_for_loop_ranges_2;
assign regfile2out_0_for_loop_ranges[3] = regfile2out_0_for_loop_ranges_3;
assign regfile2out_0_for_loop_ranges2[0] = regfile2out_0_for_loop_ranges2_0;
assign regfile2out_0_for_loop_ranges2[1] = regfile2out_0_for_loop_ranges2_1;
assign regfile2out_0_addr_gen_strides2[0] = regfile2out_0_addr_gen_strides2_0;
assign regfile2out_0_addr_gen_strides2[1] = regfile2out_0_addr_gen_strides2_1;
assign regfile2out_0_addr_gen_strides[0] = regfile2out_0_addr_gen_strides_0;
assign regfile2out_0_addr_gen_strides[1] = regfile2out_0_addr_gen_strides_1;
assign regfile2out_0_addr_gen_strides[2] = regfile2out_0_addr_gen_strides_2;
assign regfile2out_0_addr_gen_strides[3] = regfile2out_0_addr_gen_strides_3;
for_loop_dual_config_4_2_16 in2regfile_0_for_loop (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(in2regfile_0_for_loop_dimensionality),
  .dimensionality2(in2regfile_0_for_loop_dimensionality2),
  .flush(flush),
  .mux_sel_msb_init(in2regfile_0_for_loop_mux_sel_msb_init),
  .ranges(in2regfile_0_for_loop_ranges),
  .ranges2(in2regfile_0_for_loop_ranges2),
  .rst_n(rst_n),
  .step(write),
  .mux_sel_out(in2regfile_0_for_loop_mux_sel_out),
  .restart(in2regfile_0_for_loop_restart)
);

addr_gen_4_5_dual_config_2 in2regfile_0_addr_gen (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(in2regfile_0_for_loop_mux_sel_out),
  .mux_sel_msb_init(in2regfile_0_addr_gen_mux_sel_msb_init),
  .restart(in2regfile_0_for_loop_restart),
  .rst_n(rst_n),
  .starting_addr(in2regfile_0_addr_gen_starting_addr),
  .starting_addr2(in2regfile_0_addr_gen_starting_addr2),
  .step(write),
  .strides(in2regfile_0_addr_gen_strides),
  .strides2(in2regfile_0_addr_gen_strides2),
  .addr_out(write_addr)
);

sched_gen_4_16_dual_config_2 in2regfile_0_sched_gen (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(in2regfile_0_sched_gen_enable),
  .enable2(in2regfile_0_sched_gen_enable2),
  .finished(in2regfile_0_for_loop_restart),
  .flush(flush),
  .mux_sel(in2regfile_0_for_loop_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(in2regfile_0_sched_gen_sched_addr_gen_starting_addr),
  .sched_addr_gen_starting_addr2(in2regfile_0_sched_gen_sched_addr_gen_starting_addr2),
  .sched_addr_gen_strides2_0(in2regfile_0_sched_gen_sched_addr_gen_strides2_0),
  .sched_addr_gen_strides2_1(in2regfile_0_sched_gen_sched_addr_gen_strides2_1),
  .sched_addr_gen_strides_0(in2regfile_0_sched_gen_sched_addr_gen_strides_0),
  .sched_addr_gen_strides_1(in2regfile_0_sched_gen_sched_addr_gen_strides_1),
  .sched_addr_gen_strides_2(in2regfile_0_sched_gen_sched_addr_gen_strides_2),
  .sched_addr_gen_strides_3(in2regfile_0_sched_gen_sched_addr_gen_strides_3),
  .mux_sel_msb_init(in2regfile_0_sched_gen_mux_sel_msb_init),
  .valid_output(in2regfile_0_sched_gen_valid_output)
);

for_loop_dual_config_4_2_16 regfile2out_0_for_loop (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(regfile2out_0_for_loop_dimensionality),
  .dimensionality2(regfile2out_0_for_loop_dimensionality2),
  .flush(flush),
  .mux_sel_msb_init(regfile2out_0_for_loop_mux_sel_msb_init),
  .ranges(regfile2out_0_for_loop_ranges),
  .ranges2(regfile2out_0_for_loop_ranges2),
  .rst_n(rst_n),
  .step(read),
  .mux_sel_out(regfile2out_0_for_loop_mux_sel_out),
  .restart(regfile2out_0_for_loop_restart)
);

addr_gen_4_5_dual_config_2 regfile2out_0_addr_gen (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(regfile2out_0_for_loop_mux_sel_out),
  .mux_sel_msb_init(regfile2out_0_addr_gen_mux_sel_msb_init),
  .restart(regfile2out_0_for_loop_restart),
  .rst_n(rst_n),
  .starting_addr(regfile2out_0_addr_gen_starting_addr),
  .starting_addr2(regfile2out_0_addr_gen_starting_addr2),
  .step(read),
  .strides(regfile2out_0_addr_gen_strides),
  .strides2(regfile2out_0_addr_gen_strides2),
  .addr_out(read_addr)
);

sched_gen_4_16_dual_config_2 regfile2out_0_sched_gen (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(regfile2out_0_sched_gen_enable),
  .enable2(regfile2out_0_sched_gen_enable2),
  .finished(regfile2out_0_for_loop_restart),
  .flush(flush),
  .mux_sel(regfile2out_0_for_loop_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(regfile2out_0_sched_gen_sched_addr_gen_starting_addr),
  .sched_addr_gen_starting_addr2(regfile2out_0_sched_gen_sched_addr_gen_starting_addr2),
  .sched_addr_gen_strides2_0(regfile2out_0_sched_gen_sched_addr_gen_strides2_0),
  .sched_addr_gen_strides2_1(regfile2out_0_sched_gen_sched_addr_gen_strides2_1),
  .sched_addr_gen_strides_0(regfile2out_0_sched_gen_sched_addr_gen_strides_0),
  .sched_addr_gen_strides_1(regfile2out_0_sched_gen_sched_addr_gen_strides_1),
  .sched_addr_gen_strides_2(regfile2out_0_sched_gen_sched_addr_gen_strides_2),
  .sched_addr_gen_strides_3(regfile2out_0_sched_gen_sched_addr_gen_strides_3),
  .mux_sel_msb_init(regfile2out_0_sched_gen_mux_sel_msb_init),
  .valid_output(regfile2out_0_sched_gen_valid_output)
);

endmodule   // strg_ub_thin

module strg_ub_thin_flat (
  input logic clk,
  input logic clk_en,
  input logic [0:0] [16:0] data_in_f_0,
  input logic [0:0] [16:0] data_in_f_1,
  input logic flush,
  input logic rst_n,
  input logic [15:0] strg_ub_thin_inst_data_from_strg_lifted,
  input logic [4:0] strg_ub_thin_inst_in2regfile_0_addr_gen_starting_addr,
  input logic [4:0] strg_ub_thin_inst_in2regfile_0_addr_gen_starting_addr2,
  input logic [4:0] strg_ub_thin_inst_in2regfile_0_addr_gen_strides2_0,
  input logic [4:0] strg_ub_thin_inst_in2regfile_0_addr_gen_strides2_1,
  input logic [4:0] strg_ub_thin_inst_in2regfile_0_addr_gen_strides_0,
  input logic [4:0] strg_ub_thin_inst_in2regfile_0_addr_gen_strides_1,
  input logic [4:0] strg_ub_thin_inst_in2regfile_0_addr_gen_strides_2,
  input logic [4:0] strg_ub_thin_inst_in2regfile_0_addr_gen_strides_3,
  input logic [2:0] strg_ub_thin_inst_in2regfile_0_for_loop_dimensionality,
  input logic [1:0] strg_ub_thin_inst_in2regfile_0_for_loop_dimensionality2,
  input logic [15:0] strg_ub_thin_inst_in2regfile_0_for_loop_ranges2_0,
  input logic [15:0] strg_ub_thin_inst_in2regfile_0_for_loop_ranges2_1,
  input logic [15:0] strg_ub_thin_inst_in2regfile_0_for_loop_ranges_0,
  input logic [15:0] strg_ub_thin_inst_in2regfile_0_for_loop_ranges_1,
  input logic [15:0] strg_ub_thin_inst_in2regfile_0_for_loop_ranges_2,
  input logic [15:0] strg_ub_thin_inst_in2regfile_0_for_loop_ranges_3,
  input logic strg_ub_thin_inst_in2regfile_0_sched_gen_enable,
  input logic strg_ub_thin_inst_in2regfile_0_sched_gen_enable2,
  input logic [15:0] strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr,
  input logic [15:0] strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr2,
  input logic [15:0] strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_0,
  input logic [15:0] strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_1,
  input logic [15:0] strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_0,
  input logic [15:0] strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_1,
  input logic [15:0] strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_2,
  input logic [15:0] strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_3,
  input logic [4:0] strg_ub_thin_inst_regfile2out_0_addr_gen_starting_addr,
  input logic [4:0] strg_ub_thin_inst_regfile2out_0_addr_gen_starting_addr2,
  input logic [4:0] strg_ub_thin_inst_regfile2out_0_addr_gen_strides2_0,
  input logic [4:0] strg_ub_thin_inst_regfile2out_0_addr_gen_strides2_1,
  input logic [4:0] strg_ub_thin_inst_regfile2out_0_addr_gen_strides_0,
  input logic [4:0] strg_ub_thin_inst_regfile2out_0_addr_gen_strides_1,
  input logic [4:0] strg_ub_thin_inst_regfile2out_0_addr_gen_strides_2,
  input logic [4:0] strg_ub_thin_inst_regfile2out_0_addr_gen_strides_3,
  input logic [2:0] strg_ub_thin_inst_regfile2out_0_for_loop_dimensionality,
  input logic [1:0] strg_ub_thin_inst_regfile2out_0_for_loop_dimensionality2,
  input logic [15:0] strg_ub_thin_inst_regfile2out_0_for_loop_ranges2_0,
  input logic [15:0] strg_ub_thin_inst_regfile2out_0_for_loop_ranges2_1,
  input logic [15:0] strg_ub_thin_inst_regfile2out_0_for_loop_ranges_0,
  input logic [15:0] strg_ub_thin_inst_regfile2out_0_for_loop_ranges_1,
  input logic [15:0] strg_ub_thin_inst_regfile2out_0_for_loop_ranges_2,
  input logic [15:0] strg_ub_thin_inst_regfile2out_0_for_loop_ranges_3,
  input logic strg_ub_thin_inst_regfile2out_0_sched_gen_enable,
  input logic strg_ub_thin_inst_regfile2out_0_sched_gen_enable2,
  input logic [15:0] strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr,
  input logic [15:0] strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr2,
  input logic [15:0] strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_0,
  input logic [15:0] strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_1,
  input logic [15:0] strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_0,
  input logic [15:0] strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_1,
  input logic [15:0] strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_2,
  input logic [15:0] strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_3,
  output logic [0:0] [16:0] data_out_f_0,
  output logic [0:0] [16:0] data_out_f_1,
  output logic [15:0] strg_ub_thin_inst_data_to_strg_lifted,
  output logic [4:0] strg_ub_thin_inst_rd_addr_out_lifted,
  output logic strg_ub_thin_inst_ren_to_strg_lifted,
  output logic [4:0] strg_ub_thin_inst_tmp0_rdaddr_lifted,
  output logic strg_ub_thin_inst_tmp0_rden_lifted,
  output logic strg_ub_thin_inst_wen_to_strg_lifted,
  output logic [4:0] strg_ub_thin_inst_wr_addr_out_lifted,
  output logic valid_out_f_b_0,
  output logic valid_out_f_b_1
);

logic [1:0][16:0] strg_ub_thin_inst_data_in;
logic [1:0][16:0] strg_ub_thin_inst_data_out;
logic [1:0] strg_ub_thin_inst_valid_out;
assign strg_ub_thin_inst_data_in[0] = data_in_f_0;
assign strg_ub_thin_inst_data_in[1] = data_in_f_1;
assign valid_out_f_b_0 = strg_ub_thin_inst_valid_out[0];
assign valid_out_f_b_1 = strg_ub_thin_inst_valid_out[1];
assign data_out_f_0 = strg_ub_thin_inst_data_out[0];
assign data_out_f_1 = strg_ub_thin_inst_data_out[1];
strg_ub_thin strg_ub_thin_inst (
  .clk(clk),
  .clk_en(clk_en),
  .data_from_strg(strg_ub_thin_inst_data_from_strg_lifted),
  .data_in(strg_ub_thin_inst_data_in),
  .flush(flush),
  .in2regfile_0_addr_gen_starting_addr(strg_ub_thin_inst_in2regfile_0_addr_gen_starting_addr),
  .in2regfile_0_addr_gen_starting_addr2(strg_ub_thin_inst_in2regfile_0_addr_gen_starting_addr2),
  .in2regfile_0_addr_gen_strides2_0(strg_ub_thin_inst_in2regfile_0_addr_gen_strides2_0),
  .in2regfile_0_addr_gen_strides2_1(strg_ub_thin_inst_in2regfile_0_addr_gen_strides2_1),
  .in2regfile_0_addr_gen_strides_0(strg_ub_thin_inst_in2regfile_0_addr_gen_strides_0),
  .in2regfile_0_addr_gen_strides_1(strg_ub_thin_inst_in2regfile_0_addr_gen_strides_1),
  .in2regfile_0_addr_gen_strides_2(strg_ub_thin_inst_in2regfile_0_addr_gen_strides_2),
  .in2regfile_0_addr_gen_strides_3(strg_ub_thin_inst_in2regfile_0_addr_gen_strides_3),
  .in2regfile_0_for_loop_dimensionality(strg_ub_thin_inst_in2regfile_0_for_loop_dimensionality),
  .in2regfile_0_for_loop_dimensionality2(strg_ub_thin_inst_in2regfile_0_for_loop_dimensionality2),
  .in2regfile_0_for_loop_ranges2_0(strg_ub_thin_inst_in2regfile_0_for_loop_ranges2_0),
  .in2regfile_0_for_loop_ranges2_1(strg_ub_thin_inst_in2regfile_0_for_loop_ranges2_1),
  .in2regfile_0_for_loop_ranges_0(strg_ub_thin_inst_in2regfile_0_for_loop_ranges_0),
  .in2regfile_0_for_loop_ranges_1(strg_ub_thin_inst_in2regfile_0_for_loop_ranges_1),
  .in2regfile_0_for_loop_ranges_2(strg_ub_thin_inst_in2regfile_0_for_loop_ranges_2),
  .in2regfile_0_for_loop_ranges_3(strg_ub_thin_inst_in2regfile_0_for_loop_ranges_3),
  .in2regfile_0_sched_gen_enable(strg_ub_thin_inst_in2regfile_0_sched_gen_enable),
  .in2regfile_0_sched_gen_enable2(strg_ub_thin_inst_in2regfile_0_sched_gen_enable2),
  .in2regfile_0_sched_gen_sched_addr_gen_starting_addr(strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr),
  .in2regfile_0_sched_gen_sched_addr_gen_starting_addr2(strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_starting_addr2),
  .in2regfile_0_sched_gen_sched_addr_gen_strides2_0(strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_0),
  .in2regfile_0_sched_gen_sched_addr_gen_strides2_1(strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides2_1),
  .in2regfile_0_sched_gen_sched_addr_gen_strides_0(strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_0),
  .in2regfile_0_sched_gen_sched_addr_gen_strides_1(strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_1),
  .in2regfile_0_sched_gen_sched_addr_gen_strides_2(strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_2),
  .in2regfile_0_sched_gen_sched_addr_gen_strides_3(strg_ub_thin_inst_in2regfile_0_sched_gen_sched_addr_gen_strides_3),
  .regfile2out_0_addr_gen_starting_addr(strg_ub_thin_inst_regfile2out_0_addr_gen_starting_addr),
  .regfile2out_0_addr_gen_starting_addr2(strg_ub_thin_inst_regfile2out_0_addr_gen_starting_addr2),
  .regfile2out_0_addr_gen_strides2_0(strg_ub_thin_inst_regfile2out_0_addr_gen_strides2_0),
  .regfile2out_0_addr_gen_strides2_1(strg_ub_thin_inst_regfile2out_0_addr_gen_strides2_1),
  .regfile2out_0_addr_gen_strides_0(strg_ub_thin_inst_regfile2out_0_addr_gen_strides_0),
  .regfile2out_0_addr_gen_strides_1(strg_ub_thin_inst_regfile2out_0_addr_gen_strides_1),
  .regfile2out_0_addr_gen_strides_2(strg_ub_thin_inst_regfile2out_0_addr_gen_strides_2),
  .regfile2out_0_addr_gen_strides_3(strg_ub_thin_inst_regfile2out_0_addr_gen_strides_3),
  .regfile2out_0_for_loop_dimensionality(strg_ub_thin_inst_regfile2out_0_for_loop_dimensionality),
  .regfile2out_0_for_loop_dimensionality2(strg_ub_thin_inst_regfile2out_0_for_loop_dimensionality2),
  .regfile2out_0_for_loop_ranges2_0(strg_ub_thin_inst_regfile2out_0_for_loop_ranges2_0),
  .regfile2out_0_for_loop_ranges2_1(strg_ub_thin_inst_regfile2out_0_for_loop_ranges2_1),
  .regfile2out_0_for_loop_ranges_0(strg_ub_thin_inst_regfile2out_0_for_loop_ranges_0),
  .regfile2out_0_for_loop_ranges_1(strg_ub_thin_inst_regfile2out_0_for_loop_ranges_1),
  .regfile2out_0_for_loop_ranges_2(strg_ub_thin_inst_regfile2out_0_for_loop_ranges_2),
  .regfile2out_0_for_loop_ranges_3(strg_ub_thin_inst_regfile2out_0_for_loop_ranges_3),
  .regfile2out_0_sched_gen_enable(strg_ub_thin_inst_regfile2out_0_sched_gen_enable),
  .regfile2out_0_sched_gen_enable2(strg_ub_thin_inst_regfile2out_0_sched_gen_enable2),
  .regfile2out_0_sched_gen_sched_addr_gen_starting_addr(strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr),
  .regfile2out_0_sched_gen_sched_addr_gen_starting_addr2(strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_starting_addr2),
  .regfile2out_0_sched_gen_sched_addr_gen_strides2_0(strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_0),
  .regfile2out_0_sched_gen_sched_addr_gen_strides2_1(strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides2_1),
  .regfile2out_0_sched_gen_sched_addr_gen_strides_0(strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_0),
  .regfile2out_0_sched_gen_sched_addr_gen_strides_1(strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_1),
  .regfile2out_0_sched_gen_sched_addr_gen_strides_2(strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_2),
  .regfile2out_0_sched_gen_sched_addr_gen_strides_3(strg_ub_thin_inst_regfile2out_0_sched_gen_sched_addr_gen_strides_3),
  .rst_n(rst_n),
  .data_out(strg_ub_thin_inst_data_out),
  .data_to_strg(strg_ub_thin_inst_data_to_strg_lifted),
  .rd_addr_out(strg_ub_thin_inst_rd_addr_out_lifted),
  .ren_to_strg(strg_ub_thin_inst_ren_to_strg_lifted),
  .tmp0_rdaddr(strg_ub_thin_inst_tmp0_rdaddr_lifted),
  .tmp0_rden(strg_ub_thin_inst_tmp0_rden_lifted),
  .valid_out(strg_ub_thin_inst_valid_out),
  .wen_to_strg(strg_ub_thin_inst_wen_to_strg_lifted),
  .wr_addr_out(strg_ub_thin_inst_wr_addr_out_lifted)
);

endmodule   // strg_ub_thin_flat


module PE_inner (
  input logic [31:0] CONFIG_SPACE_0,
  input logic [31:0] CONFIG_SPACE_1,
  input logic [21:0] CONFIG_SPACE_2,
  input logic [0:0] [16:0] PE_input_width_17_num_0,
  input logic PE_input_width_17_num_0_dense,
  input logic PE_input_width_17_num_0_valid,
  input logic [0:0] [16:0] PE_input_width_17_num_1,
  input logic PE_input_width_17_num_1_dense,
  input logic PE_input_width_17_num_1_valid,
  input logic [0:0] [16:0] PE_input_width_17_num_2,
  input logic PE_input_width_17_num_2_valid,
  input logic [0:0] [16:0] PE_input_width_17_num_3,
  input logic PE_input_width_17_num_3_valid,
  input logic PE_input_width_1_num_0,
  input logic PE_input_width_1_num_1,
  input logic PE_input_width_1_num_2,
  input logic PE_output_width_17_num_0_dense,
  input logic PE_output_width_17_num_0_ready,
  input logic PE_output_width_17_num_1_ready,
  input logic PE_output_width_17_num_2_ready,
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [2:0] mode,
  input logic rst_n,
  input logic tile_en,
  output logic PE_input_width_17_num_0_ready,
  output logic PE_input_width_17_num_1_ready,
  output logic PE_input_width_17_num_2_ready,
  output logic PE_input_width_17_num_3_ready,
  output logic [15:0] PE_onyx_inst_onyxpeintf_O2,
  output logic [15:0] PE_onyx_inst_onyxpeintf_O3,
  output logic [15:0] PE_onyx_inst_onyxpeintf_O4,
  output logic [0:0] [16:0] PE_output_width_17_num_0,
  output logic PE_output_width_17_num_0_valid,
  output logic [0:0] [16:0] PE_output_width_17_num_1,
  output logic PE_output_width_17_num_1_valid,
  output logic [0:0] [16:0] PE_output_width_17_num_2,
  output logic PE_output_width_17_num_2_valid,
  output logic PE_output_width_1_num_0
);

logic [85:0] CONFIG_SPACE;
logic gclk;
logic [0:0][16:0] input_width_17_num_0_fifo_out;
logic input_width_17_num_0_fifo_out_ready;
logic input_width_17_num_0_fifo_out_valid;
logic input_width_17_num_0_input_fifo_empty;
logic input_width_17_num_0_input_fifo_full;
logic [0:0][16:0] input_width_17_num_1_fifo_out;
logic input_width_17_num_1_fifo_out_ready;
logic input_width_17_num_1_fifo_out_valid;
logic input_width_17_num_1_input_fifo_empty;
logic input_width_17_num_1_input_fifo_full;
logic [0:0][16:0] input_width_17_num_2_fifo_out;
logic input_width_17_num_2_fifo_out_ready;
logic input_width_17_num_2_fifo_out_valid;
logic input_width_17_num_2_input_fifo_empty;
logic input_width_17_num_2_input_fifo_full;
logic [0:0][16:0] input_width_17_num_3_fifo_out;
logic input_width_17_num_3_fifo_out_ready;
logic input_width_17_num_3_fifo_out_valid;
logic input_width_17_num_3_input_fifo_empty;
logic input_width_17_num_3_input_fifo_full;
logic mem_ctrl_PE_onyx_flat_PE_onyx_inst_dense_mode;
logic [83:0] mem_ctrl_PE_onyx_flat_PE_onyx_inst_onyxpeintf_inst;
logic mem_ctrl_PE_onyx_flat_PE_onyx_inst_tile_en;
logic mem_ctrl_PE_onyx_flat_clk;
logic [0:0][16:0] mem_ctrl_PE_onyx_flat_data0_f_;
logic mem_ctrl_PE_onyx_flat_data0_ready_f_;
logic mem_ctrl_PE_onyx_flat_data0_valid_f_;
logic [0:0][16:0] mem_ctrl_PE_onyx_flat_data1_f_;
logic mem_ctrl_PE_onyx_flat_data1_ready_f_;
logic mem_ctrl_PE_onyx_flat_data1_valid_f_;
logic [0:0][16:0] mem_ctrl_PE_onyx_flat_res_f_;
logic mem_ctrl_PE_onyx_flat_res_p_f_;
logic mem_ctrl_PE_onyx_flat_res_ready_f_;
logic mem_ctrl_PE_onyx_flat_res_valid_f_;
logic [15:0] mem_ctrl_RepeatSignalGenerator_flat_RepeatSignalGenerator_inst_stop_lvl;
logic mem_ctrl_RepeatSignalGenerator_flat_RepeatSignalGenerator_inst_tile_en;
logic mem_ctrl_RepeatSignalGenerator_flat_base_data_in_ready_f_;
logic mem_ctrl_RepeatSignalGenerator_flat_clk;
logic [0:0][16:0] mem_ctrl_RepeatSignalGenerator_flat_repsig_data_out_f_;
logic mem_ctrl_RepeatSignalGenerator_flat_repsig_data_out_valid_f_;
logic mem_ctrl_Repeat_flat_Repeat_inst_root;
logic mem_ctrl_Repeat_flat_Repeat_inst_spacc_mode;
logic [15:0] mem_ctrl_Repeat_flat_Repeat_inst_stop_lvl;
logic mem_ctrl_Repeat_flat_Repeat_inst_tile_en;
logic mem_ctrl_Repeat_flat_clk;
logic mem_ctrl_Repeat_flat_proc_data_in_ready_f_;
logic [0:0][16:0] mem_ctrl_Repeat_flat_ref_data_out_f_;
logic mem_ctrl_Repeat_flat_ref_data_out_valid_f_;
logic mem_ctrl_Repeat_flat_repsig_data_in_ready_f_;
logic mem_ctrl_crddrop_flat_clk;
logic mem_ctrl_crddrop_flat_cmrg_coord_in_0_ready_f_;
logic mem_ctrl_crddrop_flat_cmrg_coord_in_1_ready_f_;
logic [0:0][16:0] mem_ctrl_crddrop_flat_cmrg_coord_out_0_f_;
logic mem_ctrl_crddrop_flat_cmrg_coord_out_0_valid_f_;
logic [0:0][16:0] mem_ctrl_crddrop_flat_cmrg_coord_out_1_f_;
logic mem_ctrl_crddrop_flat_cmrg_coord_out_1_valid_f_;
logic mem_ctrl_crddrop_flat_crddrop_inst_cmrg_enable;
logic [15:0] mem_ctrl_crddrop_flat_crddrop_inst_cmrg_stop_lvl;
logic mem_ctrl_crddrop_flat_crddrop_inst_tile_en;
logic mem_ctrl_crdhold_flat_clk;
logic mem_ctrl_crdhold_flat_cmrg_coord_in_0_ready_f_;
logic mem_ctrl_crdhold_flat_cmrg_coord_in_1_ready_f_;
logic [0:0][16:0] mem_ctrl_crdhold_flat_cmrg_coord_out_0_f_;
logic mem_ctrl_crdhold_flat_cmrg_coord_out_0_valid_f_;
logic [0:0][16:0] mem_ctrl_crdhold_flat_cmrg_coord_out_1_f_;
logic mem_ctrl_crdhold_flat_cmrg_coord_out_1_valid_f_;
logic mem_ctrl_crdhold_flat_crdhold_inst_cmrg_enable;
logic [15:0] mem_ctrl_crdhold_flat_crdhold_inst_cmrg_stop_lvl;
logic mem_ctrl_crdhold_flat_crdhold_inst_tile_en;
logic mem_ctrl_intersect_unit_flat_clk;
logic mem_ctrl_intersect_unit_flat_coord_in_0_ready_f_;
logic mem_ctrl_intersect_unit_flat_coord_in_1_ready_f_;
logic [0:0][16:0] mem_ctrl_intersect_unit_flat_coord_out_f_;
logic mem_ctrl_intersect_unit_flat_coord_out_valid_f_;
logic mem_ctrl_intersect_unit_flat_intersect_unit_inst_joiner_op;
logic mem_ctrl_intersect_unit_flat_intersect_unit_inst_tile_en;
logic mem_ctrl_intersect_unit_flat_pos_in_0_ready_f_;
logic mem_ctrl_intersect_unit_flat_pos_in_1_ready_f_;
logic [0:0][16:0] mem_ctrl_intersect_unit_flat_pos_out_0_f_;
logic mem_ctrl_intersect_unit_flat_pos_out_0_valid_f_;
logic [0:0][16:0] mem_ctrl_intersect_unit_flat_pos_out_1_f_;
logic mem_ctrl_intersect_unit_flat_pos_out_1_valid_f_;
logic mem_ctrl_reg_cr_flat_clk;
logic mem_ctrl_reg_cr_flat_data_in_ready_f_;
logic [0:0][16:0] mem_ctrl_reg_cr_flat_data_out_f_;
logic mem_ctrl_reg_cr_flat_data_out_valid_f_;
logic [15:0] mem_ctrl_reg_cr_flat_reg_cr_inst_default_value;
logic [15:0] mem_ctrl_reg_cr_flat_reg_cr_inst_stop_lvl;
logic mem_ctrl_reg_cr_flat_reg_cr_inst_tile_en;
logic [0:0][16:0] output_width_17_num_0_fifo_in;
logic output_width_17_num_0_fifo_in_ready;
logic output_width_17_num_0_fifo_in_valid;
logic [0:0][16:0] output_width_17_num_0_output_fifo_data_out;
logic output_width_17_num_0_output_fifo_empty;
logic output_width_17_num_0_output_fifo_full;
logic [0:0][16:0] output_width_17_num_1_fifo_in;
logic output_width_17_num_1_fifo_in_ready;
logic output_width_17_num_1_fifo_in_valid;
logic [0:0][16:0] output_width_17_num_1_output_fifo_data_out;
logic output_width_17_num_1_output_fifo_empty;
logic output_width_17_num_1_output_fifo_full;
logic [0:0][16:0] output_width_17_num_2_fifo_in;
logic output_width_17_num_2_fifo_in_ready;
logic output_width_17_num_2_fifo_in_valid;
logic [0:0][16:0] output_width_17_num_2_output_fifo_data_out;
logic output_width_17_num_2_output_fifo_empty;
logic output_width_17_num_2_output_fifo_full;
assign gclk = clk & tile_en;
assign mem_ctrl_intersect_unit_flat_clk = gclk & (mode == 3'h0);
assign mem_ctrl_crddrop_flat_clk = gclk & (mode == 3'h1);
assign mem_ctrl_crdhold_flat_clk = gclk & (mode == 3'h2);
assign mem_ctrl_PE_onyx_flat_clk = gclk & (mode == 3'h3);
assign mem_ctrl_Repeat_flat_clk = gclk & (mode == 3'h4);
assign mem_ctrl_RepeatSignalGenerator_flat_clk = gclk & (mode == 3'h5);
assign mem_ctrl_reg_cr_flat_clk = gclk & (mode == 3'h6);
assign input_width_17_num_0_fifo_out_valid = ~input_width_17_num_0_input_fifo_empty;
always_comb begin
  input_width_17_num_0_fifo_out_ready = 1'h1;
  if (mode == 3'h0) begin
    input_width_17_num_0_fifo_out_ready = mem_ctrl_intersect_unit_flat_coord_in_0_ready_f_;
  end
  else if (mode == 3'h1) begin
    input_width_17_num_0_fifo_out_ready = mem_ctrl_crddrop_flat_cmrg_coord_in_0_ready_f_;
  end
  else if (mode == 3'h2) begin
    input_width_17_num_0_fifo_out_ready = mem_ctrl_crdhold_flat_cmrg_coord_in_0_ready_f_;
  end
  else if (mode == 3'h3) begin
    input_width_17_num_0_fifo_out_ready = mem_ctrl_PE_onyx_flat_data0_ready_f_;
  end
  else if (mode == 3'h4) begin
    input_width_17_num_0_fifo_out_ready = mem_ctrl_Repeat_flat_proc_data_in_ready_f_;
  end
  else if (mode == 3'h5) begin
    input_width_17_num_0_fifo_out_ready = mem_ctrl_RepeatSignalGenerator_flat_base_data_in_ready_f_;
  end
  else if (mode == 3'h6) begin
    input_width_17_num_0_fifo_out_ready = mem_ctrl_reg_cr_flat_data_in_ready_f_;
  end
end
assign mem_ctrl_PE_onyx_flat_data0_f_ = PE_input_width_17_num_0_dense ? PE_input_width_17_num_0:
    input_width_17_num_0_fifo_out;
assign mem_ctrl_PE_onyx_flat_data0_valid_f_ = PE_input_width_17_num_0_dense ? 1'h1: input_width_17_num_0_fifo_out_valid;
always_comb begin
  PE_input_width_17_num_0_ready = 1'h1;
  if (mode == 3'h0) begin
    PE_input_width_17_num_0_ready = ~input_width_17_num_0_input_fifo_full;
  end
  else if (mode == 3'h1) begin
    PE_input_width_17_num_0_ready = ~input_width_17_num_0_input_fifo_full;
  end
  else if (mode == 3'h2) begin
    PE_input_width_17_num_0_ready = ~input_width_17_num_0_input_fifo_full;
  end
  else if (mode == 3'h3) begin
    PE_input_width_17_num_0_ready = PE_input_width_17_num_0_dense ? 1'h1: ~input_width_17_num_0_input_fifo_full;
  end
  else if (mode == 3'h4) begin
    PE_input_width_17_num_0_ready = ~input_width_17_num_0_input_fifo_full;
  end
  else if (mode == 3'h5) begin
    PE_input_width_17_num_0_ready = ~input_width_17_num_0_input_fifo_full;
  end
  else if (mode == 3'h6) begin
    PE_input_width_17_num_0_ready = ~input_width_17_num_0_input_fifo_full;
  end
end
assign input_width_17_num_1_fifo_out_valid = ~input_width_17_num_1_input_fifo_empty;
always_comb begin
  input_width_17_num_1_fifo_out_ready = 1'h1;
  if (mode == 3'h0) begin
    input_width_17_num_1_fifo_out_ready = mem_ctrl_intersect_unit_flat_coord_in_1_ready_f_;
  end
  else if (mode == 3'h1) begin
    input_width_17_num_1_fifo_out_ready = mem_ctrl_crddrop_flat_cmrg_coord_in_1_ready_f_;
  end
  else if (mode == 3'h2) begin
    input_width_17_num_1_fifo_out_ready = mem_ctrl_crdhold_flat_cmrg_coord_in_1_ready_f_;
  end
  else if (mode == 3'h3) begin
    input_width_17_num_1_fifo_out_ready = mem_ctrl_PE_onyx_flat_data1_ready_f_;
  end
  else if (mode == 3'h4) begin
    input_width_17_num_1_fifo_out_ready = mem_ctrl_Repeat_flat_repsig_data_in_ready_f_;
  end
end
assign mem_ctrl_PE_onyx_flat_data1_f_ = PE_input_width_17_num_1_dense ? PE_input_width_17_num_1:
    input_width_17_num_1_fifo_out;
assign mem_ctrl_PE_onyx_flat_data1_valid_f_ = PE_input_width_17_num_1_dense ? 1'h1: input_width_17_num_1_fifo_out_valid;
always_comb begin
  PE_input_width_17_num_1_ready = 1'h1;
  if (mode == 3'h0) begin
    PE_input_width_17_num_1_ready = ~input_width_17_num_1_input_fifo_full;
  end
  else if (mode == 3'h1) begin
    PE_input_width_17_num_1_ready = ~input_width_17_num_1_input_fifo_full;
  end
  else if (mode == 3'h2) begin
    PE_input_width_17_num_1_ready = ~input_width_17_num_1_input_fifo_full;
  end
  else if (mode == 3'h3) begin
    PE_input_width_17_num_1_ready = PE_input_width_17_num_1_dense ? 1'h1: ~input_width_17_num_1_input_fifo_full;
  end
  else if (mode == 3'h4) begin
    PE_input_width_17_num_1_ready = ~input_width_17_num_1_input_fifo_full;
  end
end
assign input_width_17_num_2_fifo_out_valid = ~input_width_17_num_2_input_fifo_empty;
always_comb begin
  input_width_17_num_2_fifo_out_ready = 1'h1;
  if (mode == 3'h0) begin
    input_width_17_num_2_fifo_out_ready = mem_ctrl_intersect_unit_flat_pos_in_0_ready_f_;
  end
  else input_width_17_num_2_fifo_out_ready = 1'h1;
end
always_comb begin
  PE_input_width_17_num_2_ready = 1'h1;
  if (mode == 3'h0) begin
    PE_input_width_17_num_2_ready = ~input_width_17_num_2_input_fifo_full;
  end
  else if (mode == 3'h3) begin
    PE_input_width_17_num_2_ready = 1'h1;
  end
end
assign input_width_17_num_3_fifo_out_valid = ~input_width_17_num_3_input_fifo_empty;
always_comb begin
  input_width_17_num_3_fifo_out_ready = 1'h1;
  if (mode == 3'h0) begin
    input_width_17_num_3_fifo_out_ready = mem_ctrl_intersect_unit_flat_pos_in_1_ready_f_;
  end
  else input_width_17_num_3_fifo_out_ready = 1'h1;
end
always_comb begin
  PE_input_width_17_num_3_ready = 1'h1;
  if (mode == 3'h0) begin
    PE_input_width_17_num_3_ready = ~input_width_17_num_3_input_fifo_full;
  end
  else PE_input_width_17_num_3_ready = 1'h1;
end
assign output_width_17_num_0_fifo_in_ready = ~output_width_17_num_0_output_fifo_full;
always_comb begin
  output_width_17_num_0_fifo_in = 17'h0;
  output_width_17_num_0_fifo_in_valid = 1'h0;
  if (mode == 3'h0) begin
    output_width_17_num_0_fifo_in = mem_ctrl_intersect_unit_flat_coord_out_f_;
    output_width_17_num_0_fifo_in_valid = mem_ctrl_intersect_unit_flat_coord_out_valid_f_;
  end
  else if (mode == 3'h1) begin
    output_width_17_num_0_fifo_in = mem_ctrl_crddrop_flat_cmrg_coord_out_0_f_;
    output_width_17_num_0_fifo_in_valid = mem_ctrl_crddrop_flat_cmrg_coord_out_0_valid_f_;
  end
  else if (mode == 3'h2) begin
    output_width_17_num_0_fifo_in = mem_ctrl_crdhold_flat_cmrg_coord_out_0_f_;
    output_width_17_num_0_fifo_in_valid = mem_ctrl_crdhold_flat_cmrg_coord_out_0_valid_f_;
  end
  else if (mode == 3'h3) begin
    output_width_17_num_0_fifo_in = mem_ctrl_PE_onyx_flat_res_f_;
    output_width_17_num_0_fifo_in_valid = mem_ctrl_PE_onyx_flat_res_valid_f_;
  end
  else if (mode == 3'h4) begin
    output_width_17_num_0_fifo_in = mem_ctrl_Repeat_flat_ref_data_out_f_;
    output_width_17_num_0_fifo_in_valid = mem_ctrl_Repeat_flat_ref_data_out_valid_f_;
  end
  else if (mode == 3'h5) begin
    output_width_17_num_0_fifo_in = mem_ctrl_RepeatSignalGenerator_flat_repsig_data_out_f_;
    output_width_17_num_0_fifo_in_valid = mem_ctrl_RepeatSignalGenerator_flat_repsig_data_out_valid_f_;
  end
  else if (mode == 3'h6) begin
    output_width_17_num_0_fifo_in = mem_ctrl_reg_cr_flat_data_out_f_;
    output_width_17_num_0_fifo_in_valid = mem_ctrl_reg_cr_flat_data_out_valid_f_;
  end
end
assign mem_ctrl_PE_onyx_flat_res_ready_f_ = PE_output_width_17_num_0_dense ? 1'h1: output_width_17_num_0_fifo_in_ready;
always_comb begin
  PE_output_width_17_num_0 = 17'h0;
  if (mode == 3'h0) begin
    PE_output_width_17_num_0 = output_width_17_num_0_output_fifo_data_out;
  end
  else if (mode == 3'h1) begin
    PE_output_width_17_num_0 = output_width_17_num_0_output_fifo_data_out;
  end
  else if (mode == 3'h2) begin
    PE_output_width_17_num_0 = output_width_17_num_0_output_fifo_data_out;
  end
  else if (mode == 3'h3) begin
    PE_output_width_17_num_0 = PE_output_width_17_num_0_dense ? mem_ctrl_PE_onyx_flat_res_f_:
        output_width_17_num_0_output_fifo_data_out;
  end
  else if (mode == 3'h4) begin
    PE_output_width_17_num_0 = output_width_17_num_0_output_fifo_data_out;
  end
  else if (mode == 3'h5) begin
    PE_output_width_17_num_0 = output_width_17_num_0_output_fifo_data_out;
  end
  else if (mode == 3'h6) begin
    PE_output_width_17_num_0 = output_width_17_num_0_output_fifo_data_out;
  end
end
always_comb begin
  PE_output_width_17_num_0_valid = 1'h0;
  if (mode == 3'h0) begin
    PE_output_width_17_num_0_valid = ~output_width_17_num_0_output_fifo_empty;
  end
  else if (mode == 3'h1) begin
    PE_output_width_17_num_0_valid = ~output_width_17_num_0_output_fifo_empty;
  end
  else if (mode == 3'h2) begin
    PE_output_width_17_num_0_valid = ~output_width_17_num_0_output_fifo_empty;
  end
  else if (mode == 3'h3) begin
    PE_output_width_17_num_0_valid = PE_output_width_17_num_0_dense ? 1'h1: ~output_width_17_num_0_output_fifo_empty;
  end
  else if (mode == 3'h4) begin
    PE_output_width_17_num_0_valid = ~output_width_17_num_0_output_fifo_empty;
  end
  else if (mode == 3'h5) begin
    PE_output_width_17_num_0_valid = ~output_width_17_num_0_output_fifo_empty;
  end
  else if (mode == 3'h6) begin
    PE_output_width_17_num_0_valid = ~output_width_17_num_0_output_fifo_empty;
  end
end
assign output_width_17_num_1_fifo_in_ready = ~output_width_17_num_1_output_fifo_full;
always_comb begin
  output_width_17_num_1_fifo_in = 17'h0;
  output_width_17_num_1_fifo_in_valid = 1'h0;
  if (mode == 3'h0) begin
    output_width_17_num_1_fifo_in = mem_ctrl_intersect_unit_flat_pos_out_0_f_;
    output_width_17_num_1_fifo_in_valid = mem_ctrl_intersect_unit_flat_pos_out_0_valid_f_;
  end
  else if (mode == 3'h1) begin
    output_width_17_num_1_fifo_in = mem_ctrl_crddrop_flat_cmrg_coord_out_1_f_;
    output_width_17_num_1_fifo_in_valid = mem_ctrl_crddrop_flat_cmrg_coord_out_1_valid_f_;
  end
  else if (mode == 3'h2) begin
    output_width_17_num_1_fifo_in = mem_ctrl_crdhold_flat_cmrg_coord_out_1_f_;
    output_width_17_num_1_fifo_in_valid = mem_ctrl_crdhold_flat_cmrg_coord_out_1_valid_f_;
  end
end
always_comb begin
  PE_output_width_17_num_1 = 17'h0;
  if (mode == 3'h0) begin
    PE_output_width_17_num_1 = output_width_17_num_1_output_fifo_data_out;
  end
  else if (mode == 3'h1) begin
    PE_output_width_17_num_1 = output_width_17_num_1_output_fifo_data_out;
  end
  else if (mode == 3'h2) begin
    PE_output_width_17_num_1 = output_width_17_num_1_output_fifo_data_out;
  end
end
always_comb begin
  PE_output_width_17_num_1_valid = 1'h0;
  if (mode == 3'h0) begin
    PE_output_width_17_num_1_valid = ~output_width_17_num_1_output_fifo_empty;
  end
  else if (mode == 3'h1) begin
    PE_output_width_17_num_1_valid = ~output_width_17_num_1_output_fifo_empty;
  end
  else if (mode == 3'h2) begin
    PE_output_width_17_num_1_valid = ~output_width_17_num_1_output_fifo_empty;
  end
end
assign output_width_17_num_2_fifo_in_ready = ~output_width_17_num_2_output_fifo_full;
always_comb begin
  output_width_17_num_2_fifo_in = 17'h0;
  output_width_17_num_2_fifo_in_valid = 1'h0;
  output_width_17_num_2_fifo_in = mem_ctrl_intersect_unit_flat_pos_out_1_f_;
  output_width_17_num_2_fifo_in_valid = mem_ctrl_intersect_unit_flat_pos_out_1_valid_f_;
end
always_comb begin
  PE_output_width_17_num_2 = 17'h0;
  if (mode == 3'h0) begin
    PE_output_width_17_num_2 = output_width_17_num_2_output_fifo_data_out;
  end
  else PE_output_width_17_num_2 = 17'h0;
end
always_comb begin
  PE_output_width_17_num_2_valid = 1'h0;
  if (mode == 3'h0) begin
    PE_output_width_17_num_2_valid = ~output_width_17_num_2_output_fifo_empty;
  end
  else PE_output_width_17_num_2_valid = 1'h0;
end
always_comb begin
  PE_output_width_1_num_0 = 1'h0;
  if (mode == 3'h3) begin
    PE_output_width_1_num_0 = mem_ctrl_PE_onyx_flat_res_p_f_;
  end
  else PE_output_width_1_num_0 = 1'h0;
end
assign {mem_ctrl_intersect_unit_flat_intersect_unit_inst_joiner_op, mem_ctrl_intersect_unit_flat_intersect_unit_inst_tile_en} = CONFIG_SPACE[1:0];
assign {mem_ctrl_crddrop_flat_crddrop_inst_cmrg_enable, mem_ctrl_crddrop_flat_crddrop_inst_cmrg_stop_lvl, mem_ctrl_crddrop_flat_crddrop_inst_tile_en} = CONFIG_SPACE[17:0];
assign {mem_ctrl_crdhold_flat_crdhold_inst_cmrg_enable, mem_ctrl_crdhold_flat_crdhold_inst_cmrg_stop_lvl, mem_ctrl_crdhold_flat_crdhold_inst_tile_en} = CONFIG_SPACE[17:0];
assign {mem_ctrl_PE_onyx_flat_PE_onyx_inst_dense_mode, mem_ctrl_PE_onyx_flat_PE_onyx_inst_onyxpeintf_inst, mem_ctrl_PE_onyx_flat_PE_onyx_inst_tile_en} = CONFIG_SPACE[85:0];
assign {mem_ctrl_Repeat_flat_Repeat_inst_root, mem_ctrl_Repeat_flat_Repeat_inst_spacc_mode, mem_ctrl_Repeat_flat_Repeat_inst_stop_lvl, mem_ctrl_Repeat_flat_Repeat_inst_tile_en} = CONFIG_SPACE[18:0];
assign {mem_ctrl_RepeatSignalGenerator_flat_RepeatSignalGenerator_inst_stop_lvl, mem_ctrl_RepeatSignalGenerator_flat_RepeatSignalGenerator_inst_tile_en} = CONFIG_SPACE[16:0];
assign {mem_ctrl_reg_cr_flat_reg_cr_inst_default_value, mem_ctrl_reg_cr_flat_reg_cr_inst_stop_lvl, mem_ctrl_reg_cr_flat_reg_cr_inst_tile_en} = CONFIG_SPACE[32:0];
assign CONFIG_SPACE[31:0] = CONFIG_SPACE_0;
assign CONFIG_SPACE[63:32] = CONFIG_SPACE_1;
assign CONFIG_SPACE[85:64] = CONFIG_SPACE_2;
intersect_unit_flat mem_ctrl_intersect_unit_flat (
  .clk(mem_ctrl_intersect_unit_flat_clk),
  .clk_en(clk_en),
  .coord_in_0_f_(input_width_17_num_0_fifo_out),
  .coord_in_0_valid_f_(input_width_17_num_0_fifo_out_valid),
  .coord_in_1_f_(input_width_17_num_1_fifo_out),
  .coord_in_1_valid_f_(input_width_17_num_1_fifo_out_valid),
  .coord_out_ready_f_(output_width_17_num_0_fifo_in_ready),
  .flush(flush),
  .intersect_unit_inst_joiner_op(mem_ctrl_intersect_unit_flat_intersect_unit_inst_joiner_op),
  .intersect_unit_inst_tile_en(mem_ctrl_intersect_unit_flat_intersect_unit_inst_tile_en),
  .pos_in_0_f_(input_width_17_num_2_fifo_out),
  .pos_in_0_valid_f_(input_width_17_num_2_fifo_out_valid),
  .pos_in_1_f_(input_width_17_num_3_fifo_out),
  .pos_in_1_valid_f_(input_width_17_num_3_fifo_out_valid),
  .pos_out_0_ready_f_(output_width_17_num_1_fifo_in_ready),
  .pos_out_1_ready_f_(output_width_17_num_2_fifo_in_ready),
  .rst_n(rst_n),
  .coord_in_0_ready_f_(mem_ctrl_intersect_unit_flat_coord_in_0_ready_f_),
  .coord_in_1_ready_f_(mem_ctrl_intersect_unit_flat_coord_in_1_ready_f_),
  .coord_out_f_(mem_ctrl_intersect_unit_flat_coord_out_f_),
  .coord_out_valid_f_(mem_ctrl_intersect_unit_flat_coord_out_valid_f_),
  .pos_in_0_ready_f_(mem_ctrl_intersect_unit_flat_pos_in_0_ready_f_),
  .pos_in_1_ready_f_(mem_ctrl_intersect_unit_flat_pos_in_1_ready_f_),
  .pos_out_0_f_(mem_ctrl_intersect_unit_flat_pos_out_0_f_),
  .pos_out_0_valid_f_(mem_ctrl_intersect_unit_flat_pos_out_0_valid_f_),
  .pos_out_1_f_(mem_ctrl_intersect_unit_flat_pos_out_1_f_),
  .pos_out_1_valid_f_(mem_ctrl_intersect_unit_flat_pos_out_1_valid_f_)
);

crddrop_flat mem_ctrl_crddrop_flat (
  .clk(mem_ctrl_crddrop_flat_clk),
  .clk_en(clk_en),
  .cmrg_coord_in_0_f_(input_width_17_num_0_fifo_out),
  .cmrg_coord_in_0_valid_f_(input_width_17_num_0_fifo_out_valid),
  .cmrg_coord_in_1_f_(input_width_17_num_1_fifo_out),
  .cmrg_coord_in_1_valid_f_(input_width_17_num_1_fifo_out_valid),
  .cmrg_coord_out_0_ready_f_(output_width_17_num_0_fifo_in_ready),
  .cmrg_coord_out_1_ready_f_(output_width_17_num_1_fifo_in_ready),
  .crddrop_inst_cmrg_enable(mem_ctrl_crddrop_flat_crddrop_inst_cmrg_enable),
  .crddrop_inst_cmrg_stop_lvl(mem_ctrl_crddrop_flat_crddrop_inst_cmrg_stop_lvl),
  .crddrop_inst_tile_en(mem_ctrl_crddrop_flat_crddrop_inst_tile_en),
  .flush(flush),
  .rst_n(rst_n),
  .cmrg_coord_in_0_ready_f_(mem_ctrl_crddrop_flat_cmrg_coord_in_0_ready_f_),
  .cmrg_coord_in_1_ready_f_(mem_ctrl_crddrop_flat_cmrg_coord_in_1_ready_f_),
  .cmrg_coord_out_0_f_(mem_ctrl_crddrop_flat_cmrg_coord_out_0_f_),
  .cmrg_coord_out_0_valid_f_(mem_ctrl_crddrop_flat_cmrg_coord_out_0_valid_f_),
  .cmrg_coord_out_1_f_(mem_ctrl_crddrop_flat_cmrg_coord_out_1_f_),
  .cmrg_coord_out_1_valid_f_(mem_ctrl_crddrop_flat_cmrg_coord_out_1_valid_f_)
);

crdhold_flat mem_ctrl_crdhold_flat (
  .clk(mem_ctrl_crdhold_flat_clk),
  .clk_en(clk_en),
  .cmrg_coord_in_0_f_(input_width_17_num_0_fifo_out),
  .cmrg_coord_in_0_valid_f_(input_width_17_num_0_fifo_out_valid),
  .cmrg_coord_in_1_f_(input_width_17_num_1_fifo_out),
  .cmrg_coord_in_1_valid_f_(input_width_17_num_1_fifo_out_valid),
  .cmrg_coord_out_0_ready_f_(output_width_17_num_0_fifo_in_ready),
  .cmrg_coord_out_1_ready_f_(output_width_17_num_1_fifo_in_ready),
  .crdhold_inst_cmrg_enable(mem_ctrl_crdhold_flat_crdhold_inst_cmrg_enable),
  .crdhold_inst_cmrg_stop_lvl(mem_ctrl_crdhold_flat_crdhold_inst_cmrg_stop_lvl),
  .crdhold_inst_tile_en(mem_ctrl_crdhold_flat_crdhold_inst_tile_en),
  .flush(flush),
  .rst_n(rst_n),
  .cmrg_coord_in_0_ready_f_(mem_ctrl_crdhold_flat_cmrg_coord_in_0_ready_f_),
  .cmrg_coord_in_1_ready_f_(mem_ctrl_crdhold_flat_cmrg_coord_in_1_ready_f_),
  .cmrg_coord_out_0_f_(mem_ctrl_crdhold_flat_cmrg_coord_out_0_f_),
  .cmrg_coord_out_0_valid_f_(mem_ctrl_crdhold_flat_cmrg_coord_out_0_valid_f_),
  .cmrg_coord_out_1_f_(mem_ctrl_crdhold_flat_cmrg_coord_out_1_f_),
  .cmrg_coord_out_1_valid_f_(mem_ctrl_crdhold_flat_cmrg_coord_out_1_valid_f_)
);

PE_onyx_flat mem_ctrl_PE_onyx_flat (
  .PE_onyx_inst_dense_mode(mem_ctrl_PE_onyx_flat_PE_onyx_inst_dense_mode),
  .PE_onyx_inst_onyxpeintf_inst(mem_ctrl_PE_onyx_flat_PE_onyx_inst_onyxpeintf_inst),
  .PE_onyx_inst_tile_en(mem_ctrl_PE_onyx_flat_PE_onyx_inst_tile_en),
  .bit0_f_(PE_input_width_1_num_0),
  .bit1_f_(PE_input_width_1_num_1),
  .bit2_f_(PE_input_width_1_num_2),
  .clk(mem_ctrl_PE_onyx_flat_clk),
  .clk_en(clk_en),
  .data0_f_(mem_ctrl_PE_onyx_flat_data0_f_),
  .data0_valid_f_(mem_ctrl_PE_onyx_flat_data0_valid_f_),
  .data1_f_(mem_ctrl_PE_onyx_flat_data1_f_),
  .data1_valid_f_(mem_ctrl_PE_onyx_flat_data1_valid_f_),
  .data2_f_(PE_input_width_17_num_2),
  .flush(flush),
  .res_ready_f_(mem_ctrl_PE_onyx_flat_res_ready_f_),
  .rst_n(rst_n),
  .PE_onyx_inst_onyxpeintf_O2(PE_onyx_inst_onyxpeintf_O2),
  .PE_onyx_inst_onyxpeintf_O3(PE_onyx_inst_onyxpeintf_O3),
  .PE_onyx_inst_onyxpeintf_O4(PE_onyx_inst_onyxpeintf_O4),
  .data0_ready_f_(mem_ctrl_PE_onyx_flat_data0_ready_f_),
  .data1_ready_f_(mem_ctrl_PE_onyx_flat_data1_ready_f_),
  .res_f_(mem_ctrl_PE_onyx_flat_res_f_),
  .res_p_f_(mem_ctrl_PE_onyx_flat_res_p_f_),
  .res_valid_f_(mem_ctrl_PE_onyx_flat_res_valid_f_)
);

Repeat_flat mem_ctrl_Repeat_flat (
  .Repeat_inst_root(mem_ctrl_Repeat_flat_Repeat_inst_root),
  .Repeat_inst_spacc_mode(mem_ctrl_Repeat_flat_Repeat_inst_spacc_mode),
  .Repeat_inst_stop_lvl(mem_ctrl_Repeat_flat_Repeat_inst_stop_lvl),
  .Repeat_inst_tile_en(mem_ctrl_Repeat_flat_Repeat_inst_tile_en),
  .clk(mem_ctrl_Repeat_flat_clk),
  .clk_en(clk_en),
  .flush(flush),
  .proc_data_in_f_(input_width_17_num_0_fifo_out),
  .proc_data_in_valid_f_(input_width_17_num_0_fifo_out_valid),
  .ref_data_out_ready_f_(output_width_17_num_0_fifo_in_ready),
  .repsig_data_in_f_(input_width_17_num_1_fifo_out),
  .repsig_data_in_valid_f_(input_width_17_num_1_fifo_out_valid),
  .rst_n(rst_n),
  .proc_data_in_ready_f_(mem_ctrl_Repeat_flat_proc_data_in_ready_f_),
  .ref_data_out_f_(mem_ctrl_Repeat_flat_ref_data_out_f_),
  .ref_data_out_valid_f_(mem_ctrl_Repeat_flat_ref_data_out_valid_f_),
  .repsig_data_in_ready_f_(mem_ctrl_Repeat_flat_repsig_data_in_ready_f_)
);

RepeatSignalGenerator_flat mem_ctrl_RepeatSignalGenerator_flat (
  .RepeatSignalGenerator_inst_stop_lvl(mem_ctrl_RepeatSignalGenerator_flat_RepeatSignalGenerator_inst_stop_lvl),
  .RepeatSignalGenerator_inst_tile_en(mem_ctrl_RepeatSignalGenerator_flat_RepeatSignalGenerator_inst_tile_en),
  .base_data_in_f_(input_width_17_num_0_fifo_out),
  .base_data_in_valid_f_(input_width_17_num_0_fifo_out_valid),
  .clk(mem_ctrl_RepeatSignalGenerator_flat_clk),
  .clk_en(clk_en),
  .flush(flush),
  .repsig_data_out_ready_f_(output_width_17_num_0_fifo_in_ready),
  .rst_n(rst_n),
  .base_data_in_ready_f_(mem_ctrl_RepeatSignalGenerator_flat_base_data_in_ready_f_),
  .repsig_data_out_f_(mem_ctrl_RepeatSignalGenerator_flat_repsig_data_out_f_),
  .repsig_data_out_valid_f_(mem_ctrl_RepeatSignalGenerator_flat_repsig_data_out_valid_f_)
);

reg_cr_flat mem_ctrl_reg_cr_flat (
  .clk(mem_ctrl_reg_cr_flat_clk),
  .clk_en(clk_en),
  .data_in_f_(input_width_17_num_0_fifo_out),
  .data_in_valid_f_(input_width_17_num_0_fifo_out_valid),
  .data_out_ready_f_(output_width_17_num_0_fifo_in_ready),
  .flush(flush),
  .reg_cr_inst_default_value(mem_ctrl_reg_cr_flat_reg_cr_inst_default_value),
  .reg_cr_inst_stop_lvl(mem_ctrl_reg_cr_flat_reg_cr_inst_stop_lvl),
  .reg_cr_inst_tile_en(mem_ctrl_reg_cr_flat_reg_cr_inst_tile_en),
  .rst_n(rst_n),
  .data_in_ready_f_(mem_ctrl_reg_cr_flat_data_in_ready_f_),
  .data_out_f_(mem_ctrl_reg_cr_flat_data_out_f_),
  .data_out_valid_f_(mem_ctrl_reg_cr_flat_data_out_valid_f_)
);

reg_fifo_depth_2_w_17_afd_2 input_width_17_num_0_input_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(PE_input_width_17_num_0),
  .flush(flush),
  .pop(input_width_17_num_0_fifo_out_ready),
  .push(PE_input_width_17_num_0_valid),
  .rst_n(rst_n),
  .data_out(input_width_17_num_0_fifo_out),
  .empty(input_width_17_num_0_input_fifo_empty),
  .full(input_width_17_num_0_input_fifo_full)
);

reg_fifo_depth_2_w_17_afd_2 input_width_17_num_1_input_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(PE_input_width_17_num_1),
  .flush(flush),
  .pop(input_width_17_num_1_fifo_out_ready),
  .push(PE_input_width_17_num_1_valid),
  .rst_n(rst_n),
  .data_out(input_width_17_num_1_fifo_out),
  .empty(input_width_17_num_1_input_fifo_empty),
  .full(input_width_17_num_1_input_fifo_full)
);

reg_fifo_depth_2_w_17_afd_2 input_width_17_num_2_input_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(PE_input_width_17_num_2),
  .flush(flush),
  .pop(input_width_17_num_2_fifo_out_ready),
  .push(PE_input_width_17_num_2_valid),
  .rst_n(rst_n),
  .data_out(input_width_17_num_2_fifo_out),
  .empty(input_width_17_num_2_input_fifo_empty),
  .full(input_width_17_num_2_input_fifo_full)
);

reg_fifo_depth_2_w_17_afd_2 input_width_17_num_3_input_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(PE_input_width_17_num_3),
  .flush(flush),
  .pop(input_width_17_num_3_fifo_out_ready),
  .push(PE_input_width_17_num_3_valid),
  .rst_n(rst_n),
  .data_out(input_width_17_num_3_fifo_out),
  .empty(input_width_17_num_3_input_fifo_empty),
  .full(input_width_17_num_3_input_fifo_full)
);

reg_fifo_depth_2_w_17_afd_2 output_width_17_num_0_output_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(output_width_17_num_0_fifo_in),
  .flush(flush),
  .pop(PE_output_width_17_num_0_ready),
  .push(output_width_17_num_0_fifo_in_valid),
  .rst_n(rst_n),
  .data_out(output_width_17_num_0_output_fifo_data_out),
  .empty(output_width_17_num_0_output_fifo_empty),
  .full(output_width_17_num_0_output_fifo_full)
);

reg_fifo_depth_2_w_17_afd_2 output_width_17_num_1_output_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(output_width_17_num_1_fifo_in),
  .flush(flush),
  .pop(PE_output_width_17_num_1_ready),
  .push(output_width_17_num_1_fifo_in_valid),
  .rst_n(rst_n),
  .data_out(output_width_17_num_1_output_fifo_data_out),
  .empty(output_width_17_num_1_output_fifo_empty),
  .full(output_width_17_num_1_output_fifo_full)
);

reg_fifo_depth_2_w_17_afd_2 output_width_17_num_2_output_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(output_width_17_num_2_fifo_in),
  .flush(flush),
  .pop(PE_output_width_17_num_2_ready),
  .push(output_width_17_num_2_fifo_in_valid),
  .rst_n(rst_n),
  .data_out(output_width_17_num_2_output_fifo_data_out),
  .empty(output_width_17_num_2_output_fifo_empty),
  .full(output_width_17_num_2_output_fifo_full)
);

endmodule   // PE_inner

module PE_inner_W (
  input logic [31:0] CONFIG_SPACE_0,
  input logic [31:0] CONFIG_SPACE_1,
  input logic [21:0] CONFIG_SPACE_2,
  input logic [0:0] [16:0] PE_input_width_17_num_0,
  input logic PE_input_width_17_num_0_dense,
  input logic PE_input_width_17_num_0_valid,
  input logic [0:0] [16:0] PE_input_width_17_num_1,
  input logic PE_input_width_17_num_1_dense,
  input logic PE_input_width_17_num_1_valid,
  input logic [0:0] [16:0] PE_input_width_17_num_2,
  input logic PE_input_width_17_num_2_valid,
  input logic [0:0] [16:0] PE_input_width_17_num_3,
  input logic PE_input_width_17_num_3_valid,
  input logic PE_input_width_1_num_0,
  input logic PE_input_width_1_num_1,
  input logic PE_input_width_1_num_2,
  input logic PE_output_width_17_num_0_dense,
  input logic PE_output_width_17_num_0_ready,
  input logic PE_output_width_17_num_1_ready,
  input logic PE_output_width_17_num_2_ready,
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [2:0] mode,
  input logic rst_n,
  input logic tile_en,
  output logic PE_input_width_17_num_0_ready,
  output logic PE_input_width_17_num_1_ready,
  output logic PE_input_width_17_num_2_ready,
  output logic PE_input_width_17_num_3_ready,
  output logic [15:0] PE_onyx_inst_onyxpeintf_O2,
  output logic [15:0] PE_onyx_inst_onyxpeintf_O3,
  output logic [15:0] PE_onyx_inst_onyxpeintf_O4,
  output logic [0:0] [16:0] PE_output_width_17_num_0,
  output logic PE_output_width_17_num_0_valid,
  output logic [0:0] [16:0] PE_output_width_17_num_1,
  output logic PE_output_width_17_num_1_valid,
  output logic [0:0] [16:0] PE_output_width_17_num_2,
  output logic PE_output_width_17_num_2_valid,
  output logic PE_output_width_1_num_0
);

PE_inner PE_inner (
  .CONFIG_SPACE_0(CONFIG_SPACE_0),
  .CONFIG_SPACE_1(CONFIG_SPACE_1),
  .CONFIG_SPACE_2(CONFIG_SPACE_2),
  .PE_input_width_17_num_0(PE_input_width_17_num_0),
  .PE_input_width_17_num_0_dense(PE_input_width_17_num_0_dense),
  .PE_input_width_17_num_0_valid(PE_input_width_17_num_0_valid),
  .PE_input_width_17_num_1(PE_input_width_17_num_1),
  .PE_input_width_17_num_1_dense(PE_input_width_17_num_1_dense),
  .PE_input_width_17_num_1_valid(PE_input_width_17_num_1_valid),
  .PE_input_width_17_num_2(PE_input_width_17_num_2),
  .PE_input_width_17_num_2_valid(PE_input_width_17_num_2_valid),
  .PE_input_width_17_num_3(PE_input_width_17_num_3),
  .PE_input_width_17_num_3_valid(PE_input_width_17_num_3_valid),
  .PE_input_width_1_num_0(PE_input_width_1_num_0),
  .PE_input_width_1_num_1(PE_input_width_1_num_1),
  .PE_input_width_1_num_2(PE_input_width_1_num_2),
  .PE_output_width_17_num_0_dense(PE_output_width_17_num_0_dense),
  .PE_output_width_17_num_0_ready(PE_output_width_17_num_0_ready),
  .PE_output_width_17_num_1_ready(PE_output_width_17_num_1_ready),
  .PE_output_width_17_num_2_ready(PE_output_width_17_num_2_ready),
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mode(mode),
  .rst_n(rst_n),
  .tile_en(tile_en),
  .PE_input_width_17_num_0_ready(PE_input_width_17_num_0_ready),
  .PE_input_width_17_num_1_ready(PE_input_width_17_num_1_ready),
  .PE_input_width_17_num_2_ready(PE_input_width_17_num_2_ready),
  .PE_input_width_17_num_3_ready(PE_input_width_17_num_3_ready),
  .PE_onyx_inst_onyxpeintf_O2(PE_onyx_inst_onyxpeintf_O2),
  .PE_onyx_inst_onyxpeintf_O3(PE_onyx_inst_onyxpeintf_O3),
  .PE_onyx_inst_onyxpeintf_O4(PE_onyx_inst_onyxpeintf_O4),
  .PE_output_width_17_num_0(PE_output_width_17_num_0),
  .PE_output_width_17_num_0_valid(PE_output_width_17_num_0_valid),
  .PE_output_width_17_num_1(PE_output_width_17_num_1),
  .PE_output_width_17_num_1_valid(PE_output_width_17_num_1_valid),
  .PE_output_width_17_num_2(PE_output_width_17_num_2),
  .PE_output_width_17_num_2_valid(PE_output_width_17_num_2_valid),
  .PE_output_width_1_num_0(PE_output_width_1_num_0)
);

endmodule   // PE_inner_W

module PE_onyx (
  input logic bit0,
  input logic bit1,
  input logic bit2,
  input logic clk,
  input logic clk_en,
  input logic [16:0] data0,
  input logic data0_valid,
  input logic [16:0] data1,
  input logic data1_valid,
  input logic [16:0] data2,
  input logic dense_mode,
  input logic flush,
  input logic [83:0] onyxpeintf_inst,
  input logic res_ready,
  input logic rst_n,
  input logic tile_en,
  output logic data0_ready,
  output logic data1_ready,
  output logic [15:0] onyxpeintf_O2,
  output logic [15:0] onyxpeintf_O3,
  output logic [15:0] onyxpeintf_O4,
  output logic [16:0] res,
  output logic res_p,
  output logic res_valid
);

logic [15:0] data_to_fifo;
logic gclk;
logic [1:0][16:0] infifo_in_packed;
logic [1:0][15:0] infifo_out_data;
logic [1:0] infifo_out_eos;
logic infifo_out_maybe_0;
logic infifo_out_maybe_1;
logic [1:0][16:0] infifo_out_packed;
logic [1:0] infifo_out_valid;
logic [1:0] infifo_pop;
logic infifo_push_0;
logic infifo_push_1;
logic [0:0][16:0] input_fifo_0_data_out;
logic input_fifo_0_empty;
logic input_fifo_0_full;
logic [0:0][16:0] input_fifo_1_data_out;
logic input_fifo_1_empty;
logic input_fifo_1_full;
logic onyxpeintf_ASYNCRESET;
logic [15:0] onyxpeintf_data0;
logic [15:0] onyxpeintf_data1;
logic outfifo_full;
logic outfifo_in_eos;
logic [16:0] outfifo_in_packed;
logic [16:0] outfifo_out_packed;
logic outfifo_pop;
logic outfifo_push;
logic output_fifo_empty;
logic [15:0] pe_output;
assign gclk = clk & tile_en;
assign data0_ready = dense_mode ? 1'h1: ~input_fifo_0_full;
assign data1_ready = dense_mode ? 1'h1: ~input_fifo_1_full;
assign infifo_in_packed[0] = data0;
assign infifo_out_eos[0] = infifo_out_packed[0][16];
assign infifo_out_data[0] = infifo_out_packed[0][15:0];
assign infifo_in_packed[1] = data1;
assign infifo_out_eos[1] = infifo_out_packed[1][16];
assign infifo_out_data[1] = infifo_out_packed[1][15:0];
assign infifo_push_0 = data0_valid;
assign infifo_push_1 = data1_valid;
assign infifo_out_packed[0] = input_fifo_0_data_out;
assign infifo_out_packed[1] = input_fifo_1_data_out;
assign infifo_out_valid[0] = ~input_fifo_0_empty;
assign infifo_out_valid[1] = ~input_fifo_1_empty;
assign outfifo_in_packed[16] = outfifo_in_eos;
assign outfifo_in_packed[15:0] = data_to_fifo;
assign res = dense_mode ? 17'(pe_output): outfifo_out_packed;
assign res_valid = dense_mode ? 1'h1: ~output_fifo_empty;
assign outfifo_pop = res_ready;
assign infifo_out_maybe_0 = infifo_out_eos[0] & infifo_out_valid[0] & (infifo_out_data[0][9:8] == 2'h2);
assign infifo_out_maybe_1 = infifo_out_eos[1] & infifo_out_valid[1] & (infifo_out_data[1][9:8] == 2'h2);
assign onyxpeintf_ASYNCRESET = ~rst_n;
assign onyxpeintf_data0 = dense_mode ? data0[15:0]: infifo_out_maybe_0 ? 16'h0: infifo_out_data[0];
assign onyxpeintf_data1 = dense_mode ? data1[15:0]: infifo_out_maybe_1 ? 16'h0: infifo_out_data[1];
always_comb begin
  outfifo_push = 1'h0;
  outfifo_in_eos = 1'h0;
  data_to_fifo = 16'h0;
  infifo_pop[0] = 1'h0;
  infifo_pop[1] = 1'h0;
  if ((&infifo_out_valid) & (~outfifo_full) & (~dense_mode)) begin
    if (~(&infifo_out_eos)) begin
      outfifo_push = 1'h1;
      outfifo_in_eos = 1'h0;
      data_to_fifo = pe_output;
      infifo_pop[0] = 1'h1;
      infifo_pop[1] = 1'h1;
    end
    else begin
      outfifo_push = 1'h1;
      outfifo_in_eos = 1'h1;
      data_to_fifo = infifo_out_data[0];
      infifo_pop[0] = 1'h1;
      infifo_pop[1] = 1'h1;
    end
  end
end
reg_fifo_depth_0_w_17_afd_2 input_fifo_0 (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(infifo_in_packed[0]),
  .flush(flush),
  .pop(infifo_pop[0]),
  .push(infifo_push_0),
  .rst_n(rst_n),
  .data_out(input_fifo_0_data_out),
  .empty(input_fifo_0_empty),
  .full(input_fifo_0_full)
);

reg_fifo_depth_0_w_17_afd_2 input_fifo_1 (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(infifo_in_packed[1]),
  .flush(flush),
  .pop(infifo_pop[1]),
  .push(infifo_push_1),
  .rst_n(rst_n),
  .data_out(input_fifo_1_data_out),
  .empty(input_fifo_1_empty),
  .full(input_fifo_1_full)
);

reg_fifo_depth_2_w_17_afd_2 output_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(outfifo_in_packed),
  .flush(flush),
  .pop(outfifo_pop),
  .push(outfifo_push),
  .rst_n(rst_n),
  .data_out(outfifo_out_packed),
  .empty(output_fifo_empty),
  .full(outfifo_full)
);

PEGEN_PE onyxpeintf (
  .ASYNCRESET(onyxpeintf_ASYNCRESET),
  .CLK(gclk),
  .bit0(bit0),
  .bit1(bit1),
  .bit2(bit2),
  .clk_en(clk_en),
  .data0(onyxpeintf_data0),
  .data1(onyxpeintf_data1),
  .data2(data2[15:0]),
  .inst(onyxpeintf_inst),
  .O0(pe_output),
  .O1(res_p),
  .O2(onyxpeintf_O2),
  .O3(onyxpeintf_O3),
  .O4(onyxpeintf_O4)
);

endmodule   // PE_onyx

module PE_onyx_flat (
  input logic PE_onyx_inst_dense_mode,
  input logic [83:0] PE_onyx_inst_onyxpeintf_inst,
  input logic PE_onyx_inst_tile_en,
  input logic bit0_f_,
  input logic bit1_f_,
  input logic bit2_f_,
  input logic clk,
  input logic clk_en,
  input logic [0:0] [16:0] data0_f_,
  input logic data0_valid_f_,
  input logic [0:0] [16:0] data1_f_,
  input logic data1_valid_f_,
  input logic [0:0] [16:0] data2_f_,
  input logic flush,
  input logic res_ready_f_,
  input logic rst_n,
  output logic [15:0] PE_onyx_inst_onyxpeintf_O2,
  output logic [15:0] PE_onyx_inst_onyxpeintf_O3,
  output logic [15:0] PE_onyx_inst_onyxpeintf_O4,
  output logic data0_ready_f_,
  output logic data1_ready_f_,
  output logic [0:0] [16:0] res_f_,
  output logic res_p_f_,
  output logic res_valid_f_
);

PE_onyx PE_onyx_inst (
  .bit0(bit0_f_),
  .bit1(bit1_f_),
  .bit2(bit2_f_),
  .clk(clk),
  .clk_en(clk_en),
  .data0(data0_f_),
  .data0_valid(data0_valid_f_),
  .data1(data1_f_),
  .data1_valid(data1_valid_f_),
  .data2(data2_f_),
  .dense_mode(PE_onyx_inst_dense_mode),
  .flush(flush),
  .onyxpeintf_inst(PE_onyx_inst_onyxpeintf_inst),
  .res_ready(res_ready_f_),
  .rst_n(rst_n),
  .tile_en(PE_onyx_inst_tile_en),
  .data0_ready(data0_ready_f_),
  .data1_ready(data1_ready_f_),
  .onyxpeintf_O2(PE_onyx_inst_onyxpeintf_O2),
  .onyxpeintf_O3(PE_onyx_inst_onyxpeintf_O3),
  .onyxpeintf_O4(PE_onyx_inst_onyxpeintf_O4),
  .res(res_f_),
  .res_p(res_p_f_),
  .res_valid(res_valid_f_)
);

endmodule   // PE_onyx_flat

module Repeat (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [16:0] proc_data_in,
  input logic proc_data_in_valid,
  input logic ref_data_out_ready,
  input logic [16:0] repsig_data_in,
  input logic repsig_data_in_valid,
  input logic root,
  input logic rst_n,
  input logic spacc_mode,
  input logic [15:0] stop_lvl,
  input logic tile_en,
  output logic proc_data_in_ready,
  output logic [16:0] ref_data_out,
  output logic ref_data_out_valid,
  output logic repsig_data_in_ready
);

typedef enum logic[2:0] {
  DONE = 3'h0,
  INJECT0 = 3'h1,
  INJECT1 = 3'h2,
  PASS_REPEAT = 3'h3,
  PASS_STOP = 3'h4,
  START = 3'h5
} repeat_fsm_state;
logic clr_last_pushed_data;
logic gclk;
logic proc_done;
logic proc_fifo_full;
logic [15:0] proc_fifo_inject_data;
logic proc_fifo_inject_eos;
logic proc_fifo_inject_push;
logic [15:0] proc_fifo_out_data;
logic proc_fifo_out_eos;
logic proc_fifo_pop;
logic proc_fifo_push;
logic proc_fifo_valid;
logic [0:0][16:0] proc_in_fifo_data_in;
logic [0:0][16:0] proc_in_fifo_data_out;
logic proc_in_fifo_empty;
logic proc_in_fifo_full;
logic proc_stop;
logic ref_fifo_full;
logic [15:0] ref_fifo_in_data;
logic ref_fifo_in_eos;
logic ref_fifo_push;
logic ref_maybe;
logic [0:0][16:0] ref_out_fifo_data_in;
logic ref_out_fifo_empty;
repeat_fsm_state repeat_fsm_current_state;
repeat_fsm_state repeat_fsm_next_state;
logic repsig_done;
logic [15:0] repsig_fifo_out_data;
logic repsig_fifo_out_eos;
logic repsig_fifo_pop;
logic repsig_fifo_valid;
logic [0:0][16:0] repsig_in_fifo_data_out;
logic repsig_in_fifo_empty;
logic repsig_in_fifo_full;
logic repsig_stop;
logic seen_root_eos_sticky;
logic seen_root_eos_was_high;
logic set_last_pushed_data;
logic set_last_pushed_data_sticky;
logic set_last_pushed_data_was_high;
assign gclk = clk & tile_en;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    set_last_pushed_data_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      set_last_pushed_data_was_high <= 1'h0;
    end
    else if (clr_last_pushed_data) begin
      set_last_pushed_data_was_high <= 1'h0;
    end
    else if (set_last_pushed_data) begin
      set_last_pushed_data_was_high <= 1'h1;
    end
  end
end
assign set_last_pushed_data_sticky = set_last_pushed_data_was_high;
assign {repsig_fifo_out_eos, repsig_fifo_out_data} = repsig_in_fifo_data_out;
assign repsig_data_in_ready = ~repsig_in_fifo_full;
assign repsig_fifo_valid = ~repsig_in_fifo_empty;
assign proc_fifo_push = root ? proc_fifo_inject_push: proc_data_in_valid;
assign proc_in_fifo_data_in = root ? {proc_fifo_inject_eos, proc_fifo_inject_data}: proc_data_in;
assign {proc_fifo_out_eos, proc_fifo_out_data} = proc_in_fifo_data_out;
assign proc_data_in_ready = ~proc_in_fifo_full;
assign proc_fifo_full = proc_in_fifo_full;
assign proc_fifo_valid = ~proc_in_fifo_empty;
assign ref_out_fifo_data_in = {ref_fifo_in_eos, ref_fifo_in_data};
assign ref_data_out_valid = ~ref_out_fifo_empty;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    seen_root_eos_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      seen_root_eos_was_high <= 1'h0;
    end
    else if (1'h0) begin
      seen_root_eos_was_high <= 1'h0;
    end
    else if ((proc_fifo_out_data == 16'h0) & proc_fifo_out_eos & proc_fifo_valid) begin
      seen_root_eos_was_high <= 1'h1;
    end
  end
end
assign seen_root_eos_sticky = ((proc_fifo_out_data == 16'h0) & proc_fifo_out_eos & proc_fifo_valid) |
    seen_root_eos_was_high;
assign proc_stop = (proc_fifo_out_data[9:8] == 2'h0) & proc_fifo_out_eos & proc_fifo_valid;
assign proc_done = (proc_fifo_out_data[9:8] == 2'h1) & proc_fifo_out_eos & proc_fifo_valid;
assign repsig_stop = (repsig_fifo_out_data[9:8] == 2'h0) & repsig_fifo_out_eos & repsig_fifo_valid;
assign repsig_done = (repsig_fifo_out_data[9:8] == 2'h1) & repsig_fifo_out_eos & repsig_fifo_valid;
assign ref_maybe = proc_fifo_valid & proc_fifo_out_eos & (proc_fifo_out_data[9:8] == 2'h2);

always_ff @(posedge clk, negedge rst_n) begin
  if (!rst_n) begin
    repeat_fsm_current_state <= START;
  end
  else if (clk_en) begin
    if (flush) begin
      repeat_fsm_current_state <= START;
    end
    else repeat_fsm_current_state <= repeat_fsm_next_state;
  end
end
always_comb begin
  repeat_fsm_next_state = repeat_fsm_current_state;
  unique case (repeat_fsm_current_state)
    DONE: begin
        if ((~ref_fifo_full) & proc_done & repsig_done) begin
          repeat_fsm_next_state = START;
        end
      end
    INJECT0: begin
        if (~proc_fifo_full) begin
          repeat_fsm_next_state = INJECT1;
        end
        else repeat_fsm_next_state = INJECT0;
      end
    INJECT1: begin
        if (~proc_fifo_full) begin
          repeat_fsm_next_state = PASS_REPEAT;
        end
        else repeat_fsm_next_state = INJECT1;
      end
    PASS_REPEAT: begin
        if (proc_done) begin
          repeat_fsm_next_state = DONE;
        end
        else if (repsig_fifo_out_eos & repsig_fifo_valid & (repsig_fifo_out_data[9:8] == 2'h0)) begin
          repeat_fsm_next_state = PASS_STOP;
        end
        else repeat_fsm_next_state = PASS_REPEAT;
      end
    PASS_STOP: begin
        if (proc_fifo_valid & (~proc_stop) & (~ref_fifo_full)) begin
          repeat_fsm_next_state = PASS_REPEAT;
        end
        else repeat_fsm_next_state = PASS_STOP;
      end
    START: begin
        if (root & tile_en) begin
          repeat_fsm_next_state = INJECT0;
        end
        else if ((~root) & tile_en) begin
          repeat_fsm_next_state = PASS_REPEAT;
        end
        else repeat_fsm_next_state = START;
      end
    default: repeat_fsm_next_state = repeat_fsm_current_state;
  endcase
end
always_comb begin
  unique case (repeat_fsm_current_state)
    DONE: begin :repeat_fsm_DONE_Output
        ref_fifo_in_data = proc_fifo_out_data;
        ref_fifo_in_eos = 1'h1;
        ref_fifo_push = (~ref_fifo_full) & proc_done & repsig_done;
        proc_fifo_pop = (~ref_fifo_full) & proc_done & repsig_done;
        repsig_fifo_pop = (~ref_fifo_full) & proc_done & repsig_done;
        proc_fifo_inject_push = 1'h0;
        proc_fifo_inject_data = 16'h0;
        proc_fifo_inject_eos = 1'h0;
      end :repeat_fsm_DONE_Output
    INJECT0: begin :repeat_fsm_INJECT0_Output
        ref_fifo_in_data = 16'h0;
        ref_fifo_in_eos = 1'h0;
        ref_fifo_push = 1'h0;
        proc_fifo_pop = 1'h0;
        repsig_fifo_pop = 1'h0;
        proc_fifo_inject_push = 1'h1;
        proc_fifo_inject_data = 16'h0;
        proc_fifo_inject_eos = 1'h0;
      end :repeat_fsm_INJECT0_Output
    INJECT1: begin :repeat_fsm_INJECT1_Output
        ref_fifo_in_data = 16'h0;
        ref_fifo_in_eos = 1'h0;
        ref_fifo_push = 1'h0;
        proc_fifo_pop = 1'h0;
        repsig_fifo_pop = 1'h0;
        proc_fifo_inject_push = 1'h1;
        proc_fifo_inject_data = 16'h100;
        proc_fifo_inject_eos = 1'h1;
      end :repeat_fsm_INJECT1_Output
    PASS_REPEAT: begin :repeat_fsm_PASS_REPEAT_Output
        ref_fifo_in_data = proc_fifo_out_data;
        ref_fifo_in_eos = ref_maybe;
        ref_fifo_push = repsig_fifo_valid & proc_fifo_valid & (~repsig_fifo_out_eos) & (~proc_done) &
            (~ref_fifo_full);
        proc_fifo_pop = ((repsig_fifo_valid & repsig_fifo_out_eos & (~spacc_mode)) | (spacc_mode &
            repsig_done)) & (~proc_done);
        repsig_fifo_pop = (~ref_fifo_full) & repsig_fifo_valid & (~repsig_fifo_out_eos) & proc_fifo_valid
            & (~proc_done);
        proc_fifo_inject_push = 1'h0;
        proc_fifo_inject_data = 16'h0;
        proc_fifo_inject_eos = 1'h0;
      end :repeat_fsm_PASS_REPEAT_Output
    PASS_STOP: begin :repeat_fsm_PASS_STOP_Output
        ref_fifo_in_data = repsig_fifo_out_data;
        ref_fifo_in_eos = 1'h1;
        ref_fifo_push = repsig_stop & proc_fifo_valid & (~ref_fifo_full);
        proc_fifo_pop = repsig_fifo_valid & proc_stop & (~ref_fifo_full);
        repsig_fifo_pop = repsig_stop & proc_fifo_valid & (~ref_fifo_full);
        proc_fifo_inject_push = 1'h0;
        proc_fifo_inject_data = 16'h0;
        proc_fifo_inject_eos = 1'h0;
      end :repeat_fsm_PASS_STOP_Output
    START: begin :repeat_fsm_START_Output
        ref_fifo_in_data = 16'h0;
        ref_fifo_in_eos = 1'h0;
        ref_fifo_push = 1'h0;
        proc_fifo_pop = 1'h0;
        repsig_fifo_pop = 1'h0;
        proc_fifo_inject_push = 1'h0;
        proc_fifo_inject_data = 16'h0;
        proc_fifo_inject_eos = 1'h0;
      end :repeat_fsm_START_Output
    default: begin :repeat_fsm_default_Output
        ref_fifo_in_data = 16'h0;
        ref_fifo_in_eos = 1'h0;
        ref_fifo_push = 1'h0;
        proc_fifo_pop = 1'h0;
        repsig_fifo_pop = 1'h0;
        proc_fifo_inject_push = 1'h0;
        proc_fifo_inject_data = 16'h0;
        proc_fifo_inject_eos = 1'h0;
      end :repeat_fsm_default_Output
  endcase
end
reg_fifo_depth_0_w_17_afd_2 repsig_in_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(repsig_data_in),
  .flush(flush),
  .pop(repsig_fifo_pop),
  .push(repsig_data_in_valid),
  .rst_n(rst_n),
  .data_out(repsig_in_fifo_data_out),
  .empty(repsig_in_fifo_empty),
  .full(repsig_in_fifo_full)
);

reg_fifo_depth_2_w_17_afd_2 proc_in_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(proc_in_fifo_data_in),
  .flush(flush),
  .pop(proc_fifo_pop),
  .push(proc_fifo_push),
  .rst_n(rst_n),
  .data_out(proc_in_fifo_data_out),
  .empty(proc_in_fifo_empty),
  .full(proc_in_fifo_full)
);

reg_fifo_depth_0_w_17_afd_2 ref_out_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(ref_out_fifo_data_in),
  .flush(flush),
  .pop(ref_data_out_ready),
  .push(ref_fifo_push),
  .rst_n(rst_n),
  .data_out(ref_data_out),
  .empty(ref_out_fifo_empty),
  .full(ref_fifo_full)
);

endmodule   // Repeat

module RepeatSignalGenerator (
  input logic [16:0] base_data_in,
  input logic base_data_in_valid,
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic repsig_data_out_ready,
  input logic rst_n,
  input logic [15:0] stop_lvl,
  input logic tile_en,
  output logic base_data_in_ready,
  output logic [16:0] repsig_data_out,
  output logic repsig_data_out_valid
);

typedef enum logic[1:0] {
  DONE = 2'h0,
  PASS_REPEAT = 2'h1,
  PASS_STOP = 2'h2,
  START = 2'h3
} rsg_fsm_state;
logic already_pushed_repsig_eos_sticky;
logic already_pushed_repsig_eos_was_high;
logic [15:0] base_fifo_out_data;
logic base_fifo_out_eos;
logic base_fifo_pop;
logic base_fifo_valid;
logic [0:0][16:0] base_in_fifo_data_out;
logic base_in_fifo_empty;
logic base_in_fifo_full;
logic clr_already_pushed_repsig_eos;
logic gclk;
logic repsig_fifo_full;
logic [15:0] repsig_fifo_in_data;
logic repsig_fifo_in_eos;
logic repsig_fifo_push;
logic [0:0][16:0] repsig_out_fifo_data_in;
logic repsig_out_fifo_empty;
rsg_fsm_state rsg_fsm_current_state;
rsg_fsm_state rsg_fsm_next_state;
logic seen_root_eos_sticky;
logic seen_root_eos_was_high;
assign gclk = clk & tile_en;
assign {base_fifo_out_eos, base_fifo_out_data} = base_in_fifo_data_out;
assign base_data_in_ready = ~base_in_fifo_full;
assign base_fifo_valid = ~base_in_fifo_empty;
assign repsig_out_fifo_data_in = {repsig_fifo_in_eos, repsig_fifo_in_data};
assign repsig_data_out_valid = ~repsig_out_fifo_empty;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    seen_root_eos_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      seen_root_eos_was_high <= 1'h0;
    end
    else if (1'h0) begin
      seen_root_eos_was_high <= 1'h0;
    end
    else if ((base_fifo_out_data[9:8] == 2'h1) & base_fifo_out_eos & base_fifo_valid) begin
      seen_root_eos_was_high <= 1'h1;
    end
  end
end
assign seen_root_eos_sticky = ((base_fifo_out_data[9:8] == 2'h1) & base_fifo_out_eos & base_fifo_valid) |
    seen_root_eos_was_high;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    already_pushed_repsig_eos_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      already_pushed_repsig_eos_was_high <= 1'h0;
    end
    else if (clr_already_pushed_repsig_eos) begin
      already_pushed_repsig_eos_was_high <= 1'h0;
    end
    else if (repsig_fifo_push & (~repsig_fifo_full)) begin
      already_pushed_repsig_eos_was_high <= 1'h1;
    end
  end
end
assign already_pushed_repsig_eos_sticky = already_pushed_repsig_eos_was_high;

always_ff @(posedge clk, negedge rst_n) begin
  if (!rst_n) begin
    rsg_fsm_current_state <= START;
  end
  else if (clk_en) begin
    if (flush) begin
      rsg_fsm_current_state <= START;
    end
    else rsg_fsm_current_state <= rsg_fsm_next_state;
  end
end
always_comb begin
  rsg_fsm_next_state = rsg_fsm_current_state;
  unique case (rsg_fsm_current_state)
    DONE: rsg_fsm_next_state = START;
    PASS_REPEAT: begin
        if (base_fifo_out_eos & base_fifo_valid) begin
          rsg_fsm_next_state = PASS_STOP;
        end
        else rsg_fsm_next_state = PASS_REPEAT;
      end
    PASS_STOP: begin
        if (base_fifo_valid & base_fifo_out_eos & (base_fifo_out_data[9:8] == 2'h1) & (~repsig_fifo_full)) begin
          rsg_fsm_next_state = DONE;
        end
        else if (base_fifo_valid & (~base_fifo_out_eos)) begin
          rsg_fsm_next_state = PASS_REPEAT;
        end
        else rsg_fsm_next_state = PASS_STOP;
      end
    START: begin
        if (tile_en) begin
          rsg_fsm_next_state = PASS_REPEAT;
        end
        else rsg_fsm_next_state = START;
      end
    default: begin end
  endcase
end
always_comb begin
  unique case (rsg_fsm_current_state)
    DONE: begin :rsg_fsm_DONE_Output
        repsig_fifo_in_data = 16'h0;
        repsig_fifo_in_eos = 1'h0;
        repsig_fifo_push = 1'h0;
        base_fifo_pop = 1'h0;
        clr_already_pushed_repsig_eos = 1'h0;
      end :rsg_fsm_DONE_Output
    PASS_REPEAT: begin :rsg_fsm_PASS_REPEAT_Output
        repsig_fifo_in_data = 16'h1;
        repsig_fifo_in_eos = 1'h0;
        repsig_fifo_push = (~base_fifo_out_eos) & base_fifo_valid;
        clr_already_pushed_repsig_eos = 1'h1;
        base_fifo_pop = (~base_fifo_out_eos) & base_fifo_valid & (~repsig_fifo_full);
      end :rsg_fsm_PASS_REPEAT_Output
    PASS_STOP: begin :rsg_fsm_PASS_STOP_Output
        repsig_fifo_in_data = (base_fifo_out_data[9:8] == 2'h1) ? base_fifo_out_data: base_fifo_out_data;
        repsig_fifo_in_eos = 1'h1;
        repsig_fifo_push = base_fifo_out_eos & base_fifo_valid;
        clr_already_pushed_repsig_eos = 1'h0;
        base_fifo_pop = base_fifo_out_eos & base_fifo_valid & (~repsig_fifo_full);
      end :rsg_fsm_PASS_STOP_Output
    START: begin :rsg_fsm_START_Output
        repsig_fifo_in_data = 16'h0;
        repsig_fifo_in_eos = 1'h0;
        repsig_fifo_push = 1'h0;
        base_fifo_pop = 1'h0;
        clr_already_pushed_repsig_eos = 1'h0;
      end :rsg_fsm_START_Output
    default: begin end
  endcase
end
reg_fifo_depth_0_w_17_afd_2 base_in_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(base_data_in),
  .flush(flush),
  .pop(base_fifo_pop),
  .push(base_data_in_valid),
  .rst_n(rst_n),
  .data_out(base_in_fifo_data_out),
  .empty(base_in_fifo_empty),
  .full(base_in_fifo_full)
);

reg_fifo_depth_0_w_17_afd_2 repsig_out_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(repsig_out_fifo_data_in),
  .flush(flush),
  .pop(repsig_data_out_ready),
  .push(repsig_fifo_push),
  .rst_n(rst_n),
  .data_out(repsig_data_out),
  .empty(repsig_out_fifo_empty),
  .full(repsig_fifo_full)
);

endmodule   // RepeatSignalGenerator

module RepeatSignalGenerator_flat (
  input logic [15:0] RepeatSignalGenerator_inst_stop_lvl,
  input logic RepeatSignalGenerator_inst_tile_en,
  input logic [0:0] [16:0] base_data_in_f_,
  input logic base_data_in_valid_f_,
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic repsig_data_out_ready_f_,
  input logic rst_n,
  output logic base_data_in_ready_f_,
  output logic [0:0] [16:0] repsig_data_out_f_,
  output logic repsig_data_out_valid_f_
);

RepeatSignalGenerator RepeatSignalGenerator_inst (
  .base_data_in(base_data_in_f_),
  .base_data_in_valid(base_data_in_valid_f_),
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .repsig_data_out_ready(repsig_data_out_ready_f_),
  .rst_n(rst_n),
  .stop_lvl(RepeatSignalGenerator_inst_stop_lvl),
  .tile_en(RepeatSignalGenerator_inst_tile_en),
  .base_data_in_ready(base_data_in_ready_f_),
  .repsig_data_out(repsig_data_out_f_),
  .repsig_data_out_valid(repsig_data_out_valid_f_)
);

endmodule   // RepeatSignalGenerator_flat

module Repeat_flat (
  input logic Repeat_inst_root,
  input logic Repeat_inst_spacc_mode,
  input logic [15:0] Repeat_inst_stop_lvl,
  input logic Repeat_inst_tile_en,
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [0:0] [16:0] proc_data_in_f_,
  input logic proc_data_in_valid_f_,
  input logic ref_data_out_ready_f_,
  input logic [0:0] [16:0] repsig_data_in_f_,
  input logic repsig_data_in_valid_f_,
  input logic rst_n,
  output logic proc_data_in_ready_f_,
  output logic [0:0] [16:0] ref_data_out_f_,
  output logic ref_data_out_valid_f_,
  output logic repsig_data_in_ready_f_
);

Repeat Repeat_inst (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .proc_data_in(proc_data_in_f_),
  .proc_data_in_valid(proc_data_in_valid_f_),
  .ref_data_out_ready(ref_data_out_ready_f_),
  .repsig_data_in(repsig_data_in_f_),
  .repsig_data_in_valid(repsig_data_in_valid_f_),
  .root(Repeat_inst_root),
  .rst_n(rst_n),
  .spacc_mode(Repeat_inst_spacc_mode),
  .stop_lvl(Repeat_inst_stop_lvl),
  .tile_en(Repeat_inst_tile_en),
  .proc_data_in_ready(proc_data_in_ready_f_),
  .ref_data_out(ref_data_out_f_),
  .ref_data_out_valid(ref_data_out_valid_f_),
  .repsig_data_in_ready(repsig_data_in_ready_f_)
);

endmodule   // Repeat_flat

module crddrop (
  input logic clk,
  input logic clk_en,
  input logic [16:0] cmrg_coord_in_0,
  input logic cmrg_coord_in_0_valid,
  input logic [16:0] cmrg_coord_in_1,
  input logic cmrg_coord_in_1_valid,
  input logic cmrg_coord_out_0_ready,
  input logic cmrg_coord_out_1_ready,
  input logic cmrg_enable,
  input logic [15:0] cmrg_stop_lvl,
  input logic flush,
  input logic rst_n,
  input logic tile_en,
  output logic cmrg_coord_in_0_ready,
  output logic cmrg_coord_in_1_ready,
  output logic [16:0] cmrg_coord_out_0,
  output logic cmrg_coord_out_0_valid,
  output logic [16:0] cmrg_coord_out_1,
  output logic cmrg_coord_out_1_valid
);

typedef enum logic {
  PROCESS = 1'h0,
  START = 1'h1
} proc_seq_state;
logic base_data_seen;
logic base_done;
logic base_done_seen;
logic base_eos_seen;
logic base_infifo_empty;
logic base_infifo_full;
logic [15:0] base_infifo_in_data;
logic base_infifo_in_eos;
logic [16:0] base_infifo_in_packed;
logic base_infifo_in_valid;
logic [16:0] base_infifo_out_packed;
logic base_outfifo_empty;
logic base_outfifo_full;
logic [16:0] base_outfifo_in_packed;
logic [16:0] base_outfifo_out_packed;
logic both_done;
logic clr_pushed_data_lower;
logic clr_pushed_proc;
logic clr_pushed_stop_lvl;
logic cmrg_coord_in_0_eos;
logic cmrg_coord_in_1_eos;
logic [1:0] cmrg_fifo_pop;
logic [1:0] cmrg_fifo_push;
logic gclk;
logic proc_data_seen;
logic proc_done;
logic proc_infifo_empty;
logic proc_infifo_full;
logic [15:0] proc_infifo_in_data;
logic proc_infifo_in_eos;
logic [16:0] proc_infifo_in_packed;
logic proc_infifo_in_valid;
logic [16:0] proc_infifo_out_packed;
logic proc_outfifo_empty;
logic proc_outfifo_full;
logic [16:0] proc_outfifo_in_packed;
logic [16:0] proc_outfifo_out_packed;
proc_seq_state proc_seq_current_state;
proc_seq_state proc_seq_next_state;
logic pushed_data_sticky_sticky;
logic pushed_data_sticky_was_high;
logic pushed_proc_sticky;
logic pushed_proc_was_high;
logic pushed_stop_lvl_sticky;
logic pushed_stop_lvl_was_high;
logic pushing_done;
logic set_pushed_data_lower;
assign gclk = clk & tile_en;
assign cmrg_coord_in_0_eos = cmrg_coord_in_0[16];
assign cmrg_coord_in_1_eos = cmrg_coord_in_1[16];
assign base_infifo_in_packed[16] = cmrg_coord_in_0_eos;
assign base_infifo_in_packed[15:0] = cmrg_coord_in_0[15:0];
assign base_infifo_in_eos = base_infifo_out_packed[16];
assign base_infifo_in_data = base_infifo_out_packed[15:0];
assign base_infifo_in_valid = ~base_infifo_empty;
assign cmrg_coord_in_0_ready = ~base_infifo_full;
assign proc_infifo_in_packed[16] = cmrg_coord_in_1_eos;
assign proc_infifo_in_packed[15:0] = cmrg_coord_in_1[15:0];
assign proc_infifo_in_eos = proc_infifo_out_packed[16];
assign proc_infifo_in_data = proc_infifo_out_packed[15:0];
assign proc_infifo_in_valid = ~proc_infifo_empty;
assign cmrg_coord_in_1_ready = ~proc_infifo_full;
assign base_data_seen = base_infifo_in_valid & (~base_infifo_in_eos);
assign proc_data_seen = proc_infifo_in_valid & (~proc_infifo_in_eos);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    pushed_data_sticky_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      pushed_data_sticky_was_high <= 1'h0;
    end
    else if (clr_pushed_data_lower) begin
      pushed_data_sticky_was_high <= 1'h0;
    end
    else if (set_pushed_data_lower) begin
      pushed_data_sticky_was_high <= 1'h1;
    end
  end
end
assign pushed_data_sticky_sticky = pushed_data_sticky_was_high;
assign base_eos_seen = base_infifo_in_valid & base_infifo_in_eos & (base_infifo_in_data[9:8] == 2'h0);
assign base_done_seen = base_infifo_in_valid & base_infifo_in_eos & (base_infifo_in_data[9:8] == 2'h1);
assign base_done = base_infifo_in_valid & base_infifo_in_eos & (base_infifo_in_data[9:8] == 2'h1);
assign proc_done = proc_infifo_in_valid & proc_infifo_in_eos & (proc_infifo_in_data[9:8] == 2'h1);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    pushed_proc_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      pushed_proc_was_high <= 1'h0;
    end
    else if (clr_pushed_proc) begin
      pushed_proc_was_high <= 1'h0;
    end
    else if (cmrg_fifo_push[1]) begin
      pushed_proc_was_high <= 1'h1;
    end
  end
end
assign pushed_proc_sticky = pushed_proc_was_high;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    pushed_stop_lvl_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      pushed_stop_lvl_was_high <= 1'h0;
    end
    else if (clr_pushed_stop_lvl) begin
      pushed_stop_lvl_was_high <= 1'h0;
    end
    else if (cmrg_fifo_push[0] & base_infifo_in_valid & base_infifo_in_eos) begin
      pushed_stop_lvl_was_high <= 1'h1;
    end
  end
end
assign pushed_stop_lvl_sticky = pushed_stop_lvl_was_high;
assign both_done = base_infifo_in_valid & base_infifo_in_eos & proc_infifo_in_valid &
    proc_infifo_in_eos & (base_infifo_in_data[9:8] == 2'h1) &
    (proc_infifo_in_data[9:8] == 2'h1);
assign pushing_done = base_infifo_in_valid & base_infifo_in_eos & proc_infifo_in_valid &
    proc_infifo_in_eos & (base_infifo_in_data[9:8] == 2'h1) &
    (proc_infifo_in_data[9:8] == 2'h1) & (~base_outfifo_full) & (~proc_outfifo_full);
assign base_outfifo_in_packed[16] = base_infifo_in_eos;
assign base_outfifo_in_packed[15:0] = base_infifo_in_data;
assign cmrg_coord_out_0[16] = base_outfifo_out_packed[16];
assign cmrg_coord_out_0[15:0] = base_outfifo_out_packed[15:0];
assign cmrg_coord_out_0_valid = ~base_outfifo_empty;
assign proc_outfifo_in_packed[16] = proc_infifo_in_eos;
assign proc_outfifo_in_packed[15:0] = proc_infifo_in_data;
assign cmrg_coord_out_1[16] = proc_outfifo_out_packed[16];
assign cmrg_coord_out_1[15:0] = proc_outfifo_out_packed[15:0];
assign cmrg_coord_out_1_valid = ~proc_outfifo_empty;

always_ff @(posedge clk, negedge rst_n) begin
  if (!rst_n) begin
    proc_seq_current_state <= START;
  end
  else if (clk_en) begin
    if (flush) begin
      proc_seq_current_state <= START;
    end
    else proc_seq_current_state <= proc_seq_next_state;
  end
end
always_comb begin
  proc_seq_next_state = proc_seq_current_state;
  unique case (proc_seq_current_state)
    PROCESS: proc_seq_next_state = PROCESS;
    START: begin
        if (tile_en) begin
          proc_seq_next_state = PROCESS;
        end
        else proc_seq_next_state = START;
      end
    default: begin end
  endcase
end
always_comb begin
  unique case (proc_seq_current_state)
    PROCESS: begin :proc_seq_PROCESS_Output
        cmrg_fifo_pop[0] = base_done ? proc_done & (~base_outfifo_full) & (~proc_outfifo_full):
            (base_infifo_in_valid & (~base_infifo_in_eos)) ? ~base_outfifo_full:
            (base_infifo_in_valid & base_infifo_in_eos) ? (proc_done | (proc_infifo_in_valid
            & (~proc_infifo_in_eos))) & (~base_outfifo_full) & (~proc_outfifo_full): 1'h0;
        cmrg_fifo_pop[1] = proc_done ? base_done & (~base_outfifo_full) & (~proc_outfifo_full):
            (base_infifo_in_valid & base_infifo_in_eos & proc_infifo_in_valid &
            (~proc_infifo_in_eos)) ? (~base_outfifo_full) & ((~proc_outfifo_full) |
            (~pushed_data_sticky_sticky)): (proc_infifo_in_valid & proc_infifo_in_eos) ?
            ~proc_outfifo_full: 1'h0;
        cmrg_fifo_push[0] = base_done ? proc_done: (base_infifo_in_valid & (~base_infifo_in_eos)) ?
            ~base_outfifo_full: (base_infifo_in_valid & base_infifo_in_eos) ? (proc_done |
            (proc_infifo_in_valid & (~proc_infifo_in_eos) & pushed_data_sticky_sticky)) &
            (~base_outfifo_full) & (~proc_outfifo_full): 1'h0;
        cmrg_fifo_push[1] = proc_done ? base_done: (base_infifo_in_valid & base_infifo_in_eos &
            proc_infifo_in_valid & (~proc_infifo_in_eos)) ? (~base_outfifo_full) &
            (~proc_outfifo_full) & pushed_data_sticky_sticky: (proc_infifo_in_valid &
            proc_infifo_in_eos) ? ~proc_outfifo_full: 1'h0;
        clr_pushed_proc = 1'h0;
        clr_pushed_stop_lvl = 1'h0;
        set_pushed_data_lower = base_infifo_in_valid & (~base_infifo_in_eos) & (~base_outfifo_full);
        clr_pushed_data_lower = base_done | (base_infifo_in_valid & base_infifo_in_eos & proc_infifo_in_valid &
            (~proc_infifo_in_eos) & (~base_outfifo_full) & (~proc_outfifo_full));
      end :proc_seq_PROCESS_Output
    START: begin :proc_seq_START_Output
        cmrg_fifo_pop[0] = 1'h0;
        cmrg_fifo_pop[1] = 1'h0;
        cmrg_fifo_push[0] = 1'h0;
        cmrg_fifo_push[1] = 1'h0;
        clr_pushed_proc = 1'h1;
        clr_pushed_stop_lvl = 1'h1;
        set_pushed_data_lower = 1'h0;
        clr_pushed_data_lower = 1'h1;
      end :proc_seq_START_Output
    default: begin end
  endcase
end
reg_fifo_depth_0_w_17_afd_2 base_infifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(base_infifo_in_packed),
  .flush(flush),
  .pop(cmrg_fifo_pop[0]),
  .push(cmrg_coord_in_0_valid),
  .rst_n(rst_n),
  .data_out(base_infifo_out_packed),
  .empty(base_infifo_empty),
  .full(base_infifo_full)
);

reg_fifo_depth_0_w_17_afd_2 proc_infifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(proc_infifo_in_packed),
  .flush(flush),
  .pop(cmrg_fifo_pop[1]),
  .push(cmrg_coord_in_1_valid),
  .rst_n(rst_n),
  .data_out(proc_infifo_out_packed),
  .empty(proc_infifo_empty),
  .full(proc_infifo_full)
);

reg_fifo_depth_0_w_17_afd_2 base_outfifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(base_outfifo_in_packed),
  .flush(flush),
  .pop(cmrg_coord_out_0_ready),
  .push(cmrg_fifo_push[0]),
  .rst_n(rst_n),
  .data_out(base_outfifo_out_packed),
  .empty(base_outfifo_empty),
  .full(base_outfifo_full)
);

reg_fifo_depth_0_w_17_afd_2 proc_outfifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(proc_outfifo_in_packed),
  .flush(flush),
  .pop(cmrg_coord_out_1_ready),
  .push(cmrg_fifo_push[1]),
  .rst_n(rst_n),
  .data_out(proc_outfifo_out_packed),
  .empty(proc_outfifo_empty),
  .full(proc_outfifo_full)
);

endmodule   // crddrop

module crddrop_flat (
  input logic clk,
  input logic clk_en,
  input logic [0:0] [16:0] cmrg_coord_in_0_f_,
  input logic cmrg_coord_in_0_valid_f_,
  input logic [0:0] [16:0] cmrg_coord_in_1_f_,
  input logic cmrg_coord_in_1_valid_f_,
  input logic cmrg_coord_out_0_ready_f_,
  input logic cmrg_coord_out_1_ready_f_,
  input logic crddrop_inst_cmrg_enable,
  input logic [15:0] crddrop_inst_cmrg_stop_lvl,
  input logic crddrop_inst_tile_en,
  input logic flush,
  input logic rst_n,
  output logic cmrg_coord_in_0_ready_f_,
  output logic cmrg_coord_in_1_ready_f_,
  output logic [0:0] [16:0] cmrg_coord_out_0_f_,
  output logic cmrg_coord_out_0_valid_f_,
  output logic [0:0] [16:0] cmrg_coord_out_1_f_,
  output logic cmrg_coord_out_1_valid_f_
);

crddrop crddrop_inst (
  .clk(clk),
  .clk_en(clk_en),
  .cmrg_coord_in_0(cmrg_coord_in_0_f_),
  .cmrg_coord_in_0_valid(cmrg_coord_in_0_valid_f_),
  .cmrg_coord_in_1(cmrg_coord_in_1_f_),
  .cmrg_coord_in_1_valid(cmrg_coord_in_1_valid_f_),
  .cmrg_coord_out_0_ready(cmrg_coord_out_0_ready_f_),
  .cmrg_coord_out_1_ready(cmrg_coord_out_1_ready_f_),
  .cmrg_enable(crddrop_inst_cmrg_enable),
  .cmrg_stop_lvl(crddrop_inst_cmrg_stop_lvl),
  .flush(flush),
  .rst_n(rst_n),
  .tile_en(crddrop_inst_tile_en),
  .cmrg_coord_in_0_ready(cmrg_coord_in_0_ready_f_),
  .cmrg_coord_in_1_ready(cmrg_coord_in_1_ready_f_),
  .cmrg_coord_out_0(cmrg_coord_out_0_f_),
  .cmrg_coord_out_0_valid(cmrg_coord_out_0_valid_f_),
  .cmrg_coord_out_1(cmrg_coord_out_1_f_),
  .cmrg_coord_out_1_valid(cmrg_coord_out_1_valid_f_)
);

endmodule   // crddrop_flat

module crdhold (
  input logic clk,
  input logic clk_en,
  input logic [16:0] cmrg_coord_in_0,
  input logic cmrg_coord_in_0_valid,
  input logic [16:0] cmrg_coord_in_1,
  input logic cmrg_coord_in_1_valid,
  input logic cmrg_coord_out_0_ready,
  input logic cmrg_coord_out_1_ready,
  input logic cmrg_enable,
  input logic [15:0] cmrg_stop_lvl,
  input logic flush,
  input logic rst_n,
  input logic tile_en,
  output logic cmrg_coord_in_0_ready,
  output logic cmrg_coord_in_1_ready,
  output logic [16:0] cmrg_coord_out_0,
  output logic cmrg_coord_out_0_valid,
  output logic [16:0] cmrg_coord_out_1,
  output logic cmrg_coord_out_1_valid
);

typedef enum logic[1:0] {
  DATA_SEEN = 2'h0,
  DONE = 2'h1,
  START = 2'h2
} proc_seq_state;
logic base_data_seen;
logic base_done_seen;
logic base_eos_seen;
logic base_infifo_empty;
logic base_infifo_full;
logic [15:0] base_infifo_in_data;
logic base_infifo_in_eos;
logic [16:0] base_infifo_in_packed;
logic base_infifo_in_valid;
logic [16:0] base_infifo_out_packed;
logic base_outfifo_empty;
logic base_outfifo_full;
logic [16:0] base_outfifo_in_packed;
logic [16:0] base_outfifo_out_packed;
logic both_done;
logic clr_pushed_base;
logic clr_pushed_proc;
logic cmrg_coord_in_0_eos;
logic cmrg_coord_in_1_eos;
logic [1:0] cmrg_fifo_pop;
logic [1:0] cmrg_fifo_push;
logic [15:0] data_to_fifo;
logic eos_to_fifo;
logic gclk;
logic [15:0] hold_reg;
logic proc_data_seen;
logic proc_done_seen;
logic proc_eos_seen;
logic proc_infifo_empty;
logic proc_infifo_full;
logic [15:0] proc_infifo_in_data;
logic proc_infifo_in_eos;
logic [16:0] proc_infifo_in_packed;
logic proc_infifo_in_valid;
logic [16:0] proc_infifo_out_packed;
logic proc_outfifo_empty;
logic proc_outfifo_full;
logic [16:0] proc_outfifo_in_packed;
logic [16:0] proc_outfifo_out_packed;
proc_seq_state proc_seq_current_state;
proc_seq_state proc_seq_next_state;
logic pushed_base_sticky;
logic pushed_base_was_high;
logic pushed_proc_sticky;
logic pushed_proc_was_high;
logic pushing_done;
logic reg_clr;
logic reg_hold;
assign gclk = clk & tile_en;
assign cmrg_coord_in_0_eos = cmrg_coord_in_0[16];
assign cmrg_coord_in_1_eos = cmrg_coord_in_1[16];
assign base_infifo_in_packed[16] = cmrg_coord_in_0_eos;
assign base_infifo_in_packed[15:0] = cmrg_coord_in_0[15:0];
assign base_infifo_in_eos = base_infifo_out_packed[16];
assign base_infifo_in_data = base_infifo_out_packed[15:0];
assign base_infifo_in_valid = ~base_infifo_empty;
assign cmrg_coord_in_0_ready = ~base_infifo_full;
assign proc_infifo_in_packed[16] = cmrg_coord_in_1_eos;
assign proc_infifo_in_packed[15:0] = cmrg_coord_in_1[15:0];
assign proc_infifo_in_eos = proc_infifo_out_packed[16];
assign proc_infifo_in_data = proc_infifo_out_packed[15:0];
assign proc_infifo_in_valid = ~proc_infifo_empty;
assign cmrg_coord_in_1_ready = ~proc_infifo_full;
assign base_data_seen = base_infifo_in_valid & (~base_infifo_in_eos);
assign proc_data_seen = proc_infifo_in_valid & (~proc_infifo_in_eos);
assign base_eos_seen = base_infifo_in_valid & base_infifo_in_eos & (base_infifo_in_data[9:8] == 2'h0);
assign proc_eos_seen = proc_infifo_in_valid & proc_infifo_in_eos & (proc_infifo_in_data[9:8] == 2'h0);
assign base_done_seen = base_infifo_in_valid & base_infifo_in_eos & (base_infifo_in_data[9:8] == 2'h1);
assign proc_done_seen = proc_infifo_in_valid & proc_infifo_in_eos & (proc_infifo_in_data[9:8] == 2'h1);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    pushed_proc_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      pushed_proc_was_high <= 1'h0;
    end
    else if (clr_pushed_proc) begin
      pushed_proc_was_high <= 1'h0;
    end
    else if (cmrg_fifo_push[1]) begin
      pushed_proc_was_high <= 1'h1;
    end
  end
end
assign pushed_proc_sticky = pushed_proc_was_high;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    pushed_base_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      pushed_base_was_high <= 1'h0;
    end
    else if (clr_pushed_base) begin
      pushed_base_was_high <= 1'h0;
    end
    else if (cmrg_fifo_push[0]) begin
      pushed_base_was_high <= 1'h1;
    end
  end
end
assign pushed_base_sticky = pushed_base_was_high;
assign both_done = base_infifo_in_valid & base_infifo_in_eos & proc_infifo_in_valid &
    proc_infifo_in_eos & (base_infifo_in_data[9:8] == 2'h1) &
    (proc_infifo_in_data[9:8] == 2'h1);
assign pushing_done = base_infifo_in_valid & base_infifo_in_eos & proc_infifo_in_valid &
    proc_infifo_in_eos & (base_infifo_in_data[9:8] == 2'h1) &
    (proc_infifo_in_data[9:8] == 2'h1) & (~base_outfifo_full) & (~proc_outfifo_full);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    hold_reg <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      hold_reg <= 16'h0;
    end
    else if (reg_clr) begin
      hold_reg <= 16'h0;
    end
    else if (reg_hold) begin
      hold_reg <= proc_infifo_in_data;
    end
  end
end
assign base_outfifo_in_packed[16] = base_infifo_in_eos;
assign base_outfifo_in_packed[15:0] = base_infifo_in_data;
assign cmrg_coord_out_0[16] = base_outfifo_out_packed[16];
assign cmrg_coord_out_0[15:0] = base_outfifo_out_packed[15:0];
assign cmrg_coord_out_0_valid = ~base_outfifo_empty;
assign proc_outfifo_in_packed[16] = eos_to_fifo;
assign proc_outfifo_in_packed[15:0] = data_to_fifo;
assign cmrg_coord_out_1[16] = proc_outfifo_out_packed[16];
assign cmrg_coord_out_1[15:0] = proc_outfifo_out_packed[15:0];
assign cmrg_coord_out_1_valid = ~proc_outfifo_empty;

always_ff @(posedge clk, negedge rst_n) begin
  if (!rst_n) begin
    proc_seq_current_state <= START;
  end
  else if (clk_en) begin
    if (flush) begin
      proc_seq_current_state <= START;
    end
    else proc_seq_current_state <= proc_seq_next_state;
  end
end
always_comb begin
  proc_seq_next_state = proc_seq_current_state;
  unique case (proc_seq_current_state)
    DATA_SEEN: begin
        if (both_done) begin
          proc_seq_next_state = DONE;
        end
        else proc_seq_next_state = DATA_SEEN;
      end
    DONE: begin
        if ((~base_outfifo_full) & (~proc_outfifo_full)) begin
          proc_seq_next_state = START;
        end
      end
    START: begin
        if (tile_en) begin
          proc_seq_next_state = DATA_SEEN;
        end
        else proc_seq_next_state = START;
      end
    default: proc_seq_next_state = proc_seq_current_state;
  endcase
end
always_comb begin
  unique case (proc_seq_current_state)
    DATA_SEEN: begin :proc_seq_DATA_SEEN_Output
        cmrg_fifo_pop[0] = (base_eos_seen ? 1'h1: base_infifo_in_valid & (~base_infifo_in_eos) &
            proc_infifo_in_valid & (~proc_infifo_in_eos)) & (~base_outfifo_full) &
            (~proc_outfifo_full) & (~base_done_seen);
        cmrg_fifo_pop[1] = (proc_eos_seen ? 1'h1: base_eos_seen & (~base_outfifo_full) &
            (~proc_outfifo_full)) & (~proc_done_seen);
        cmrg_fifo_push[0] = (base_eos_seen ? 1'h1: base_infifo_in_valid & (~base_infifo_in_eos) &
            proc_infifo_in_valid & (~proc_infifo_in_eos)) & (~base_outfifo_full) &
            (~proc_outfifo_full) & (~base_done_seen);
        cmrg_fifo_push[1] = (base_eos_seen ? 1'h1: base_infifo_in_valid & (~base_infifo_in_eos) &
            proc_infifo_in_valid & (~proc_infifo_in_eos)) & (~base_outfifo_full) &
            (~proc_outfifo_full) & (~base_done_seen);
        data_to_fifo = base_infifo_in_eos ? base_infifo_in_data: proc_infifo_in_data;
        eos_to_fifo = base_infifo_in_eos;
        clr_pushed_proc = 1'h1;
        clr_pushed_base = 1'h1;
        reg_clr = 1'h1;
        reg_hold = 1'h0;
      end :proc_seq_DATA_SEEN_Output
    DONE: begin :proc_seq_DONE_Output
        cmrg_fifo_pop[0] = (~proc_outfifo_full) & (~base_outfifo_full);
        cmrg_fifo_pop[1] = (~proc_outfifo_full) & (~base_outfifo_full);
        cmrg_fifo_push[0] = (~proc_outfifo_full) & (~base_outfifo_full);
        cmrg_fifo_push[1] = (~proc_outfifo_full) & (~base_outfifo_full);
        data_to_fifo = base_infifo_in_data;
        eos_to_fifo = 1'h1;
        clr_pushed_proc = 1'h1;
        clr_pushed_base = 1'h1;
        reg_clr = 1'h1;
        reg_hold = 1'h0;
      end :proc_seq_DONE_Output
    START: begin :proc_seq_START_Output
        cmrg_fifo_pop[0] = 1'h0;
        cmrg_fifo_pop[1] = 1'h0;
        cmrg_fifo_push[0] = 1'h0;
        cmrg_fifo_push[1] = 1'h0;
        data_to_fifo = 16'h0;
        eos_to_fifo = 1'h0;
        clr_pushed_proc = 1'h1;
        clr_pushed_base = 1'h1;
        reg_clr = 1'h0;
        reg_hold = 1'h0;
      end :proc_seq_START_Output
    default: begin :proc_seq_default_Output
        cmrg_fifo_pop[0] = 1'h0;
        cmrg_fifo_pop[1] = 1'h0;
        cmrg_fifo_push[0] = 1'h0;
        cmrg_fifo_push[1] = 1'h0;
        data_to_fifo = 16'h0;
        eos_to_fifo = 1'h0;
        clr_pushed_proc = 1'h1;
        clr_pushed_base = 1'h1;
        reg_clr = 1'h0;
        reg_hold = 1'h0;
      end :proc_seq_default_Output
  endcase
end
reg_fifo_depth_0_w_17_afd_2 base_infifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(base_infifo_in_packed),
  .flush(flush),
  .pop(cmrg_fifo_pop[0]),
  .push(cmrg_coord_in_0_valid),
  .rst_n(rst_n),
  .data_out(base_infifo_out_packed),
  .empty(base_infifo_empty),
  .full(base_infifo_full)
);

reg_fifo_depth_0_w_17_afd_2 proc_infifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(proc_infifo_in_packed),
  .flush(flush),
  .pop(cmrg_fifo_pop[1]),
  .push(cmrg_coord_in_1_valid),
  .rst_n(rst_n),
  .data_out(proc_infifo_out_packed),
  .empty(proc_infifo_empty),
  .full(proc_infifo_full)
);

reg_fifo_depth_0_w_17_afd_2 base_outfifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(base_outfifo_in_packed),
  .flush(flush),
  .pop(cmrg_coord_out_0_ready),
  .push(cmrg_fifo_push[0]),
  .rst_n(rst_n),
  .data_out(base_outfifo_out_packed),
  .empty(base_outfifo_empty),
  .full(base_outfifo_full)
);

reg_fifo_depth_0_w_17_afd_2 proc_outfifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(proc_outfifo_in_packed),
  .flush(flush),
  .pop(cmrg_coord_out_1_ready),
  .push(cmrg_fifo_push[1]),
  .rst_n(rst_n),
  .data_out(proc_outfifo_out_packed),
  .empty(proc_outfifo_empty),
  .full(proc_outfifo_full)
);

endmodule   // crdhold

module crdhold_flat (
  input logic clk,
  input logic clk_en,
  input logic [0:0] [16:0] cmrg_coord_in_0_f_,
  input logic cmrg_coord_in_0_valid_f_,
  input logic [0:0] [16:0] cmrg_coord_in_1_f_,
  input logic cmrg_coord_in_1_valid_f_,
  input logic cmrg_coord_out_0_ready_f_,
  input logic cmrg_coord_out_1_ready_f_,
  input logic crdhold_inst_cmrg_enable,
  input logic [15:0] crdhold_inst_cmrg_stop_lvl,
  input logic crdhold_inst_tile_en,
  input logic flush,
  input logic rst_n,
  output logic cmrg_coord_in_0_ready_f_,
  output logic cmrg_coord_in_1_ready_f_,
  output logic [0:0] [16:0] cmrg_coord_out_0_f_,
  output logic cmrg_coord_out_0_valid_f_,
  output logic [0:0] [16:0] cmrg_coord_out_1_f_,
  output logic cmrg_coord_out_1_valid_f_
);

crdhold crdhold_inst (
  .clk(clk),
  .clk_en(clk_en),
  .cmrg_coord_in_0(cmrg_coord_in_0_f_),
  .cmrg_coord_in_0_valid(cmrg_coord_in_0_valid_f_),
  .cmrg_coord_in_1(cmrg_coord_in_1_f_),
  .cmrg_coord_in_1_valid(cmrg_coord_in_1_valid_f_),
  .cmrg_coord_out_0_ready(cmrg_coord_out_0_ready_f_),
  .cmrg_coord_out_1_ready(cmrg_coord_out_1_ready_f_),
  .cmrg_enable(crdhold_inst_cmrg_enable),
  .cmrg_stop_lvl(crdhold_inst_cmrg_stop_lvl),
  .flush(flush),
  .rst_n(rst_n),
  .tile_en(crdhold_inst_tile_en),
  .cmrg_coord_in_0_ready(cmrg_coord_in_0_ready_f_),
  .cmrg_coord_in_1_ready(cmrg_coord_in_1_ready_f_),
  .cmrg_coord_out_0(cmrg_coord_out_0_f_),
  .cmrg_coord_out_0_valid(cmrg_coord_out_0_valid_f_),
  .cmrg_coord_out_1(cmrg_coord_out_1_f_),
  .cmrg_coord_out_1_valid(cmrg_coord_out_1_valid_f_)
);

endmodule   // crdhold_flat

module intersect_unit (
  input logic clk,
  input logic clk_en,
  input logic [16:0] coord_in_0,
  input logic coord_in_0_valid,
  input logic [16:0] coord_in_1,
  input logic coord_in_1_valid,
  input logic coord_out_ready,
  input logic flush,
  input logic joiner_op,
  input logic [16:0] pos_in_0,
  input logic pos_in_0_valid,
  input logic [16:0] pos_in_1,
  input logic pos_in_1_valid,
  input logic pos_out_0_ready,
  input logic pos_out_1_ready,
  input logic rst_n,
  input logic tile_en,
  output logic coord_in_0_ready,
  output logic coord_in_1_ready,
  output logic [16:0] coord_out,
  output logic coord_out_valid,
  output logic pos_in_0_ready,
  output logic pos_in_1_ready,
  output logic [16:0] pos_out_0,
  output logic pos_out_0_valid,
  output logic [16:0] pos_out_1,
  output logic pos_out_1_valid
);

typedef enum logic[2:0] {
  ALIGN = 3'h0,
  DONE = 3'h1,
  DRAIN = 3'h2,
  IDLE = 3'h3,
  ITER = 3'h4,
  UNION = 3'h5
} intersect_seq_state;
logic all_valid;
logic all_valid_join;
logic any_eos;
logic [1:0] clr_eos_sticky;
logic [16:0] coord_fifo_in_packed;
logic [16:0] coord_fifo_out_packed;
logic coord_in_0_fifo_eos_in;
logic [16:0] coord_in_0_fifo_in;
logic coord_in_0_fifo_valid_in;
logic coord_in_1_fifo_eos_in;
logic [16:0] coord_in_1_fifo_in;
logic coord_in_1_fifo_valid_in;
logic coord_in_fifo_0_empty;
logic coord_in_fifo_0_full;
logic coord_in_fifo_1_empty;
logic coord_in_fifo_1_full;
logic [15:0] coord_to_fifo;
logic coord_to_fifo_eos;
logic coordinate_fifo_empty;
logic coordinate_fifo_full;
logic [1:0] eos_in_sticky;
logic eos_sticky_0_sticky;
logic eos_sticky_0_was_high;
logic eos_sticky_1_sticky;
logic eos_sticky_1_was_high;
logic [2:0] fifo_full;
logic fifo_push;
logic gclk;
logic [1:0] inc_pos_cnt;
intersect_seq_state intersect_seq_current_state;
intersect_seq_state intersect_seq_next_state;
logic [15:0] maybe;
logic pos0_fifo_empty;
logic pos0_fifo_full;
logic [16:0] pos0_fifo_in_packed;
logic [16:0] pos0_fifo_out_packed;
logic pos1_fifo_empty;
logic pos1_fifo_full;
logic [16:0] pos1_fifo_in_packed;
logic [16:0] pos1_fifo_out_packed;
logic [1:0][15:0] pos_cnt;
logic pos_in_0_fifo_eos_in;
logic [16:0] pos_in_0_fifo_in;
logic pos_in_0_fifo_valid_in;
logic pos_in_1_fifo_eos_in;
logic [16:0] pos_in_1_fifo_in;
logic pos_in_1_fifo_valid_in;
logic pos_in_fifo_0_empty;
logic pos_in_fifo_0_full;
logic pos_in_fifo_1_empty;
logic pos_in_fifo_1_full;
logic [1:0][15:0] pos_to_fifo;
logic [1:0] pos_to_fifo_eos;
logic [1:0] rst_pos_cnt;
assign gclk = clk & tile_en;
assign coord_in_0_fifo_eos_in = coord_in_0_fifo_in[16];
assign coord_in_0_ready = ~coord_in_fifo_0_full;
assign coord_in_0_fifo_valid_in = ~coord_in_fifo_0_empty;
assign pos_in_0_fifo_eos_in = pos_in_0_fifo_in[16];
assign pos_in_0_ready = ~pos_in_fifo_0_full;
assign pos_in_0_fifo_valid_in = ~pos_in_fifo_0_empty;
assign coord_in_1_fifo_eos_in = coord_in_1_fifo_in[16];
assign coord_in_1_ready = ~coord_in_fifo_1_full;
assign coord_in_1_fifo_valid_in = ~coord_in_fifo_1_empty;
assign pos_in_1_fifo_eos_in = pos_in_1_fifo_in[16];
assign pos_in_1_ready = ~pos_in_fifo_1_full;
assign pos_in_1_fifo_valid_in = ~pos_in_fifo_1_empty;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    eos_sticky_0_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      eos_sticky_0_was_high <= 1'h0;
    end
    else if (clr_eos_sticky[0]) begin
      eos_sticky_0_was_high <= 1'h0;
    end
    else if (coord_in_0_fifo_eos_in & coord_in_0_fifo_valid_in & pos_in_0_fifo_eos_in & pos_in_0_fifo_valid_in) begin
      eos_sticky_0_was_high <= 1'h1;
    end
  end
end
assign eos_sticky_0_sticky = (coord_in_0_fifo_eos_in & coord_in_0_fifo_valid_in & pos_in_0_fifo_eos_in &
    pos_in_0_fifo_valid_in) | eos_sticky_0_was_high;
assign eos_in_sticky[0] = eos_sticky_0_sticky;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    eos_sticky_1_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      eos_sticky_1_was_high <= 1'h0;
    end
    else if (clr_eos_sticky[1]) begin
      eos_sticky_1_was_high <= 1'h0;
    end
    else if (coord_in_1_fifo_eos_in & coord_in_1_fifo_valid_in & pos_in_1_fifo_eos_in & pos_in_1_fifo_valid_in) begin
      eos_sticky_1_was_high <= 1'h1;
    end
  end
end
assign eos_sticky_1_sticky = (coord_in_1_fifo_eos_in & coord_in_1_fifo_valid_in & pos_in_1_fifo_eos_in &
    pos_in_1_fifo_valid_in) | eos_sticky_1_was_high;
assign eos_in_sticky[1] = eos_sticky_1_sticky;
assign all_valid = (&{coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in,
    pos_in_1_fifo_valid_in}) & (~any_eos);
assign all_valid_join = &{coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in,
    pos_in_1_fifo_valid_in};
assign any_eos = |({coord_in_0_fifo_eos_in, coord_in_1_fifo_eos_in, pos_in_0_fifo_eos_in,
    pos_in_1_fifo_eos_in} & {coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in,
    pos_in_0_fifo_valid_in, pos_in_1_fifo_valid_in});
assign maybe = {6'h0, 2'h2, 8'h0};

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    pos_cnt[0] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      pos_cnt[0] <= 16'h0;
    end
    else if (rst_pos_cnt[0]) begin
      pos_cnt[0] <= 16'h0;
    end
    else if (inc_pos_cnt[0]) begin
      pos_cnt[0] <= pos_cnt[0] + 16'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    pos_cnt[1] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      pos_cnt[1] <= 16'h0;
    end
    else if (rst_pos_cnt[1]) begin
      pos_cnt[1] <= 16'h0;
    end
    else if (inc_pos_cnt[1]) begin
      pos_cnt[1] <= pos_cnt[1] + 16'h1;
    end
  end
end
assign coord_fifo_in_packed[16] = coord_to_fifo_eos;
assign coord_fifo_in_packed[15:0] = coord_to_fifo;
assign coord_out[16] = coord_fifo_out_packed[16];
assign coord_out[15:0] = coord_fifo_out_packed[15:0];
assign pos0_fifo_in_packed[16] = pos_to_fifo_eos[0];
assign pos0_fifo_in_packed[15:0] = pos_to_fifo[0];
assign pos_out_0[16] = pos0_fifo_out_packed[16];
assign pos_out_0[15:0] = pos0_fifo_out_packed[15:0];
assign pos1_fifo_in_packed[16] = pos_to_fifo_eos[1];
assign pos1_fifo_in_packed[15:0] = pos_to_fifo[1];
assign pos_out_1[16] = pos1_fifo_out_packed[16];
assign pos_out_1[15:0] = pos1_fifo_out_packed[15:0];
assign fifo_full[0] = coordinate_fifo_full;
assign fifo_full[1] = pos0_fifo_full;
assign fifo_full[2] = pos1_fifo_full;
assign coord_out_valid = ~coordinate_fifo_empty;
assign pos_out_0_valid = ~pos0_fifo_empty;
assign pos_out_1_valid = ~pos1_fifo_empty;

always_ff @(posedge clk, negedge rst_n) begin
  if (!rst_n) begin
    intersect_seq_current_state <= IDLE;
  end
  else if (clk_en) begin
    if (flush) begin
      intersect_seq_current_state <= IDLE;
    end
    else intersect_seq_current_state <= intersect_seq_next_state;
  end
end
always_comb begin
  intersect_seq_next_state = intersect_seq_current_state;
  unique case (intersect_seq_current_state)
    ALIGN: begin
        if (&eos_in_sticky) begin
          intersect_seq_next_state = DRAIN;
        end
        else intersect_seq_next_state = ALIGN;
      end
    DONE: intersect_seq_next_state = IDLE;
    DRAIN: begin
        if ((~(&({coord_in_0_fifo_eos_in, coord_in_1_fifo_eos_in, pos_in_0_fifo_eos_in, pos_in_1_fifo_eos_in} & {coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in, pos_in_1_fifo_valid_in}))) & (&{coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in, pos_in_1_fifo_valid_in})) begin
          intersect_seq_next_state = DONE;
        end
        else intersect_seq_next_state = DRAIN;
      end
    IDLE: begin
        if (all_valid_join & (joiner_op == 1'h1) & tile_en) begin
          intersect_seq_next_state = UNION;
        end
        else if (any_eos & (joiner_op == 1'h0) & tile_en) begin
          intersect_seq_next_state = ALIGN;
        end
        else if (all_valid & (joiner_op == 1'h0) & tile_en) begin
          intersect_seq_next_state = ITER;
        end
        else intersect_seq_next_state = IDLE;
      end
    ITER: begin
        if (any_eos) begin
          intersect_seq_next_state = ALIGN;
        end
        else intersect_seq_next_state = ITER;
      end
    UNION: begin
        if (&eos_in_sticky) begin
          intersect_seq_next_state = DRAIN;
        end
        else intersect_seq_next_state = UNION;
      end
    default: intersect_seq_next_state = intersect_seq_current_state;
  endcase
end
always_comb begin
  unique case (intersect_seq_current_state)
    ALIGN: begin :intersect_seq_ALIGN_Output
        inc_pos_cnt[0] = (~eos_in_sticky[0]) & coord_in_0_fifo_valid_in & pos_in_0_fifo_valid_in;
        inc_pos_cnt[1] = (~eos_in_sticky[1]) & coord_in_1_fifo_valid_in & pos_in_1_fifo_valid_in;
        rst_pos_cnt[0] = 1'h0;
        rst_pos_cnt[1] = 1'h0;
        fifo_push = 1'h0;
        clr_eos_sticky[0] = 1'h0;
        clr_eos_sticky[1] = 1'h0;
        coord_to_fifo = 16'h0;
        pos_to_fifo[0] = 16'h0;
        pos_to_fifo[1] = 16'h0;
        coord_to_fifo_eos = 1'h0;
        pos_to_fifo_eos[0] = 1'h0;
        pos_to_fifo_eos[1] = 1'h0;
      end :intersect_seq_ALIGN_Output
    DONE: begin :intersect_seq_DONE_Output
        inc_pos_cnt[0] = 1'h0;
        inc_pos_cnt[1] = 1'h0;
        rst_pos_cnt[0] = 1'h1;
        rst_pos_cnt[1] = 1'h1;
        fifo_push = 1'h0;
        clr_eos_sticky[0] = 1'h1;
        clr_eos_sticky[1] = 1'h1;
        coord_to_fifo = 16'h0;
        pos_to_fifo[0] = 16'h0;
        pos_to_fifo[1] = 16'h0;
        coord_to_fifo_eos = 1'h0;
        pos_to_fifo_eos[0] = 1'h0;
        pos_to_fifo_eos[1] = 1'h0;
      end :intersect_seq_DONE_Output
    DRAIN: begin :intersect_seq_DRAIN_Output
        inc_pos_cnt[0] = (~(|fifo_full)) & (&({coord_in_0_fifo_eos_in, coord_in_1_fifo_eos_in,
            pos_in_0_fifo_eos_in, pos_in_1_fifo_eos_in} & {coord_in_0_fifo_valid_in,
            coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in, pos_in_1_fifo_valid_in})) &
            (&{coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in,
            pos_in_1_fifo_valid_in});
        inc_pos_cnt[1] = (~(|fifo_full)) & (&({coord_in_0_fifo_eos_in, coord_in_1_fifo_eos_in,
            pos_in_0_fifo_eos_in, pos_in_1_fifo_eos_in} & {coord_in_0_fifo_valid_in,
            coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in, pos_in_1_fifo_valid_in})) &
            (&{coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in,
            pos_in_1_fifo_valid_in});
        rst_pos_cnt[0] = 1'h0;
        rst_pos_cnt[1] = 1'h0;
        fifo_push = (~(|fifo_full)) & (&({coord_in_0_fifo_eos_in, coord_in_1_fifo_eos_in,
            pos_in_0_fifo_eos_in, pos_in_1_fifo_eos_in} & {coord_in_0_fifo_valid_in,
            coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in, pos_in_1_fifo_valid_in})) &
            (&{coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in,
            pos_in_1_fifo_valid_in});
        clr_eos_sticky[0] = 1'h0;
        clr_eos_sticky[1] = 1'h0;
        coord_to_fifo = coord_in_0_fifo_in[15:0];
        pos_to_fifo[0] = coord_in_0_fifo_in[15:0];
        pos_to_fifo[1] = coord_in_0_fifo_in[15:0];
        coord_to_fifo_eos = any_eos;
        pos_to_fifo_eos[0] = any_eos;
        pos_to_fifo_eos[1] = any_eos;
      end :intersect_seq_DRAIN_Output
    IDLE: begin :intersect_seq_IDLE_Output
        inc_pos_cnt[0] = 1'h0;
        inc_pos_cnt[1] = 1'h0;
        rst_pos_cnt[0] = 1'h0;
        rst_pos_cnt[1] = 1'h0;
        fifo_push = 1'h0;
        clr_eos_sticky[0] = 1'h0;
        clr_eos_sticky[1] = 1'h0;
        coord_to_fifo = 16'h0;
        pos_to_fifo[0] = 16'h0;
        pos_to_fifo[1] = 16'h0;
        coord_to_fifo_eos = 1'h0;
        pos_to_fifo_eos[0] = 1'h0;
        pos_to_fifo_eos[1] = 1'h0;
      end :intersect_seq_IDLE_Output
    ITER: begin :intersect_seq_ITER_Output
        inc_pos_cnt[0] = all_valid & (coord_in_0_fifo_in <= coord_in_1_fifo_in) & (~(|fifo_full));
        inc_pos_cnt[1] = all_valid & (coord_in_0_fifo_in >= coord_in_1_fifo_in) & (~(|fifo_full));
        rst_pos_cnt[0] = any_eos & (~(|fifo_full));
        rst_pos_cnt[1] = any_eos & (~(|fifo_full));
        fifo_push = all_valid & (coord_in_0_fifo_in == coord_in_1_fifo_in) & (~(|fifo_full)) &
            (~any_eos);
        clr_eos_sticky[0] = 1'h0;
        clr_eos_sticky[1] = 1'h0;
        coord_to_fifo = coord_in_0_fifo_in[15:0];
        pos_to_fifo[0] = pos_in_0_fifo_in[15:0];
        pos_to_fifo[1] = pos_in_1_fifo_in[15:0];
        coord_to_fifo_eos = 1'h0;
        pos_to_fifo_eos[0] = 1'h0;
        pos_to_fifo_eos[1] = 1'h0;
      end :intersect_seq_ITER_Output
    UNION: begin :intersect_seq_UNION_Output
        inc_pos_cnt[0] = all_valid_join & ((coord_in_0_fifo_in <= coord_in_1_fifo_in) |
            coord_in_1_fifo_eos_in) & (~(|fifo_full)) & (~coord_in_0_fifo_eos_in);
        inc_pos_cnt[1] = all_valid_join & ((coord_in_0_fifo_in >= coord_in_1_fifo_in) |
            coord_in_0_fifo_eos_in) & (~(|fifo_full)) & (~coord_in_1_fifo_eos_in);
        rst_pos_cnt[0] = any_eos & (~(|fifo_full));
        rst_pos_cnt[1] = any_eos & (~(|fifo_full));
        fifo_push = all_valid_join & (~(|fifo_full)) & (~(&({coord_in_0_fifo_eos_in,
            coord_in_1_fifo_eos_in, pos_in_0_fifo_eos_in, pos_in_1_fifo_eos_in} &
            {coord_in_0_fifo_valid_in, coord_in_1_fifo_valid_in, pos_in_0_fifo_valid_in,
            pos_in_1_fifo_valid_in})));
        clr_eos_sticky[0] = 1'h0;
        clr_eos_sticky[1] = 1'h0;
        coord_to_fifo = coord_in_0_fifo_eos_in ? coord_in_1_fifo_in[15:0]: coord_in_1_fifo_eos_in ?
            coord_in_0_fifo_in[15:0]: (coord_in_0_fifo_in <= coord_in_1_fifo_in) ?
            coord_in_0_fifo_in[15:0]: coord_in_1_fifo_in[15:0];
        pos_to_fifo[0] = coord_in_0_fifo_eos_in ? maybe: coord_in_1_fifo_eos_in ? pos_in_0_fifo_in[15:0]:
            (coord_in_0_fifo_in <= coord_in_1_fifo_in) ? pos_in_0_fifo_in[15:0]: maybe;
        pos_to_fifo[1] = coord_in_1_fifo_eos_in ? maybe: coord_in_0_fifo_eos_in ? pos_in_1_fifo_in[15:0]:
            (coord_in_1_fifo_in <= coord_in_0_fifo_in) ? pos_in_1_fifo_in[15:0]: maybe;
        coord_to_fifo_eos = 1'h0;
        pos_to_fifo_eos[0] = (pos_in_0_fifo_eos_in & (~coord_in_0_fifo_eos_in)) | (coord_in_0_fifo_eos_in ?
            1'h1: coord_in_1_fifo_eos_in ? 1'h0: (coord_in_0_fifo_in <= coord_in_1_fifo_in)
            ? 1'h0: 1'h1);
        pos_to_fifo_eos[1] = (pos_in_1_fifo_eos_in & (~coord_in_1_fifo_eos_in)) | (coord_in_1_fifo_eos_in ?
            1'h1: coord_in_0_fifo_eos_in ? 1'h0: (coord_in_1_fifo_in <= coord_in_0_fifo_in)
            ? 1'h0: 1'h1);
      end :intersect_seq_UNION_Output
    default: begin :intersect_seq_default_Output
        inc_pos_cnt[0] = 1'h0;
        inc_pos_cnt[1] = 1'h0;
        rst_pos_cnt[0] = 1'h0;
        rst_pos_cnt[1] = 1'h0;
        fifo_push = 1'h0;
        clr_eos_sticky[0] = 1'h0;
        clr_eos_sticky[1] = 1'h0;
        coord_to_fifo = 16'h0;
        pos_to_fifo[0] = 16'h0;
        pos_to_fifo[1] = 16'h0;
        coord_to_fifo_eos = 1'h0;
        pos_to_fifo_eos[0] = 1'h0;
        pos_to_fifo_eos[1] = 1'h0;
      end :intersect_seq_default_Output
  endcase
end
reg_fifo_depth_0_w_17_afd_2 coord_in_fifo_0 (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(coord_in_0),
  .flush(flush),
  .pop(inc_pos_cnt[0]),
  .push(coord_in_0_valid),
  .rst_n(rst_n),
  .data_out(coord_in_0_fifo_in),
  .empty(coord_in_fifo_0_empty),
  .full(coord_in_fifo_0_full)
);

reg_fifo_depth_0_w_17_afd_2 pos_in_fifo_0 (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(pos_in_0),
  .flush(flush),
  .pop(inc_pos_cnt[0]),
  .push(pos_in_0_valid),
  .rst_n(rst_n),
  .data_out(pos_in_0_fifo_in),
  .empty(pos_in_fifo_0_empty),
  .full(pos_in_fifo_0_full)
);

reg_fifo_depth_0_w_17_afd_2 coord_in_fifo_1 (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(coord_in_1),
  .flush(flush),
  .pop(inc_pos_cnt[1]),
  .push(coord_in_1_valid),
  .rst_n(rst_n),
  .data_out(coord_in_1_fifo_in),
  .empty(coord_in_fifo_1_empty),
  .full(coord_in_fifo_1_full)
);

reg_fifo_depth_0_w_17_afd_2 pos_in_fifo_1 (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(pos_in_1),
  .flush(flush),
  .pop(inc_pos_cnt[1]),
  .push(pos_in_1_valid),
  .rst_n(rst_n),
  .data_out(pos_in_1_fifo_in),
  .empty(pos_in_fifo_1_empty),
  .full(pos_in_fifo_1_full)
);

reg_fifo_depth_0_w_17_afd_2 coordinate_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(coord_fifo_in_packed),
  .flush(flush),
  .pop(coord_out_ready),
  .push(fifo_push),
  .rst_n(rst_n),
  .data_out(coord_fifo_out_packed),
  .empty(coordinate_fifo_empty),
  .full(coordinate_fifo_full)
);

reg_fifo_depth_0_w_17_afd_2 pos0_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(pos0_fifo_in_packed),
  .flush(flush),
  .pop(pos_out_0_ready),
  .push(fifo_push),
  .rst_n(rst_n),
  .data_out(pos0_fifo_out_packed),
  .empty(pos0_fifo_empty),
  .full(pos0_fifo_full)
);

reg_fifo_depth_0_w_17_afd_2 pos1_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(pos1_fifo_in_packed),
  .flush(flush),
  .pop(pos_out_1_ready),
  .push(fifo_push),
  .rst_n(rst_n),
  .data_out(pos1_fifo_out_packed),
  .empty(pos1_fifo_empty),
  .full(pos1_fifo_full)
);

endmodule   // intersect_unit

module intersect_unit_flat (
  input logic clk,
  input logic clk_en,
  input logic [0:0] [16:0] coord_in_0_f_,
  input logic coord_in_0_valid_f_,
  input logic [0:0] [16:0] coord_in_1_f_,
  input logic coord_in_1_valid_f_,
  input logic coord_out_ready_f_,
  input logic flush,
  input logic intersect_unit_inst_joiner_op,
  input logic intersect_unit_inst_tile_en,
  input logic [0:0] [16:0] pos_in_0_f_,
  input logic pos_in_0_valid_f_,
  input logic [0:0] [16:0] pos_in_1_f_,
  input logic pos_in_1_valid_f_,
  input logic pos_out_0_ready_f_,
  input logic pos_out_1_ready_f_,
  input logic rst_n,
  output logic coord_in_0_ready_f_,
  output logic coord_in_1_ready_f_,
  output logic [0:0] [16:0] coord_out_f_,
  output logic coord_out_valid_f_,
  output logic pos_in_0_ready_f_,
  output logic pos_in_1_ready_f_,
  output logic [0:0] [16:0] pos_out_0_f_,
  output logic pos_out_0_valid_f_,
  output logic [0:0] [16:0] pos_out_1_f_,
  output logic pos_out_1_valid_f_
);

intersect_unit intersect_unit_inst (
  .clk(clk),
  .clk_en(clk_en),
  .coord_in_0(coord_in_0_f_),
  .coord_in_0_valid(coord_in_0_valid_f_),
  .coord_in_1(coord_in_1_f_),
  .coord_in_1_valid(coord_in_1_valid_f_),
  .coord_out_ready(coord_out_ready_f_),
  .flush(flush),
  .joiner_op(intersect_unit_inst_joiner_op),
  .pos_in_0(pos_in_0_f_),
  .pos_in_0_valid(pos_in_0_valid_f_),
  .pos_in_1(pos_in_1_f_),
  .pos_in_1_valid(pos_in_1_valid_f_),
  .pos_out_0_ready(pos_out_0_ready_f_),
  .pos_out_1_ready(pos_out_1_ready_f_),
  .rst_n(rst_n),
  .tile_en(intersect_unit_inst_tile_en),
  .coord_in_0_ready(coord_in_0_ready_f_),
  .coord_in_1_ready(coord_in_1_ready_f_),
  .coord_out(coord_out_f_),
  .coord_out_valid(coord_out_valid_f_),
  .pos_in_0_ready(pos_in_0_ready_f_),
  .pos_in_1_ready(pos_in_1_ready_f_),
  .pos_out_0(pos_out_0_f_),
  .pos_out_0_valid(pos_out_0_valid_f_),
  .pos_out_1(pos_out_1_f_),
  .pos_out_1_valid(pos_out_1_valid_f_)
);

endmodule   // intersect_unit_flat

module reg_cr (
  input logic clk,
  input logic clk_en,
  input logic [16:0] data_in,
  input logic data_in_valid,
  input logic data_out_ready,
  input logic [15:0] default_value,
  input logic flush,
  input logic rst_n,
  input logic [15:0] stop_lvl,
  input logic tile_en,
  output logic data_in_ready,
  output logic [16:0] data_out,
  output logic data_out_valid
);

typedef enum logic[2:0] {
  ACCUM = 3'h0,
  DONE = 3'h1,
  OUTPUT = 3'h2,
  START = 3'h3,
  STOP_PASS = 3'h4
} accum_seq_state;
logic [15:0] accum_reg;
accum_seq_state accum_seq_current_state;
accum_seq_state accum_seq_next_state;
logic clr_once_popped;
logic [15:0] data_to_fifo;
logic gclk;
logic [16:0] infifo_in_packed;
logic [15:0] infifo_out_data;
logic infifo_out_eos;
logic [16:0] infifo_out_packed;
logic infifo_out_valid;
logic infifo_pop;
logic infifo_push;
logic input_fifo_empty;
logic input_fifo_full;
logic outfifo_full;
logic outfifo_in_eos;
logic [16:0] outfifo_in_packed;
logic [16:0] outfifo_out_packed;
logic outfifo_pop;
logic outfifo_push;
logic output_fifo_empty;
logic reg_accum;
logic reg_clr;
logic set_once_popped;
logic set_once_popped_sticky;
logic set_once_popped_was_high;
assign gclk = clk & tile_en;
assign data_in_ready = ~input_fifo_full;
assign infifo_in_packed[16:0] = data_in;
assign infifo_out_eos = infifo_out_packed[16];
assign infifo_out_data = infifo_out_packed[15:0];
assign infifo_push = data_in_valid;
assign infifo_out_valid = ~input_fifo_empty;
assign outfifo_in_packed[16] = outfifo_in_eos;
assign outfifo_in_packed[15:0] = data_to_fifo;
assign data_out = outfifo_out_packed[16:0];

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    set_once_popped_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      set_once_popped_was_high <= 1'h0;
    end
    else if (clr_once_popped) begin
      set_once_popped_was_high <= 1'h0;
    end
    else if (set_once_popped) begin
      set_once_popped_was_high <= 1'h1;
    end
  end
end
assign set_once_popped_sticky = set_once_popped_was_high;
assign data_out_valid = ~output_fifo_empty;
assign outfifo_pop = data_out_ready;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    accum_reg <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      accum_reg <= 16'h0;
    end
    else if (reg_clr) begin
      accum_reg <= default_value;
    end
    else if (reg_accum) begin
      accum_reg <= accum_reg + infifo_out_data;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (!rst_n) begin
    accum_seq_current_state <= START;
  end
  else if (clk_en) begin
    if (flush) begin
      accum_seq_current_state <= START;
    end
    else accum_seq_current_state <= accum_seq_next_state;
  end
end
always_comb begin
  accum_seq_next_state = accum_seq_current_state;
  unique case (accum_seq_current_state)
    ACCUM: begin
        if (infifo_out_valid & infifo_out_eos) begin
          accum_seq_next_state = OUTPUT;
        end
        else accum_seq_next_state = ACCUM;
      end
    DONE: begin
        if (~outfifo_full) begin
          accum_seq_next_state = START;
        end
        else accum_seq_next_state = DONE;
      end
    OUTPUT: begin
        if (~outfifo_full) begin
          accum_seq_next_state = STOP_PASS;
        end
        else accum_seq_next_state = OUTPUT;
      end
    START: begin
        if (infifo_out_valid & (~infifo_out_eos)) begin
          accum_seq_next_state = ACCUM;
        end
        else if (infifo_out_valid & infifo_out_eos & (infifo_out_data[9:8] == 2'h1)) begin
          accum_seq_next_state = DONE;
        end
        else if (infifo_out_valid & infifo_out_eos & (infifo_out_data[9:8] == 2'h0)) begin
          accum_seq_next_state = OUTPUT;
        end
        else accum_seq_next_state = START;
      end
    STOP_PASS: begin
        if (~outfifo_full) begin
          accum_seq_next_state = START;
        end
        else accum_seq_next_state = STOP_PASS;
      end
    default: accum_seq_next_state = accum_seq_current_state;
  endcase
end
always_comb begin
  unique case (accum_seq_current_state)
    ACCUM: begin :accum_seq_ACCUM_Output
        infifo_pop = infifo_out_valid & (~infifo_out_eos);
        outfifo_push = 1'h0;
        reg_clr = 1'h0;
        reg_accum = infifo_out_valid & (~infifo_out_eos);
        data_to_fifo = 16'h0;
        outfifo_in_eos = 1'h0;
        set_once_popped = 1'h0;
        clr_once_popped = 1'h0;
      end :accum_seq_ACCUM_Output
    DONE: begin :accum_seq_DONE_Output
        infifo_pop = ~outfifo_full;
        outfifo_push = ~outfifo_full;
        reg_clr = 1'h1;
        reg_accum = 1'h0;
        data_to_fifo = infifo_out_data;
        outfifo_in_eos = infifo_out_eos;
        set_once_popped = 1'h0;
        clr_once_popped = 1'h1;
      end :accum_seq_DONE_Output
    OUTPUT: begin :accum_seq_OUTPUT_Output
        infifo_pop = 1'h0;
        outfifo_push = ~outfifo_full;
        reg_clr = 1'h0;
        reg_accum = 1'h0;
        data_to_fifo = accum_reg;
        outfifo_in_eos = 1'h0;
        set_once_popped = 1'h0;
        clr_once_popped = 1'h0;
      end :accum_seq_OUTPUT_Output
    START: begin :accum_seq_START_Output
        infifo_pop = 1'h0;
        outfifo_push = 1'h0;
        reg_clr = 1'h0;
        reg_accum = 1'h0;
        data_to_fifo = 16'h0;
        outfifo_in_eos = 1'h0;
        set_once_popped = 1'h0;
        clr_once_popped = 1'h0;
      end :accum_seq_START_Output
    STOP_PASS: begin :accum_seq_STOP_PASS_Output
        infifo_pop = (~outfifo_full) & infifo_out_valid & infifo_out_eos & (infifo_out_data[9:8] ==
            2'h0);
        outfifo_push = (~outfifo_full) & infifo_out_valid & infifo_out_eos & (infifo_out_data[9:8] ==
            2'h0) & (infifo_out_data[7:0] > 8'h0);
        reg_clr = 1'h1;
        reg_accum = 1'h0;
        data_to_fifo = infifo_out_data - 16'h1;
        outfifo_in_eos = 1'h1;
        set_once_popped = 1'h0;
        clr_once_popped = 1'h1;
      end :accum_seq_STOP_PASS_Output
    default: begin :accum_seq_default_Output
        infifo_pop = 1'h0;
        outfifo_push = 1'h0;
        reg_clr = 1'h0;
        reg_accum = 1'h0;
        data_to_fifo = 16'h0;
        outfifo_in_eos = 1'h0;
        set_once_popped = 1'h0;
        clr_once_popped = 1'h0;
      end :accum_seq_default_Output
  endcase
end
reg_fifo_depth_0_w_17_afd_2 input_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(infifo_in_packed),
  .flush(flush),
  .pop(infifo_pop),
  .push(infifo_push),
  .rst_n(rst_n),
  .data_out(infifo_out_packed),
  .empty(input_fifo_empty),
  .full(input_fifo_full)
);

reg_fifo_depth_0_w_17_afd_2 output_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(outfifo_in_packed),
  .flush(flush),
  .pop(outfifo_pop),
  .push(outfifo_push),
  .rst_n(rst_n),
  .data_out(outfifo_out_packed),
  .empty(output_fifo_empty),
  .full(outfifo_full)
);

endmodule   // reg_cr

module reg_cr_flat (
  input logic clk,
  input logic clk_en,
  input logic [0:0] [16:0] data_in_f_,
  input logic data_in_valid_f_,
  input logic data_out_ready_f_,
  input logic flush,
  input logic [15:0] reg_cr_inst_default_value,
  input logic [15:0] reg_cr_inst_stop_lvl,
  input logic reg_cr_inst_tile_en,
  input logic rst_n,
  output logic data_in_ready_f_,
  output logic [0:0] [16:0] data_out_f_,
  output logic data_out_valid_f_
);

reg_cr reg_cr_inst (
  .clk(clk),
  .clk_en(clk_en),
  .data_in(data_in_f_),
  .data_in_valid(data_in_valid_f_),
  .data_out_ready(data_out_ready_f_),
  .default_value(reg_cr_inst_default_value),
  .flush(flush),
  .rst_n(rst_n),
  .stop_lvl(reg_cr_inst_stop_lvl),
  .tile_en(reg_cr_inst_tile_en),
  .data_in_ready(data_in_ready_f_),
  .data_out(data_out_f_),
  .data_out_valid(data_out_valid_f_)
);

endmodule   // reg_cr_flat

module reg_fifo_depth_0_w_17_afd_2 (
  input logic clk,
  input logic clk_en,
  input logic [0:0] [16:0] data_in,
  input logic flush,
  input logic pop,
  input logic push,
  input logic rst_n,
  output logic almost_full,
  output logic [0:0] [16:0] data_out,
  output logic empty,
  output logic full,
  output logic valid
);

assign data_out = data_in;
assign valid = push;
assign empty = ~push;
assign full = ~pop;
assign almost_full = ~pop;
endmodule   // reg_fifo_depth_0_w_17_afd_2

module reg_fifo_depth_2_w_17_afd_2 (
  input logic clk,
  input logic clk_en,
  input logic [0:0] [16:0] data_in,
  input logic flush,
  input logic pop,
  input logic push,
  input logic rst_n,
  output logic almost_full,
  output logic [0:0] [16:0] data_out,
  output logic empty,
  output logic full,
  output logic valid
);

logic [1:0] num_items;
logic passthru;
logic rd_ptr;
logic read;
logic [1:0][0:0][16:0] reg_array;
logic wr_ptr;
logic write;
assign full = num_items == 2'h2;
assign almost_full = num_items >= 2'h0;
assign empty = num_items == 2'h0;
assign read = pop & (~passthru) & (~empty);
assign passthru = 1'h0;
assign write = push & (~passthru) & (~full);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_items <= 2'h0;
  end
  else if (flush) begin
    num_items <= 2'h0;
  end
  else if (clk_en) begin
    if (write & (~read)) begin
      num_items <= num_items + 2'h1;
    end
    else if ((~write) & read) begin
      num_items <= num_items - 2'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    reg_array <= 34'h0;
  end
  else if (flush) begin
    reg_array <= 34'h0;
  end
  else if (clk_en) begin
    if (write) begin
      reg_array[wr_ptr] <= data_in;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    wr_ptr <= 1'h0;
  end
  else if (flush) begin
    wr_ptr <= 1'h0;
  end
  else if (clk_en) begin
    if (write) begin
      if (wr_ptr == 1'h1) begin
        wr_ptr <= 1'h0;
      end
      else wr_ptr <= wr_ptr + 1'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    rd_ptr <= 1'h0;
  end
  else if (flush) begin
    rd_ptr <= 1'h0;
  end
  else if (clk_en) begin
    if (read) begin
      rd_ptr <= rd_ptr + 1'h1;
    end
  end
end
always_comb begin
  if (passthru) begin
    data_out = data_in;
  end
  else data_out = reg_array[rd_ptr];
end
always_comb begin
  valid = (~empty) | passthru;
end
endmodule   // reg_fifo_depth_2_w_17_afd_2


module Or4x32 (
    input [31:0] I0,
    input [31:0] I1,
    input [31:0] I2,
    input [31:0] I3,
    output [31:0] O
);
wire orr_inst0_out;
wire orr_inst1_out;
wire orr_inst10_out;
wire orr_inst11_out;
wire orr_inst12_out;
wire orr_inst13_out;
wire orr_inst14_out;
wire orr_inst15_out;
wire orr_inst16_out;
wire orr_inst17_out;
wire orr_inst18_out;
wire orr_inst19_out;
wire orr_inst2_out;
wire orr_inst20_out;
wire orr_inst21_out;
wire orr_inst22_out;
wire orr_inst23_out;
wire orr_inst24_out;
wire orr_inst25_out;
wire orr_inst26_out;
wire orr_inst27_out;
wire orr_inst28_out;
wire orr_inst29_out;
wire orr_inst3_out;
wire orr_inst30_out;
wire orr_inst31_out;
wire orr_inst4_out;
wire orr_inst5_out;
wire orr_inst6_out;
wire orr_inst7_out;
wire orr_inst8_out;
wire orr_inst9_out;
wire [3:0] orr_inst0_in;
assign orr_inst0_in = {I3[0],I2[0],I1[0],I0[0]};
coreir_orr #(
    .width(4)
) orr_inst0 (
    .in(orr_inst0_in),
    .out(orr_inst0_out)
);
wire [3:0] orr_inst1_in;
assign orr_inst1_in = {I3[1],I2[1],I1[1],I0[1]};
coreir_orr #(
    .width(4)
) orr_inst1 (
    .in(orr_inst1_in),
    .out(orr_inst1_out)
);
wire [3:0] orr_inst10_in;
assign orr_inst10_in = {I3[10],I2[10],I1[10],I0[10]};
coreir_orr #(
    .width(4)
) orr_inst10 (
    .in(orr_inst10_in),
    .out(orr_inst10_out)
);
wire [3:0] orr_inst11_in;
assign orr_inst11_in = {I3[11],I2[11],I1[11],I0[11]};
coreir_orr #(
    .width(4)
) orr_inst11 (
    .in(orr_inst11_in),
    .out(orr_inst11_out)
);
wire [3:0] orr_inst12_in;
assign orr_inst12_in = {I3[12],I2[12],I1[12],I0[12]};
coreir_orr #(
    .width(4)
) orr_inst12 (
    .in(orr_inst12_in),
    .out(orr_inst12_out)
);
wire [3:0] orr_inst13_in;
assign orr_inst13_in = {I3[13],I2[13],I1[13],I0[13]};
coreir_orr #(
    .width(4)
) orr_inst13 (
    .in(orr_inst13_in),
    .out(orr_inst13_out)
);
wire [3:0] orr_inst14_in;
assign orr_inst14_in = {I3[14],I2[14],I1[14],I0[14]};
coreir_orr #(
    .width(4)
) orr_inst14 (
    .in(orr_inst14_in),
    .out(orr_inst14_out)
);
wire [3:0] orr_inst15_in;
assign orr_inst15_in = {I3[15],I2[15],I1[15],I0[15]};
coreir_orr #(
    .width(4)
) orr_inst15 (
    .in(orr_inst15_in),
    .out(orr_inst15_out)
);
wire [3:0] orr_inst16_in;
assign orr_inst16_in = {I3[16],I2[16],I1[16],I0[16]};
coreir_orr #(
    .width(4)
) orr_inst16 (
    .in(orr_inst16_in),
    .out(orr_inst16_out)
);
wire [3:0] orr_inst17_in;
assign orr_inst17_in = {I3[17],I2[17],I1[17],I0[17]};
coreir_orr #(
    .width(4)
) orr_inst17 (
    .in(orr_inst17_in),
    .out(orr_inst17_out)
);
wire [3:0] orr_inst18_in;
assign orr_inst18_in = {I3[18],I2[18],I1[18],I0[18]};
coreir_orr #(
    .width(4)
) orr_inst18 (
    .in(orr_inst18_in),
    .out(orr_inst18_out)
);
wire [3:0] orr_inst19_in;
assign orr_inst19_in = {I3[19],I2[19],I1[19],I0[19]};
coreir_orr #(
    .width(4)
) orr_inst19 (
    .in(orr_inst19_in),
    .out(orr_inst19_out)
);
wire [3:0] orr_inst2_in;
assign orr_inst2_in = {I3[2],I2[2],I1[2],I0[2]};
coreir_orr #(
    .width(4)
) orr_inst2 (
    .in(orr_inst2_in),
    .out(orr_inst2_out)
);
wire [3:0] orr_inst20_in;
assign orr_inst20_in = {I3[20],I2[20],I1[20],I0[20]};
coreir_orr #(
    .width(4)
) orr_inst20 (
    .in(orr_inst20_in),
    .out(orr_inst20_out)
);
wire [3:0] orr_inst21_in;
assign orr_inst21_in = {I3[21],I2[21],I1[21],I0[21]};
coreir_orr #(
    .width(4)
) orr_inst21 (
    .in(orr_inst21_in),
    .out(orr_inst21_out)
);
wire [3:0] orr_inst22_in;
assign orr_inst22_in = {I3[22],I2[22],I1[22],I0[22]};
coreir_orr #(
    .width(4)
) orr_inst22 (
    .in(orr_inst22_in),
    .out(orr_inst22_out)
);
wire [3:0] orr_inst23_in;
assign orr_inst23_in = {I3[23],I2[23],I1[23],I0[23]};
coreir_orr #(
    .width(4)
) orr_inst23 (
    .in(orr_inst23_in),
    .out(orr_inst23_out)
);
wire [3:0] orr_inst24_in;
assign orr_inst24_in = {I3[24],I2[24],I1[24],I0[24]};
coreir_orr #(
    .width(4)
) orr_inst24 (
    .in(orr_inst24_in),
    .out(orr_inst24_out)
);
wire [3:0] orr_inst25_in;
assign orr_inst25_in = {I3[25],I2[25],I1[25],I0[25]};
coreir_orr #(
    .width(4)
) orr_inst25 (
    .in(orr_inst25_in),
    .out(orr_inst25_out)
);
wire [3:0] orr_inst26_in;
assign orr_inst26_in = {I3[26],I2[26],I1[26],I0[26]};
coreir_orr #(
    .width(4)
) orr_inst26 (
    .in(orr_inst26_in),
    .out(orr_inst26_out)
);
wire [3:0] orr_inst27_in;
assign orr_inst27_in = {I3[27],I2[27],I1[27],I0[27]};
coreir_orr #(
    .width(4)
) orr_inst27 (
    .in(orr_inst27_in),
    .out(orr_inst27_out)
);
wire [3:0] orr_inst28_in;
assign orr_inst28_in = {I3[28],I2[28],I1[28],I0[28]};
coreir_orr #(
    .width(4)
) orr_inst28 (
    .in(orr_inst28_in),
    .out(orr_inst28_out)
);
wire [3:0] orr_inst29_in;
assign orr_inst29_in = {I3[29],I2[29],I1[29],I0[29]};
coreir_orr #(
    .width(4)
) orr_inst29 (
    .in(orr_inst29_in),
    .out(orr_inst29_out)
);
wire [3:0] orr_inst3_in;
assign orr_inst3_in = {I3[3],I2[3],I1[3],I0[3]};
coreir_orr #(
    .width(4)
) orr_inst3 (
    .in(orr_inst3_in),
    .out(orr_inst3_out)
);
wire [3:0] orr_inst30_in;
assign orr_inst30_in = {I3[30],I2[30],I1[30],I0[30]};
coreir_orr #(
    .width(4)
) orr_inst30 (
    .in(orr_inst30_in),
    .out(orr_inst30_out)
);
wire [3:0] orr_inst31_in;
assign orr_inst31_in = {I3[31],I2[31],I1[31],I0[31]};
coreir_orr #(
    .width(4)
) orr_inst31 (
    .in(orr_inst31_in),
    .out(orr_inst31_out)
);
wire [3:0] orr_inst4_in;
assign orr_inst4_in = {I3[4],I2[4],I1[4],I0[4]};
coreir_orr #(
    .width(4)
) orr_inst4 (
    .in(orr_inst4_in),
    .out(orr_inst4_out)
);
wire [3:0] orr_inst5_in;
assign orr_inst5_in = {I3[5],I2[5],I1[5],I0[5]};
coreir_orr #(
    .width(4)
) orr_inst5 (
    .in(orr_inst5_in),
    .out(orr_inst5_out)
);
wire [3:0] orr_inst6_in;
assign orr_inst6_in = {I3[6],I2[6],I1[6],I0[6]};
coreir_orr #(
    .width(4)
) orr_inst6 (
    .in(orr_inst6_in),
    .out(orr_inst6_out)
);
wire [3:0] orr_inst7_in;
assign orr_inst7_in = {I3[7],I2[7],I1[7],I0[7]};
coreir_orr #(
    .width(4)
) orr_inst7 (
    .in(orr_inst7_in),
    .out(orr_inst7_out)
);
wire [3:0] orr_inst8_in;
assign orr_inst8_in = {I3[8],I2[8],I1[8],I0[8]};
coreir_orr #(
    .width(4)
) orr_inst8 (
    .in(orr_inst8_in),
    .out(orr_inst8_out)
);
wire [3:0] orr_inst9_in;
assign orr_inst9_in = {I3[9],I2[9],I1[9],I0[9]};
coreir_orr #(
    .width(4)
) orr_inst9 (
    .in(orr_inst9_in),
    .out(orr_inst9_out)
);
assign O = {orr_inst31_out,orr_inst30_out,orr_inst29_out,orr_inst28_out,orr_inst27_out,orr_inst26_out,orr_inst25_out,orr_inst24_out,orr_inst23_out,orr_inst22_out,orr_inst21_out,orr_inst20_out,orr_inst19_out,orr_inst18_out,orr_inst17_out,orr_inst16_out,orr_inst15_out,orr_inst14_out,orr_inst13_out,orr_inst12_out,orr_inst11_out,orr_inst10_out,orr_inst9_out,orr_inst8_out,orr_inst7_out,orr_inst6_out,orr_inst5_out,orr_inst4_out,orr_inst3_out,orr_inst2_out,orr_inst1_out,orr_inst0_out};
endmodule

module Or3x8 (
    input [7:0] I0,
    input [7:0] I1,
    input [7:0] I2,
    output [7:0] O
);
wire orr_inst0_out;
wire orr_inst1_out;
wire orr_inst2_out;
wire orr_inst3_out;
wire orr_inst4_out;
wire orr_inst5_out;
wire orr_inst6_out;
wire orr_inst7_out;
wire [2:0] orr_inst0_in;
assign orr_inst0_in = {I2[0],I1[0],I0[0]};
coreir_orr #(
    .width(3)
) orr_inst0 (
    .in(orr_inst0_in),
    .out(orr_inst0_out)
);
wire [2:0] orr_inst1_in;
assign orr_inst1_in = {I2[1],I1[1],I0[1]};
coreir_orr #(
    .width(3)
) orr_inst1 (
    .in(orr_inst1_in),
    .out(orr_inst1_out)
);
wire [2:0] orr_inst2_in;
assign orr_inst2_in = {I2[2],I1[2],I0[2]};
coreir_orr #(
    .width(3)
) orr_inst2 (
    .in(orr_inst2_in),
    .out(orr_inst2_out)
);
wire [2:0] orr_inst3_in;
assign orr_inst3_in = {I2[3],I1[3],I0[3]};
coreir_orr #(
    .width(3)
) orr_inst3 (
    .in(orr_inst3_in),
    .out(orr_inst3_out)
);
wire [2:0] orr_inst4_in;
assign orr_inst4_in = {I2[4],I1[4],I0[4]};
coreir_orr #(
    .width(3)
) orr_inst4 (
    .in(orr_inst4_in),
    .out(orr_inst4_out)
);
wire [2:0] orr_inst5_in;
assign orr_inst5_in = {I2[5],I1[5],I0[5]};
coreir_orr #(
    .width(3)
) orr_inst5 (
    .in(orr_inst5_in),
    .out(orr_inst5_out)
);
wire [2:0] orr_inst6_in;
assign orr_inst6_in = {I2[6],I1[6],I0[6]};
coreir_orr #(
    .width(3)
) orr_inst6 (
    .in(orr_inst6_in),
    .out(orr_inst6_out)
);
wire [2:0] orr_inst7_in;
assign orr_inst7_in = {I2[7],I1[7],I0[7]};
coreir_orr #(
    .width(3)
) orr_inst7 (
    .in(orr_inst7_in),
    .out(orr_inst7_out)
);
assign O = {orr_inst7_out,orr_inst6_out,orr_inst5_out,orr_inst4_out,orr_inst3_out,orr_inst2_out,orr_inst1_out,orr_inst0_out};
endmodule

module Or3x32 (
    input [31:0] I0,
    input [31:0] I1,
    input [31:0] I2,
    output [31:0] O
);
wire orr_inst0_out;
wire orr_inst1_out;
wire orr_inst10_out;
wire orr_inst11_out;
wire orr_inst12_out;
wire orr_inst13_out;
wire orr_inst14_out;
wire orr_inst15_out;
wire orr_inst16_out;
wire orr_inst17_out;
wire orr_inst18_out;
wire orr_inst19_out;
wire orr_inst2_out;
wire orr_inst20_out;
wire orr_inst21_out;
wire orr_inst22_out;
wire orr_inst23_out;
wire orr_inst24_out;
wire orr_inst25_out;
wire orr_inst26_out;
wire orr_inst27_out;
wire orr_inst28_out;
wire orr_inst29_out;
wire orr_inst3_out;
wire orr_inst30_out;
wire orr_inst31_out;
wire orr_inst4_out;
wire orr_inst5_out;
wire orr_inst6_out;
wire orr_inst7_out;
wire orr_inst8_out;
wire orr_inst9_out;
wire [2:0] orr_inst0_in;
assign orr_inst0_in = {I2[0],I1[0],I0[0]};
coreir_orr #(
    .width(3)
) orr_inst0 (
    .in(orr_inst0_in),
    .out(orr_inst0_out)
);
wire [2:0] orr_inst1_in;
assign orr_inst1_in = {I2[1],I1[1],I0[1]};
coreir_orr #(
    .width(3)
) orr_inst1 (
    .in(orr_inst1_in),
    .out(orr_inst1_out)
);
wire [2:0] orr_inst10_in;
assign orr_inst10_in = {I2[10],I1[10],I0[10]};
coreir_orr #(
    .width(3)
) orr_inst10 (
    .in(orr_inst10_in),
    .out(orr_inst10_out)
);
wire [2:0] orr_inst11_in;
assign orr_inst11_in = {I2[11],I1[11],I0[11]};
coreir_orr #(
    .width(3)
) orr_inst11 (
    .in(orr_inst11_in),
    .out(orr_inst11_out)
);
wire [2:0] orr_inst12_in;
assign orr_inst12_in = {I2[12],I1[12],I0[12]};
coreir_orr #(
    .width(3)
) orr_inst12 (
    .in(orr_inst12_in),
    .out(orr_inst12_out)
);
wire [2:0] orr_inst13_in;
assign orr_inst13_in = {I2[13],I1[13],I0[13]};
coreir_orr #(
    .width(3)
) orr_inst13 (
    .in(orr_inst13_in),
    .out(orr_inst13_out)
);
wire [2:0] orr_inst14_in;
assign orr_inst14_in = {I2[14],I1[14],I0[14]};
coreir_orr #(
    .width(3)
) orr_inst14 (
    .in(orr_inst14_in),
    .out(orr_inst14_out)
);
wire [2:0] orr_inst15_in;
assign orr_inst15_in = {I2[15],I1[15],I0[15]};
coreir_orr #(
    .width(3)
) orr_inst15 (
    .in(orr_inst15_in),
    .out(orr_inst15_out)
);
wire [2:0] orr_inst16_in;
assign orr_inst16_in = {I2[16],I1[16],I0[16]};
coreir_orr #(
    .width(3)
) orr_inst16 (
    .in(orr_inst16_in),
    .out(orr_inst16_out)
);
wire [2:0] orr_inst17_in;
assign orr_inst17_in = {I2[17],I1[17],I0[17]};
coreir_orr #(
    .width(3)
) orr_inst17 (
    .in(orr_inst17_in),
    .out(orr_inst17_out)
);
wire [2:0] orr_inst18_in;
assign orr_inst18_in = {I2[18],I1[18],I0[18]};
coreir_orr #(
    .width(3)
) orr_inst18 (
    .in(orr_inst18_in),
    .out(orr_inst18_out)
);
wire [2:0] orr_inst19_in;
assign orr_inst19_in = {I2[19],I1[19],I0[19]};
coreir_orr #(
    .width(3)
) orr_inst19 (
    .in(orr_inst19_in),
    .out(orr_inst19_out)
);
wire [2:0] orr_inst2_in;
assign orr_inst2_in = {I2[2],I1[2],I0[2]};
coreir_orr #(
    .width(3)
) orr_inst2 (
    .in(orr_inst2_in),
    .out(orr_inst2_out)
);
wire [2:0] orr_inst20_in;
assign orr_inst20_in = {I2[20],I1[20],I0[20]};
coreir_orr #(
    .width(3)
) orr_inst20 (
    .in(orr_inst20_in),
    .out(orr_inst20_out)
);
wire [2:0] orr_inst21_in;
assign orr_inst21_in = {I2[21],I1[21],I0[21]};
coreir_orr #(
    .width(3)
) orr_inst21 (
    .in(orr_inst21_in),
    .out(orr_inst21_out)
);
wire [2:0] orr_inst22_in;
assign orr_inst22_in = {I2[22],I1[22],I0[22]};
coreir_orr #(
    .width(3)
) orr_inst22 (
    .in(orr_inst22_in),
    .out(orr_inst22_out)
);
wire [2:0] orr_inst23_in;
assign orr_inst23_in = {I2[23],I1[23],I0[23]};
coreir_orr #(
    .width(3)
) orr_inst23 (
    .in(orr_inst23_in),
    .out(orr_inst23_out)
);
wire [2:0] orr_inst24_in;
assign orr_inst24_in = {I2[24],I1[24],I0[24]};
coreir_orr #(
    .width(3)
) orr_inst24 (
    .in(orr_inst24_in),
    .out(orr_inst24_out)
);
wire [2:0] orr_inst25_in;
assign orr_inst25_in = {I2[25],I1[25],I0[25]};
coreir_orr #(
    .width(3)
) orr_inst25 (
    .in(orr_inst25_in),
    .out(orr_inst25_out)
);
wire [2:0] orr_inst26_in;
assign orr_inst26_in = {I2[26],I1[26],I0[26]};
coreir_orr #(
    .width(3)
) orr_inst26 (
    .in(orr_inst26_in),
    .out(orr_inst26_out)
);
wire [2:0] orr_inst27_in;
assign orr_inst27_in = {I2[27],I1[27],I0[27]};
coreir_orr #(
    .width(3)
) orr_inst27 (
    .in(orr_inst27_in),
    .out(orr_inst27_out)
);
wire [2:0] orr_inst28_in;
assign orr_inst28_in = {I2[28],I1[28],I0[28]};
coreir_orr #(
    .width(3)
) orr_inst28 (
    .in(orr_inst28_in),
    .out(orr_inst28_out)
);
wire [2:0] orr_inst29_in;
assign orr_inst29_in = {I2[29],I1[29],I0[29]};
coreir_orr #(
    .width(3)
) orr_inst29 (
    .in(orr_inst29_in),
    .out(orr_inst29_out)
);
wire [2:0] orr_inst3_in;
assign orr_inst3_in = {I2[3],I1[3],I0[3]};
coreir_orr #(
    .width(3)
) orr_inst3 (
    .in(orr_inst3_in),
    .out(orr_inst3_out)
);
wire [2:0] orr_inst30_in;
assign orr_inst30_in = {I2[30],I1[30],I0[30]};
coreir_orr #(
    .width(3)
) orr_inst30 (
    .in(orr_inst30_in),
    .out(orr_inst30_out)
);
wire [2:0] orr_inst31_in;
assign orr_inst31_in = {I2[31],I1[31],I0[31]};
coreir_orr #(
    .width(3)
) orr_inst31 (
    .in(orr_inst31_in),
    .out(orr_inst31_out)
);
wire [2:0] orr_inst4_in;
assign orr_inst4_in = {I2[4],I1[4],I0[4]};
coreir_orr #(
    .width(3)
) orr_inst4 (
    .in(orr_inst4_in),
    .out(orr_inst4_out)
);
wire [2:0] orr_inst5_in;
assign orr_inst5_in = {I2[5],I1[5],I0[5]};
coreir_orr #(
    .width(3)
) orr_inst5 (
    .in(orr_inst5_in),
    .out(orr_inst5_out)
);
wire [2:0] orr_inst6_in;
assign orr_inst6_in = {I2[6],I1[6],I0[6]};
coreir_orr #(
    .width(3)
) orr_inst6 (
    .in(orr_inst6_in),
    .out(orr_inst6_out)
);
wire [2:0] orr_inst7_in;
assign orr_inst7_in = {I2[7],I1[7],I0[7]};
coreir_orr #(
    .width(3)
) orr_inst7 (
    .in(orr_inst7_in),
    .out(orr_inst7_out)
);
wire [2:0] orr_inst8_in;
assign orr_inst8_in = {I2[8],I1[8],I0[8]};
coreir_orr #(
    .width(3)
) orr_inst8 (
    .in(orr_inst8_in),
    .out(orr_inst8_out)
);
wire [2:0] orr_inst9_in;
assign orr_inst9_in = {I2[9],I1[9],I0[9]};
coreir_orr #(
    .width(3)
) orr_inst9 (
    .in(orr_inst9_in),
    .out(orr_inst9_out)
);
assign O = {orr_inst31_out,orr_inst30_out,orr_inst29_out,orr_inst28_out,orr_inst27_out,orr_inst26_out,orr_inst25_out,orr_inst24_out,orr_inst23_out,orr_inst22_out,orr_inst21_out,orr_inst20_out,orr_inst19_out,orr_inst18_out,orr_inst17_out,orr_inst16_out,orr_inst15_out,orr_inst14_out,orr_inst13_out,orr_inst12_out,orr_inst11_out,orr_inst10_out,orr_inst9_out,orr_inst8_out,orr_inst7_out,orr_inst6_out,orr_inst5_out,orr_inst4_out,orr_inst3_out,orr_inst2_out,orr_inst1_out,orr_inst0_out};
endmodule

module MuxWrapperAOI_1_1_RegularReadyValid (
    input [0:0] I,
    output [0:0] O,
    input ready_in,
    output ready_out,
    input valid_in,
    output valid_out
);
assign O = I;
assign ready_out = ready_in;
assign valid_out = valid_in;
endmodule

module MuxWrapperAOI_1_1_ConstReadyValid (
    input [0:0] I,
    output [0:0] O,
    input ready_in,
    output ready_out,
    input valid_in,
    output valid_out
);
assign O = I;
assign ready_out = ready_in;
assign valid_out = valid_in;
endmodule

module MuxWrapperAOI_1_17_RegularReadyValid (
    input [16:0] I,
    output [16:0] O,
    input ready_in,
    output ready_out,
    input valid_in,
    output valid_out
);
assign O = I;
assign ready_out = ready_in;
assign valid_out = valid_in;
endmodule

module MuxWrapperAOI_1_17_ConstReadyValid (
    input [16:0] I,
    output [16:0] O,
    input ready_in,
    output ready_out,
    input valid_in,
    output valid_out
);
assign O = I;
assign ready_out = ready_in;
assign valid_out = valid_in;
endmodule

module MuxWithDefaultWrapper_6_32_8_0 (
    input [31:0] I [5:0],
    input [7:0] S,
    input [0:0] EN,
    output [31:0] O
);
wire [31:0] const_0_32_out;
wire [7:0] const_6_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_ult_inst0_out;
wire [31:0] mux_aoi_2_32_inst0_O;
wire [1:0] mux_aoi_2_32_inst0_out_sel;
wire [31:0] mux_aoi_6_32_inst0_O;
wire [7:0] mux_aoi_6_32_inst0_out_sel;
coreir_const #(
    .value(32'h00000000),
    .width(32)
) const_0_32 (
    .out(const_0_32_out)
);
coreir_const #(
    .value(8'h06),
    .width(8)
) const_6_8 (
    .out(const_6_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_ult_inst0_out),
    .in1(EN[0]),
    .out(magma_Bit_and_inst0_out)
);
coreir_ult #(
    .width(8)
) magma_Bits_8_ult_inst0 (
    .in0(S),
    .in1(const_6_8_out),
    .out(magma_Bits_8_ult_inst0_out)
);
wire [31:0] mux_aoi_2_32_inst0_I [1:0];
assign mux_aoi_2_32_inst0_I[1] = mux_aoi_6_32_inst0_O;
assign mux_aoi_2_32_inst0_I[0] = const_0_32_out;
mux_aoi_2_32 mux_aoi_2_32_inst0 (
    .I(mux_aoi_2_32_inst0_I),
    .O(mux_aoi_2_32_inst0_O),
    .S(magma_Bit_and_inst0_out),
    .out_sel(mux_aoi_2_32_inst0_out_sel)
);
wire [31:0] mux_aoi_6_32_inst0_I [5:0];
assign mux_aoi_6_32_inst0_I[5] = I[5];
assign mux_aoi_6_32_inst0_I[4] = I[4];
assign mux_aoi_6_32_inst0_I[3] = I[3];
assign mux_aoi_6_32_inst0_I[2] = I[2];
assign mux_aoi_6_32_inst0_I[1] = I[1];
assign mux_aoi_6_32_inst0_I[0] = I[0];
mux_aoi_6_32 mux_aoi_6_32_inst0 (
    .I(mux_aoi_6_32_inst0_I),
    .O(mux_aoi_6_32_inst0_O),
    .S(S[2:0]),
    .out_sel(mux_aoi_6_32_inst0_out_sel)
);
assign O = mux_aoi_2_32_inst0_O;
endmodule

module MuxWithDefaultWrapper_16_32_8_0 (
    input [31:0] I [15:0],
    input [7:0] S,
    input [0:0] EN,
    output [31:0] O
);
wire [31:0] const_0_32_out;
wire [7:0] const_16_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_ult_inst0_out;
wire [31:0] mux_aoi_16_32_inst0_O;
wire [15:0] mux_aoi_16_32_inst0_out_sel;
wire [31:0] mux_aoi_2_32_inst0_O;
wire [1:0] mux_aoi_2_32_inst0_out_sel;
coreir_const #(
    .value(32'h00000000),
    .width(32)
) const_0_32 (
    .out(const_0_32_out)
);
coreir_const #(
    .value(8'h10),
    .width(8)
) const_16_8 (
    .out(const_16_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_ult_inst0_out),
    .in1(EN[0]),
    .out(magma_Bit_and_inst0_out)
);
coreir_ult #(
    .width(8)
) magma_Bits_8_ult_inst0 (
    .in0(S),
    .in1(const_16_8_out),
    .out(magma_Bits_8_ult_inst0_out)
);
wire [31:0] mux_aoi_16_32_inst0_I [15:0];
assign mux_aoi_16_32_inst0_I[15] = I[15];
assign mux_aoi_16_32_inst0_I[14] = I[14];
assign mux_aoi_16_32_inst0_I[13] = I[13];
assign mux_aoi_16_32_inst0_I[12] = I[12];
assign mux_aoi_16_32_inst0_I[11] = I[11];
assign mux_aoi_16_32_inst0_I[10] = I[10];
assign mux_aoi_16_32_inst0_I[9] = I[9];
assign mux_aoi_16_32_inst0_I[8] = I[8];
assign mux_aoi_16_32_inst0_I[7] = I[7];
assign mux_aoi_16_32_inst0_I[6] = I[6];
assign mux_aoi_16_32_inst0_I[5] = I[5];
assign mux_aoi_16_32_inst0_I[4] = I[4];
assign mux_aoi_16_32_inst0_I[3] = I[3];
assign mux_aoi_16_32_inst0_I[2] = I[2];
assign mux_aoi_16_32_inst0_I[1] = I[1];
assign mux_aoi_16_32_inst0_I[0] = I[0];
mux_aoi_16_32 mux_aoi_16_32_inst0 (
    .I(mux_aoi_16_32_inst0_I),
    .O(mux_aoi_16_32_inst0_O),
    .S(S[3:0]),
    .out_sel(mux_aoi_16_32_inst0_out_sel)
);
wire [31:0] mux_aoi_2_32_inst0_I [1:0];
assign mux_aoi_2_32_inst0_I[1] = mux_aoi_16_32_inst0_O;
assign mux_aoi_2_32_inst0_I[0] = const_0_32_out;
mux_aoi_2_32 mux_aoi_2_32_inst0 (
    .I(mux_aoi_2_32_inst0_I),
    .O(mux_aoi_2_32_inst0_O),
    .S(magma_Bit_and_inst0_out),
    .out_sel(mux_aoi_2_32_inst0_out_sel)
);
assign O = mux_aoi_2_32_inst0_O;
endmodule

module MuxWithDefaultWrapper_13_32_8_0 (
    input [31:0] I [12:0],
    input [7:0] S,
    input [0:0] EN,
    output [31:0] O
);
wire [31:0] const_0_32_out;
wire [7:0] const_13_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_ult_inst0_out;
wire [31:0] mux_aoi_13_32_inst0_O;
wire [15:0] mux_aoi_13_32_inst0_out_sel;
wire [31:0] mux_aoi_2_32_inst0_O;
wire [1:0] mux_aoi_2_32_inst0_out_sel;
coreir_const #(
    .value(32'h00000000),
    .width(32)
) const_0_32 (
    .out(const_0_32_out)
);
coreir_const #(
    .value(8'h0d),
    .width(8)
) const_13_8 (
    .out(const_13_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_ult_inst0_out),
    .in1(EN[0]),
    .out(magma_Bit_and_inst0_out)
);
coreir_ult #(
    .width(8)
) magma_Bits_8_ult_inst0 (
    .in0(S),
    .in1(const_13_8_out),
    .out(magma_Bits_8_ult_inst0_out)
);
wire [31:0] mux_aoi_13_32_inst0_I [12:0];
assign mux_aoi_13_32_inst0_I[12] = I[12];
assign mux_aoi_13_32_inst0_I[11] = I[11];
assign mux_aoi_13_32_inst0_I[10] = I[10];
assign mux_aoi_13_32_inst0_I[9] = I[9];
assign mux_aoi_13_32_inst0_I[8] = I[8];
assign mux_aoi_13_32_inst0_I[7] = I[7];
assign mux_aoi_13_32_inst0_I[6] = I[6];
assign mux_aoi_13_32_inst0_I[5] = I[5];
assign mux_aoi_13_32_inst0_I[4] = I[4];
assign mux_aoi_13_32_inst0_I[3] = I[3];
assign mux_aoi_13_32_inst0_I[2] = I[2];
assign mux_aoi_13_32_inst0_I[1] = I[1];
assign mux_aoi_13_32_inst0_I[0] = I[0];
mux_aoi_13_32 mux_aoi_13_32_inst0 (
    .I(mux_aoi_13_32_inst0_I),
    .O(mux_aoi_13_32_inst0_O),
    .S(S[3:0]),
    .out_sel(mux_aoi_13_32_inst0_out_sel)
);
wire [31:0] mux_aoi_2_32_inst0_I [1:0];
assign mux_aoi_2_32_inst0_I[1] = mux_aoi_13_32_inst0_O;
assign mux_aoi_2_32_inst0_I[0] = const_0_32_out;
mux_aoi_2_32 mux_aoi_2_32_inst0 (
    .I(mux_aoi_2_32_inst0_I),
    .O(mux_aoi_2_32_inst0_O),
    .S(magma_Bit_and_inst0_out),
    .out_sel(mux_aoi_2_32_inst0_out_sel)
);
assign O = mux_aoi_2_32_inst0_O;
endmodule

module Chain_2_16 (
  input logic [1:0] accessor_output,
  input logic [1:0] [15:0] chain_data_in,
  input logic chain_en,
  input logic clk_en,
  input logic [1:0] [15:0] curr_tile_data_out,
  input logic flush,
  output logic [1:0] [15:0] data_out_tile
);

always_comb begin
  if (accessor_output[0]) begin
    data_out_tile[0] = curr_tile_data_out[0];
  end
  else if (chain_en) begin
    data_out_tile[0] = chain_data_in[0];
  end
  else data_out_tile[0] = 16'h0;
  if (accessor_output[1]) begin
    data_out_tile[1] = curr_tile_data_out[1];
  end
  else if (chain_en) begin
    data_out_tile[1] = chain_data_in[1];
  end
  else data_out_tile[1] = 16'h0;
end
endmodule   // Chain_2_16

module MemCore_inner (
  input logic [31:0] CONFIG_SPACE_0,
  input logic [31:0] CONFIG_SPACE_1,
  input logic [31:0] CONFIG_SPACE_10,
  input logic [31:0] CONFIG_SPACE_11,
  input logic [31:0] CONFIG_SPACE_12,
  input logic [31:0] CONFIG_SPACE_13,
  input logic [31:0] CONFIG_SPACE_14,
  input logic [31:0] CONFIG_SPACE_15,
  input logic [31:0] CONFIG_SPACE_16,
  input logic [31:0] CONFIG_SPACE_17,
  input logic [31:0] CONFIG_SPACE_18,
  input logic [31:0] CONFIG_SPACE_19,
  input logic [31:0] CONFIG_SPACE_2,
  input logic [31:0] CONFIG_SPACE_20,
  input logic [31:0] CONFIG_SPACE_21,
  input logic [31:0] CONFIG_SPACE_22,
  input logic [31:0] CONFIG_SPACE_23,
  input logic [31:0] CONFIG_SPACE_24,
  input logic [31:0] CONFIG_SPACE_25,
  input logic [31:0] CONFIG_SPACE_26,
  input logic [31:0] CONFIG_SPACE_27,
  input logic [31:0] CONFIG_SPACE_28,
  input logic [31:0] CONFIG_SPACE_29,
  input logic [31:0] CONFIG_SPACE_3,
  input logic [31:0] CONFIG_SPACE_30,
  input logic [31:0] CONFIG_SPACE_31,
  input logic [31:0] CONFIG_SPACE_32,
  input logic [31:0] CONFIG_SPACE_33,
  input logic [31:0] CONFIG_SPACE_34,
  input logic [31:0] CONFIG_SPACE_35,
  input logic [31:0] CONFIG_SPACE_36,
  input logic [31:0] CONFIG_SPACE_37,
  input logic [31:0] CONFIG_SPACE_38,
  input logic [31:0] CONFIG_SPACE_39,
  input logic [31:0] CONFIG_SPACE_4,
  input logic [31:0] CONFIG_SPACE_40,
  input logic [31:0] CONFIG_SPACE_41,
  input logic [31:0] CONFIG_SPACE_42,
  input logic [31:0] CONFIG_SPACE_43,
  input logic [31:0] CONFIG_SPACE_44,
  input logic [18:0] CONFIG_SPACE_45,
  input logic [31:0] CONFIG_SPACE_5,
  input logic [31:0] CONFIG_SPACE_6,
  input logic [31:0] CONFIG_SPACE_7,
  input logic [31:0] CONFIG_SPACE_8,
  input logic [31:0] CONFIG_SPACE_9,
  input logic [0:0] [16:0] MEM_input_width_17_num_0,
  input logic MEM_input_width_17_num_0_valid,
  input logic [0:0] [16:0] MEM_input_width_17_num_1,
  input logic MEM_input_width_17_num_1_valid,
  input logic [0:0] [16:0] MEM_input_width_17_num_2,
  input logic MEM_input_width_17_num_2_valid,
  input logic [0:0] [16:0] MEM_input_width_17_num_3,
  input logic MEM_input_width_17_num_3_valid,
  input logic MEM_input_width_1_num_0,
  input logic MEM_input_width_1_num_1,
  input logic MEM_output_width_17_num_0_ready,
  input logic MEM_output_width_17_num_1_ready,
  input logic MEM_output_width_17_num_2_ready,
  input logic clk,
  input logic clk_en,
  input logic [7:0] config_addr_in,
  input logic [31:0] config_data_in,
  input logic [1:0] config_en,
  input logic config_read,
  input logic config_write,
  input logic flush,
  input logic [1:0] mode,
  input logic mode_excl,
  input logic rst_n,
  input logic tile_en,
  output logic MEM_input_width_17_num_0_ready,
  output logic MEM_input_width_17_num_1_ready,
  output logic MEM_input_width_17_num_2_ready,
  output logic MEM_input_width_17_num_3_ready,
  output logic [0:0] [16:0] MEM_output_width_17_num_0,
  output logic MEM_output_width_17_num_0_valid,
  output logic [0:0] [16:0] MEM_output_width_17_num_1,
  output logic MEM_output_width_17_num_1_valid,
  output logic [0:0] [16:0] MEM_output_width_17_num_2,
  output logic MEM_output_width_17_num_2_valid,
  output logic MEM_output_width_1_num_0,
  output logic MEM_output_width_1_num_1,
  output logic MEM_output_width_1_num_2,
  output logic [1:0] [31:0] config_data_out
);

logic [1458:0] CONFIG_SPACE;
logic [15:0] config_data_in_shrt;
logic [1:0][15:0] config_data_out_shrt;
logic [8:0] config_seq_addr_out;
logic config_seq_clk_en;
logic [0:0][3:0][15:0] config_seq_rd_data_stg;
logic config_seq_ren_out;
logic config_seq_wen_out;
logic [3:0][15:0] config_seq_wr_data;
logic gclk;
logic [0:0][16:0] input_width_17_num_0_fifo_out;
logic input_width_17_num_0_fifo_out_ready;
logic input_width_17_num_0_fifo_out_valid;
logic input_width_17_num_0_input_fifo_empty;
logic input_width_17_num_0_input_fifo_full;
logic [0:0][16:0] input_width_17_num_1_fifo_out;
logic input_width_17_num_1_fifo_out_ready;
logic input_width_17_num_1_fifo_out_valid;
logic input_width_17_num_1_input_fifo_empty;
logic input_width_17_num_1_input_fifo_full;
logic [0:0][16:0] input_width_17_num_2_fifo_out;
logic input_width_17_num_2_fifo_out_ready;
logic input_width_17_num_2_fifo_out_valid;
logic input_width_17_num_2_input_fifo_empty;
logic input_width_17_num_2_input_fifo_full;
logic [0:0][16:0] input_width_17_num_3_fifo_out;
logic input_width_17_num_3_fifo_out_ready;
logic input_width_17_num_3_fifo_out_valid;
logic input_width_17_num_3_input_fifo_empty;
logic input_width_17_num_3_input_fifo_full;
logic mem_ctrl_fiber_access_16_flat_clk;
logic [8:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_addr_to_mem_lifted_lifted;
logic [3:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_buffet_capacity_log_0;
logic [3:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_buffet_capacity_log_1;
logic [3:0][15:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_data_from_mem_lifted_lifted;
logic [3:0][15:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_data_to_mem_lifted_lifted;
logic mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_ren_to_mem_lifted_lifted;
logic mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_tile_en;
logic mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_wen_to_mem_lifted_lifted;
logic mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_block_mode;
logic mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_dense;
logic [15:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_dim_size;
logic mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_do_repeat;
logic [15:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_inner_dim_offset;
logic mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_lookup;
logic [15:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_repeat_factor;
logic mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_repeat_outer_inner_n;
logic mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_root;
logic mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_spacc_mode;
logic [15:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_stop_lvl;
logic mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_tile_en;
logic mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_tile_en;
logic mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_block_mode;
logic mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_compressed;
logic mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_init_blank;
logic mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_lowest_level;
logic mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_spacc_mode;
logic [15:0] mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_stop_lvl;
logic mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_tile_en;
logic [0:0][16:0] mem_ctrl_fiber_access_16_flat_read_scanner_block_rd_out_f_;
logic mem_ctrl_fiber_access_16_flat_read_scanner_block_rd_out_valid_f_;
logic [0:0][16:0] mem_ctrl_fiber_access_16_flat_read_scanner_coord_out_f_;
logic mem_ctrl_fiber_access_16_flat_read_scanner_coord_out_valid_f_;
logic [0:0][16:0] mem_ctrl_fiber_access_16_flat_read_scanner_pos_out_f_;
logic mem_ctrl_fiber_access_16_flat_read_scanner_pos_out_valid_f_;
logic mem_ctrl_fiber_access_16_flat_read_scanner_us_pos_in_ready_f_;
logic mem_ctrl_fiber_access_16_flat_write_scanner_addr_in_ready_f_;
logic mem_ctrl_fiber_access_16_flat_write_scanner_block_wr_in_ready_f_;
logic mem_ctrl_fiber_access_16_flat_write_scanner_data_in_ready_f_;
logic mem_ctrl_stencil_valid_flat_clk;
logic mem_ctrl_stencil_valid_flat_stencil_valid_f_;
logic [3:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality;
logic [10:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0;
logic [10:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1;
logic [10:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2;
logic [10:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3;
logic [10:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4;
logic [10:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5;
logic mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable;
logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr;
logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0;
logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1;
logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2;
logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3;
logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4;
logic [15:0] mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5;
logic mem_ctrl_strg_ram_64_512_delay1_flat_clk;
logic [0:0][16:0] mem_ctrl_strg_ram_64_512_delay1_flat_data_out_f_;
logic mem_ctrl_strg_ram_64_512_delay1_flat_ready_f_;
logic [0:0][8:0] mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_addr_out_lifted;
logic [0:0][3:0][15:0] mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_data_from_strg_lifted;
logic [0:0][3:0][15:0] mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_data_to_strg_lifted;
logic mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_ren_to_strg_lifted;
logic mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_wen_to_strg_lifted;
logic mem_ctrl_strg_ram_64_512_delay1_flat_valid_out_f_;
logic mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_0;
logic mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_1;
logic mem_ctrl_strg_ub_vec_flat_clk;
logic [0:0][16:0] mem_ctrl_strg_ub_vec_flat_data_out_f_0;
logic [0:0][16:0] mem_ctrl_strg_ub_vec_flat_data_out_f_1;
logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_addr_out_lifted;
logic [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr;
logic [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0;
logic [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1;
logic [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2;
logic [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr;
logic [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0;
logic [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1;
logic [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2;
logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2;
logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2;
logic [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2;
logic [2:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2;
logic [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_agg_read_padding;
logic [7:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_agg_read_padding;
logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr;
logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr;
logic [1:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_mode_0;
logic [1:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_mode_1;
logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en;
logic [3:0][15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_data_from_strg_lifted;
logic [3:0][15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_data_to_strg_lifted;
logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_ren_to_strg_lifted;
logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr;
logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0;
logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1;
logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2;
logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3;
logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4;
logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5;
logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr;
logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0;
logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1;
logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2;
logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3;
logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4;
logic [8:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5;
logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable;
logic [9:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5;
logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable;
logic [9:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4;
logic [10:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5;
logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_shared_tb_0;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5;
logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable;
logic [9:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_delay;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5;
logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable;
logic [9:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_delay;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4;
logic [15:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4;
logic [3:0] mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5;
logic mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_wen_to_strg_lifted;
logic memory_0_clk_en;
logic [63:0] memory_0_data_in_p0;
logic [63:0] memory_0_data_out_p0;
logic [8:0] memory_0_read_addr_p0;
logic memory_0_read_enable_p0;
logic [8:0] memory_0_write_addr_p0;
logic memory_0_write_enable_p0;
logic [0:0][16:0] output_width_17_num_0_fifo_in;
logic output_width_17_num_0_fifo_in_ready;
logic output_width_17_num_0_fifo_in_valid;
logic [0:0][16:0] output_width_17_num_0_output_fifo_data_out;
logic output_width_17_num_0_output_fifo_empty;
logic output_width_17_num_0_output_fifo_full;
logic [0:0][16:0] output_width_17_num_1_fifo_in;
logic output_width_17_num_1_fifo_in_ready;
logic output_width_17_num_1_fifo_in_valid;
logic [0:0][16:0] output_width_17_num_1_output_fifo_data_out;
logic output_width_17_num_1_output_fifo_empty;
logic output_width_17_num_1_output_fifo_full;
logic [0:0][16:0] output_width_17_num_2_fifo_in;
logic output_width_17_num_2_fifo_in_ready;
logic output_width_17_num_2_fifo_in_valid;
logic [0:0][16:0] output_width_17_num_2_output_fifo_data_out;
logic output_width_17_num_2_output_fifo_empty;
logic output_width_17_num_2_output_fifo_full;
assign gclk = clk & tile_en;
assign mem_ctrl_fiber_access_16_flat_clk = gclk & (mode == 2'h0);
assign mem_ctrl_strg_ub_vec_flat_clk = gclk & (mode == 2'h1);
assign mem_ctrl_strg_ram_64_512_delay1_flat_clk = gclk & (mode == 2'h2);
assign mem_ctrl_stencil_valid_flat_clk = gclk;
assign input_width_17_num_0_fifo_out_valid = ~input_width_17_num_0_input_fifo_empty;
always_comb begin
  input_width_17_num_0_fifo_out_ready = 1'h1;
  if (mode == 2'h0) begin
    input_width_17_num_0_fifo_out_ready = mem_ctrl_fiber_access_16_flat_read_scanner_us_pos_in_ready_f_;
  end
  else input_width_17_num_0_fifo_out_ready = 1'h1;
end
always_comb begin
  MEM_input_width_17_num_0_ready = 1'h1;
  if (mode == 2'h0) begin
    MEM_input_width_17_num_0_ready = ~input_width_17_num_0_input_fifo_full;
  end
  else if (mode == 2'h1) begin
    MEM_input_width_17_num_0_ready = 1'h1;
  end
  else if (mode == 2'h2) begin
    MEM_input_width_17_num_0_ready = 1'h1;
  end
end
assign input_width_17_num_1_fifo_out_valid = ~input_width_17_num_1_input_fifo_empty;
always_comb begin
  input_width_17_num_1_fifo_out_ready = 1'h1;
  if (mode == 2'h0) begin
    input_width_17_num_1_fifo_out_ready = mem_ctrl_fiber_access_16_flat_write_scanner_addr_in_ready_f_;
  end
  else input_width_17_num_1_fifo_out_ready = 1'h1;
end
always_comb begin
  MEM_input_width_17_num_1_ready = 1'h1;
  if (mode == 2'h0) begin
    MEM_input_width_17_num_1_ready = ~input_width_17_num_1_input_fifo_full;
  end
  else if (mode == 2'h1) begin
    MEM_input_width_17_num_1_ready = 1'h1;
  end
  else if (mode == 2'h2) begin
    MEM_input_width_17_num_1_ready = 1'h1;
  end
end
assign input_width_17_num_2_fifo_out_valid = ~input_width_17_num_2_input_fifo_empty;
always_comb begin
  input_width_17_num_2_fifo_out_ready = 1'h1;
  if (mode == 2'h0) begin
    input_width_17_num_2_fifo_out_ready = mem_ctrl_fiber_access_16_flat_write_scanner_block_wr_in_ready_f_;
  end
  else input_width_17_num_2_fifo_out_ready = 1'h1;
end
always_comb begin
  MEM_input_width_17_num_2_ready = 1'h1;
  if (mode == 2'h0) begin
    MEM_input_width_17_num_2_ready = ~input_width_17_num_2_input_fifo_full;
  end
  else if (mode == 2'h1) begin
    MEM_input_width_17_num_2_ready = 1'h1;
  end
  else if (mode == 2'h2) begin
    MEM_input_width_17_num_2_ready = 1'h1;
  end
end
assign input_width_17_num_3_fifo_out_valid = ~input_width_17_num_3_input_fifo_empty;
always_comb begin
  input_width_17_num_3_fifo_out_ready = 1'h1;
  if (mode == 2'h0) begin
    input_width_17_num_3_fifo_out_ready = mem_ctrl_fiber_access_16_flat_write_scanner_data_in_ready_f_;
  end
  else input_width_17_num_3_fifo_out_ready = 1'h1;
end
always_comb begin
  MEM_input_width_17_num_3_ready = 1'h1;
  if (mode == 2'h0) begin
    MEM_input_width_17_num_3_ready = ~input_width_17_num_3_input_fifo_full;
  end
  else if (mode == 2'h1) begin
    MEM_input_width_17_num_3_ready = 1'h1;
  end
end
assign output_width_17_num_0_fifo_in_ready = ~output_width_17_num_0_output_fifo_full;
always_comb begin
  output_width_17_num_0_fifo_in = 17'h0;
  output_width_17_num_0_fifo_in_valid = 1'h0;
  output_width_17_num_0_fifo_in = mem_ctrl_fiber_access_16_flat_read_scanner_block_rd_out_f_;
  output_width_17_num_0_fifo_in_valid = mem_ctrl_fiber_access_16_flat_read_scanner_block_rd_out_valid_f_;
end
always_comb begin
  MEM_output_width_17_num_0 = 17'h0;
  if (mode == 2'h0) begin
    MEM_output_width_17_num_0 = output_width_17_num_0_output_fifo_data_out;
  end
  else if (mode == 2'h1) begin
    MEM_output_width_17_num_0 = mem_ctrl_strg_ub_vec_flat_data_out_f_0;
  end
  else if (mode == 2'h2) begin
    MEM_output_width_17_num_0 = mem_ctrl_strg_ram_64_512_delay1_flat_data_out_f_;
  end
end
always_comb begin
  MEM_output_width_17_num_0_valid = 1'h0;
  if (mode == 2'h0) begin
    MEM_output_width_17_num_0_valid = ~output_width_17_num_0_output_fifo_empty;
  end
  else if (mode == 2'h1) begin
    MEM_output_width_17_num_0_valid = 1'h1;
  end
  else if (mode == 2'h2) begin
    MEM_output_width_17_num_0_valid = 1'h1;
  end
end
assign output_width_17_num_1_fifo_in_ready = ~output_width_17_num_1_output_fifo_full;
always_comb begin
  output_width_17_num_1_fifo_in = 17'h0;
  output_width_17_num_1_fifo_in_valid = 1'h0;
  output_width_17_num_1_fifo_in = mem_ctrl_fiber_access_16_flat_read_scanner_coord_out_f_;
  output_width_17_num_1_fifo_in_valid = mem_ctrl_fiber_access_16_flat_read_scanner_coord_out_valid_f_;
end
always_comb begin
  MEM_output_width_17_num_1 = 17'h0;
  if (mode == 2'h0) begin
    MEM_output_width_17_num_1 = output_width_17_num_1_output_fifo_data_out;
  end
  else if (mode == 2'h1) begin
    MEM_output_width_17_num_1 = mem_ctrl_strg_ub_vec_flat_data_out_f_1;
  end
end
always_comb begin
  MEM_output_width_17_num_1_valid = 1'h0;
  if (mode == 2'h0) begin
    MEM_output_width_17_num_1_valid = ~output_width_17_num_1_output_fifo_empty;
  end
  else if (mode == 2'h1) begin
    MEM_output_width_17_num_1_valid = 1'h1;
  end
end
assign output_width_17_num_2_fifo_in_ready = ~output_width_17_num_2_output_fifo_full;
always_comb begin
  output_width_17_num_2_fifo_in = 17'h0;
  output_width_17_num_2_fifo_in_valid = 1'h0;
  output_width_17_num_2_fifo_in = mem_ctrl_fiber_access_16_flat_read_scanner_pos_out_f_;
  output_width_17_num_2_fifo_in_valid = mem_ctrl_fiber_access_16_flat_read_scanner_pos_out_valid_f_;
end
always_comb begin
  MEM_output_width_17_num_2 = 17'h0;
  if (mode == 2'h0) begin
    MEM_output_width_17_num_2 = output_width_17_num_2_output_fifo_data_out;
  end
  else MEM_output_width_17_num_2 = 17'h0;
end
always_comb begin
  MEM_output_width_17_num_2_valid = 1'h0;
  if (mode == 2'h0) begin
    MEM_output_width_17_num_2_valid = ~output_width_17_num_2_output_fifo_empty;
  end
  else MEM_output_width_17_num_2_valid = 1'h0;
end
always_comb begin
  MEM_output_width_1_num_0 = 1'h0;
  if (mode == 2'h1) begin
    MEM_output_width_1_num_0 = mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_0;
  end
  else if (mode == 2'h2) begin
    MEM_output_width_1_num_0 = mem_ctrl_strg_ram_64_512_delay1_flat_ready_f_;
  end
end
always_comb begin
  MEM_output_width_1_num_1 = 1'h0;
  if (mode == 2'h1) begin
    MEM_output_width_1_num_1 = mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_1;
  end
  else if (mode == 2'h2) begin
    MEM_output_width_1_num_1 = mem_ctrl_strg_ram_64_512_delay1_flat_valid_out_f_;
  end
end
always_comb begin
  MEM_output_width_1_num_2 = 1'h0;
  if (mode_excl == 1'h1) begin
    MEM_output_width_1_num_2 = mem_ctrl_stencil_valid_flat_stencil_valid_f_;
  end
  else MEM_output_width_1_num_2 = 1'h0;
end
always_comb begin
  memory_0_data_in_p0 = 64'h0;
  memory_0_write_addr_p0 = 9'h0;
  memory_0_write_enable_p0 = 1'h0;
  memory_0_read_addr_p0 = 9'h0;
  memory_0_read_enable_p0 = 1'h0;
  if (|config_en) begin
    memory_0_data_in_p0 = config_seq_wr_data;
    memory_0_write_addr_p0 = config_seq_addr_out;
    memory_0_write_enable_p0 = config_seq_wen_out;
    memory_0_read_addr_p0 = config_seq_addr_out;
    memory_0_read_enable_p0 = config_seq_ren_out;
  end
  else if (mode == 2'h0) begin
    memory_0_data_in_p0 = mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_data_to_mem_lifted_lifted;
    memory_0_write_addr_p0 = mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_addr_to_mem_lifted_lifted;
    memory_0_write_enable_p0 = mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_wen_to_mem_lifted_lifted;
    memory_0_read_addr_p0 = mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_addr_to_mem_lifted_lifted;
    memory_0_read_enable_p0 = mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_ren_to_mem_lifted_lifted;
  end
  else if (mode == 2'h1) begin
    memory_0_data_in_p0 = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_data_to_strg_lifted;
    memory_0_write_addr_p0 = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_addr_out_lifted;
    memory_0_write_enable_p0 = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_wen_to_strg_lifted;
    memory_0_read_addr_p0 = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_addr_out_lifted;
    memory_0_read_enable_p0 = mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_ren_to_strg_lifted;
  end
  else if (mode == 2'h2) begin
    memory_0_data_in_p0 = mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_data_to_strg_lifted;
    memory_0_write_addr_p0 = mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_addr_out_lifted;
    memory_0_write_enable_p0 = mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_wen_to_strg_lifted;
    memory_0_read_addr_p0 = mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_addr_out_lifted;
    memory_0_read_enable_p0 = mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_ren_to_strg_lifted;
  end
end
always_comb begin
  mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_data_from_mem_lifted_lifted = memory_0_data_out_p0;
  mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_data_from_strg_lifted = memory_0_data_out_p0;
  mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_data_from_strg_lifted = memory_0_data_out_p0;
  config_seq_rd_data_stg = memory_0_data_out_p0;
end
assign config_data_in_shrt = config_data_in[15:0];
assign config_data_out[0] = 32'(config_data_out_shrt[0]);
assign config_data_out[1] = 32'(config_data_out_shrt[1]);
assign config_seq_clk_en = clk_en | (|config_en);
assign memory_0_clk_en = clk_en | (|config_en);
assign {mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_buffet_capacity_log_0, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_buffet_capacity_log_1, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_tile_en, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_block_mode, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_dense, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_dim_size, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_do_repeat, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_inner_dim_offset, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_lookup, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_repeat_factor, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_repeat_outer_inner_n, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_root, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_spacc_mode, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_stop_lvl, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_tile_en, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_tile_en, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_block_mode, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_compressed, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_init_blank, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_lowest_level, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_spacc_mode, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_stop_lvl, mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_tile_en} = CONFIG_SPACE[103:0];
assign {mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_agg_read_padding, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_agg_read_padding, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_mode_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_mode_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_shared_tb_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_delay, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_delay, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4, mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5} = CONFIG_SPACE[1275:0];
assign {mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality, mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0, mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1, mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2, mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3, mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4, mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5, mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable, mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr, mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0, mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1, mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2, mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3, mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4, mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5} = CONFIG_SPACE[1458:1276];
assign CONFIG_SPACE[31:0] = CONFIG_SPACE_0;
assign CONFIG_SPACE[63:32] = CONFIG_SPACE_1;
assign CONFIG_SPACE[95:64] = CONFIG_SPACE_2;
assign CONFIG_SPACE[127:96] = CONFIG_SPACE_3;
assign CONFIG_SPACE[159:128] = CONFIG_SPACE_4;
assign CONFIG_SPACE[191:160] = CONFIG_SPACE_5;
assign CONFIG_SPACE[223:192] = CONFIG_SPACE_6;
assign CONFIG_SPACE[255:224] = CONFIG_SPACE_7;
assign CONFIG_SPACE[287:256] = CONFIG_SPACE_8;
assign CONFIG_SPACE[319:288] = CONFIG_SPACE_9;
assign CONFIG_SPACE[351:320] = CONFIG_SPACE_10;
assign CONFIG_SPACE[383:352] = CONFIG_SPACE_11;
assign CONFIG_SPACE[415:384] = CONFIG_SPACE_12;
assign CONFIG_SPACE[447:416] = CONFIG_SPACE_13;
assign CONFIG_SPACE[479:448] = CONFIG_SPACE_14;
assign CONFIG_SPACE[511:480] = CONFIG_SPACE_15;
assign CONFIG_SPACE[543:512] = CONFIG_SPACE_16;
assign CONFIG_SPACE[575:544] = CONFIG_SPACE_17;
assign CONFIG_SPACE[607:576] = CONFIG_SPACE_18;
assign CONFIG_SPACE[639:608] = CONFIG_SPACE_19;
assign CONFIG_SPACE[671:640] = CONFIG_SPACE_20;
assign CONFIG_SPACE[703:672] = CONFIG_SPACE_21;
assign CONFIG_SPACE[735:704] = CONFIG_SPACE_22;
assign CONFIG_SPACE[767:736] = CONFIG_SPACE_23;
assign CONFIG_SPACE[799:768] = CONFIG_SPACE_24;
assign CONFIG_SPACE[831:800] = CONFIG_SPACE_25;
assign CONFIG_SPACE[863:832] = CONFIG_SPACE_26;
assign CONFIG_SPACE[895:864] = CONFIG_SPACE_27;
assign CONFIG_SPACE[927:896] = CONFIG_SPACE_28;
assign CONFIG_SPACE[959:928] = CONFIG_SPACE_29;
assign CONFIG_SPACE[991:960] = CONFIG_SPACE_30;
assign CONFIG_SPACE[1023:992] = CONFIG_SPACE_31;
assign CONFIG_SPACE[1055:1024] = CONFIG_SPACE_32;
assign CONFIG_SPACE[1087:1056] = CONFIG_SPACE_33;
assign CONFIG_SPACE[1119:1088] = CONFIG_SPACE_34;
assign CONFIG_SPACE[1151:1120] = CONFIG_SPACE_35;
assign CONFIG_SPACE[1183:1152] = CONFIG_SPACE_36;
assign CONFIG_SPACE[1215:1184] = CONFIG_SPACE_37;
assign CONFIG_SPACE[1247:1216] = CONFIG_SPACE_38;
assign CONFIG_SPACE[1279:1248] = CONFIG_SPACE_39;
assign CONFIG_SPACE[1311:1280] = CONFIG_SPACE_40;
assign CONFIG_SPACE[1343:1312] = CONFIG_SPACE_41;
assign CONFIG_SPACE[1375:1344] = CONFIG_SPACE_42;
assign CONFIG_SPACE[1407:1376] = CONFIG_SPACE_43;
assign CONFIG_SPACE[1439:1408] = CONFIG_SPACE_44;
assign CONFIG_SPACE[1458:1440] = CONFIG_SPACE_45;
fiber_access_16_flat mem_ctrl_fiber_access_16_flat (
  .clk(mem_ctrl_fiber_access_16_flat_clk),
  .clk_en(clk_en),
  .fiber_access_16_inst_buffet_buffet_capacity_log_0(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_buffet_capacity_log_0),
  .fiber_access_16_inst_buffet_buffet_capacity_log_1(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_buffet_capacity_log_1),
  .fiber_access_16_inst_buffet_data_from_mem_lifted_lifted(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_data_from_mem_lifted_lifted),
  .fiber_access_16_inst_buffet_tile_en(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_tile_en),
  .fiber_access_16_inst_read_scanner_block_mode(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_block_mode),
  .fiber_access_16_inst_read_scanner_dense(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_dense),
  .fiber_access_16_inst_read_scanner_dim_size(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_dim_size),
  .fiber_access_16_inst_read_scanner_do_repeat(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_do_repeat),
  .fiber_access_16_inst_read_scanner_inner_dim_offset(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_inner_dim_offset),
  .fiber_access_16_inst_read_scanner_lookup(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_lookup),
  .fiber_access_16_inst_read_scanner_repeat_factor(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_repeat_factor),
  .fiber_access_16_inst_read_scanner_repeat_outer_inner_n(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_repeat_outer_inner_n),
  .fiber_access_16_inst_read_scanner_root(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_root),
  .fiber_access_16_inst_read_scanner_spacc_mode(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_spacc_mode),
  .fiber_access_16_inst_read_scanner_stop_lvl(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_stop_lvl),
  .fiber_access_16_inst_read_scanner_tile_en(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_read_scanner_tile_en),
  .fiber_access_16_inst_tile_en(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_tile_en),
  .fiber_access_16_inst_write_scanner_block_mode(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_block_mode),
  .fiber_access_16_inst_write_scanner_compressed(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_compressed),
  .fiber_access_16_inst_write_scanner_init_blank(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_init_blank),
  .fiber_access_16_inst_write_scanner_lowest_level(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_lowest_level),
  .fiber_access_16_inst_write_scanner_spacc_mode(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_spacc_mode),
  .fiber_access_16_inst_write_scanner_stop_lvl(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_stop_lvl),
  .fiber_access_16_inst_write_scanner_tile_en(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_write_scanner_tile_en),
  .flush(flush),
  .read_scanner_block_rd_out_ready_f_(output_width_17_num_0_fifo_in_ready),
  .read_scanner_coord_out_ready_f_(output_width_17_num_1_fifo_in_ready),
  .read_scanner_pos_out_ready_f_(output_width_17_num_2_fifo_in_ready),
  .read_scanner_us_pos_in_f_(input_width_17_num_0_fifo_out),
  .read_scanner_us_pos_in_valid_f_(input_width_17_num_0_fifo_out_valid),
  .rst_n(rst_n),
  .write_scanner_addr_in_f_(input_width_17_num_1_fifo_out),
  .write_scanner_addr_in_valid_f_(input_width_17_num_1_fifo_out_valid),
  .write_scanner_block_wr_in_f_(input_width_17_num_2_fifo_out),
  .write_scanner_block_wr_in_valid_f_(input_width_17_num_2_fifo_out_valid),
  .write_scanner_data_in_f_(input_width_17_num_3_fifo_out),
  .write_scanner_data_in_valid_f_(input_width_17_num_3_fifo_out_valid),
  .fiber_access_16_inst_buffet_addr_to_mem_lifted_lifted(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_addr_to_mem_lifted_lifted),
  .fiber_access_16_inst_buffet_data_to_mem_lifted_lifted(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_data_to_mem_lifted_lifted),
  .fiber_access_16_inst_buffet_ren_to_mem_lifted_lifted(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_ren_to_mem_lifted_lifted),
  .fiber_access_16_inst_buffet_wen_to_mem_lifted_lifted(mem_ctrl_fiber_access_16_flat_fiber_access_16_inst_buffet_wen_to_mem_lifted_lifted),
  .read_scanner_block_rd_out_f_(mem_ctrl_fiber_access_16_flat_read_scanner_block_rd_out_f_),
  .read_scanner_block_rd_out_valid_f_(mem_ctrl_fiber_access_16_flat_read_scanner_block_rd_out_valid_f_),
  .read_scanner_coord_out_f_(mem_ctrl_fiber_access_16_flat_read_scanner_coord_out_f_),
  .read_scanner_coord_out_valid_f_(mem_ctrl_fiber_access_16_flat_read_scanner_coord_out_valid_f_),
  .read_scanner_pos_out_f_(mem_ctrl_fiber_access_16_flat_read_scanner_pos_out_f_),
  .read_scanner_pos_out_valid_f_(mem_ctrl_fiber_access_16_flat_read_scanner_pos_out_valid_f_),
  .read_scanner_us_pos_in_ready_f_(mem_ctrl_fiber_access_16_flat_read_scanner_us_pos_in_ready_f_),
  .write_scanner_addr_in_ready_f_(mem_ctrl_fiber_access_16_flat_write_scanner_addr_in_ready_f_),
  .write_scanner_block_wr_in_ready_f_(mem_ctrl_fiber_access_16_flat_write_scanner_block_wr_in_ready_f_),
  .write_scanner_data_in_ready_f_(mem_ctrl_fiber_access_16_flat_write_scanner_data_in_ready_f_)
);

strg_ub_vec_flat mem_ctrl_strg_ub_vec_flat (
  .chain_data_in_f_0(MEM_input_width_17_num_0),
  .chain_data_in_f_1(MEM_input_width_17_num_1),
  .clk(mem_ctrl_strg_ub_vec_flat_clk),
  .clk_en(clk_en),
  .data_in_f_0(MEM_input_width_17_num_2),
  .data_in_f_1(MEM_input_width_17_num_3),
  .flush(flush),
  .rst_n(rst_n),
  .strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr),
  .strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0),
  .strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1),
  .strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2),
  .strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr),
  .strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0),
  .strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1),
  .strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2),
  .strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable),
  .strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr),
  .strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0),
  .strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1),
  .strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2),
  .strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable),
  .strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr),
  .strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0),
  .strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1),
  .strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2),
  .strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality),
  .strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0),
  .strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1),
  .strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2),
  .strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality),
  .strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0),
  .strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1),
  .strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2),
  .strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_agg_read_padding(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_agg_read_padding),
  .strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_agg_read_padding(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_agg_read_padding),
  .strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr),
  .strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr),
  .strg_ub_vec_inst_agg_sram_shared_mode_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_mode_0),
  .strg_ub_vec_inst_agg_sram_shared_mode_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_agg_sram_shared_mode_1),
  .strg_ub_vec_inst_chain_chain_en(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_chain_chain_en),
  .strg_ub_vec_inst_data_from_strg_lifted(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_data_from_strg_lifted),
  .strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr),
  .strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0),
  .strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1),
  .strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2),
  .strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3),
  .strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4),
  .strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5),
  .strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr),
  .strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0),
  .strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1),
  .strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2),
  .strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3),
  .strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4),
  .strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5),
  .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality),
  .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0),
  .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1),
  .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2),
  .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3),
  .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4),
  .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5),
  .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality),
  .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0),
  .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1),
  .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2),
  .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3),
  .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4),
  .strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4),
  .strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5),
  .strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality),
  .strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0),
  .strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1),
  .strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2),
  .strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3),
  .strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4),
  .strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5),
  .strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality),
  .strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0),
  .strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1),
  .strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2),
  .strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3),
  .strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4),
  .strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5),
  .strg_ub_vec_inst_tb_only_shared_tb_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_shared_tb_0),
  .strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr),
  .strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0),
  .strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1),
  .strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2),
  .strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3),
  .strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4),
  .strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5),
  .strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr),
  .strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0),
  .strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1),
  .strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2),
  .strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3),
  .strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4),
  .strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_delay(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_delay),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_delay(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_delay),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4),
  .strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5),
  .strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr),
  .strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0),
  .strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1),
  .strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2),
  .strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3),
  .strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4),
  .strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5),
  .strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr),
  .strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0),
  .strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1),
  .strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2),
  .strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3),
  .strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4),
  .strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5),
  .accessor_output_f_b_0(mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_0),
  .accessor_output_f_b_1(mem_ctrl_strg_ub_vec_flat_accessor_output_f_b_1),
  .data_out_f_0(mem_ctrl_strg_ub_vec_flat_data_out_f_0),
  .data_out_f_1(mem_ctrl_strg_ub_vec_flat_data_out_f_1),
  .strg_ub_vec_inst_addr_out_lifted(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_addr_out_lifted),
  .strg_ub_vec_inst_data_to_strg_lifted(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_data_to_strg_lifted),
  .strg_ub_vec_inst_ren_to_strg_lifted(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_ren_to_strg_lifted),
  .strg_ub_vec_inst_wen_to_strg_lifted(mem_ctrl_strg_ub_vec_flat_strg_ub_vec_inst_wen_to_strg_lifted)
);

strg_ram_64_512_delay1_flat mem_ctrl_strg_ram_64_512_delay1_flat (
  .clk(mem_ctrl_strg_ram_64_512_delay1_flat_clk),
  .clk_en(clk_en),
  .data_in_f_(MEM_input_width_17_num_0),
  .flush(flush),
  .rd_addr_in_f_(MEM_input_width_17_num_1),
  .ren_f_(MEM_input_width_1_num_0),
  .rst_n(rst_n),
  .strg_ram_64_512_delay1_inst_data_from_strg_lifted(mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_data_from_strg_lifted),
  .wen_f_(MEM_input_width_1_num_1),
  .wr_addr_in_f_(MEM_input_width_17_num_2),
  .data_out_f_(mem_ctrl_strg_ram_64_512_delay1_flat_data_out_f_),
  .ready_f_(mem_ctrl_strg_ram_64_512_delay1_flat_ready_f_),
  .strg_ram_64_512_delay1_inst_addr_out_lifted(mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_addr_out_lifted),
  .strg_ram_64_512_delay1_inst_data_to_strg_lifted(mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_data_to_strg_lifted),
  .strg_ram_64_512_delay1_inst_ren_to_strg_lifted(mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_ren_to_strg_lifted),
  .strg_ram_64_512_delay1_inst_wen_to_strg_lifted(mem_ctrl_strg_ram_64_512_delay1_flat_strg_ram_64_512_delay1_inst_wen_to_strg_lifted),
  .valid_out_f_(mem_ctrl_strg_ram_64_512_delay1_flat_valid_out_f_)
);

stencil_valid_flat mem_ctrl_stencil_valid_flat (
  .clk(mem_ctrl_stencil_valid_flat_clk),
  .clk_en(clk_en),
  .flush(flush),
  .rst_n(rst_n),
  .stencil_valid_inst_loops_stencil_valid_dimensionality(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_dimensionality),
  .stencil_valid_inst_loops_stencil_valid_ranges_0(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_0),
  .stencil_valid_inst_loops_stencil_valid_ranges_1(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_1),
  .stencil_valid_inst_loops_stencil_valid_ranges_2(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_2),
  .stencil_valid_inst_loops_stencil_valid_ranges_3(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_3),
  .stencil_valid_inst_loops_stencil_valid_ranges_4(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_4),
  .stencil_valid_inst_loops_stencil_valid_ranges_5(mem_ctrl_stencil_valid_flat_stencil_valid_inst_loops_stencil_valid_ranges_5),
  .stencil_valid_inst_stencil_valid_sched_gen_enable(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_enable),
  .stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr),
  .stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0),
  .stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1),
  .stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2),
  .stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3),
  .stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4),
  .stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5(mem_ctrl_stencil_valid_flat_stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5),
  .stencil_valid_f_(mem_ctrl_stencil_valid_flat_stencil_valid_f_)
);

reg_fifo_depth_2_w_17_afd_2 input_width_17_num_0_input_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(MEM_input_width_17_num_0),
  .flush(flush),
  .pop(input_width_17_num_0_fifo_out_ready),
  .push(MEM_input_width_17_num_0_valid),
  .rst_n(rst_n),
  .data_out(input_width_17_num_0_fifo_out),
  .empty(input_width_17_num_0_input_fifo_empty),
  .full(input_width_17_num_0_input_fifo_full)
);

reg_fifo_depth_2_w_17_afd_2 input_width_17_num_1_input_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(MEM_input_width_17_num_1),
  .flush(flush),
  .pop(input_width_17_num_1_fifo_out_ready),
  .push(MEM_input_width_17_num_1_valid),
  .rst_n(rst_n),
  .data_out(input_width_17_num_1_fifo_out),
  .empty(input_width_17_num_1_input_fifo_empty),
  .full(input_width_17_num_1_input_fifo_full)
);

reg_fifo_depth_2_w_17_afd_2 input_width_17_num_2_input_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(MEM_input_width_17_num_2),
  .flush(flush),
  .pop(input_width_17_num_2_fifo_out_ready),
  .push(MEM_input_width_17_num_2_valid),
  .rst_n(rst_n),
  .data_out(input_width_17_num_2_fifo_out),
  .empty(input_width_17_num_2_input_fifo_empty),
  .full(input_width_17_num_2_input_fifo_full)
);

reg_fifo_depth_2_w_17_afd_2 input_width_17_num_3_input_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(MEM_input_width_17_num_3),
  .flush(flush),
  .pop(input_width_17_num_3_fifo_out_ready),
  .push(MEM_input_width_17_num_3_valid),
  .rst_n(rst_n),
  .data_out(input_width_17_num_3_fifo_out),
  .empty(input_width_17_num_3_input_fifo_empty),
  .full(input_width_17_num_3_input_fifo_full)
);

reg_fifo_depth_2_w_17_afd_2 output_width_17_num_0_output_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(output_width_17_num_0_fifo_in),
  .flush(flush),
  .pop(MEM_output_width_17_num_0_ready),
  .push(output_width_17_num_0_fifo_in_valid),
  .rst_n(rst_n),
  .data_out(output_width_17_num_0_output_fifo_data_out),
  .empty(output_width_17_num_0_output_fifo_empty),
  .full(output_width_17_num_0_output_fifo_full)
);

reg_fifo_depth_2_w_17_afd_2 output_width_17_num_1_output_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(output_width_17_num_1_fifo_in),
  .flush(flush),
  .pop(MEM_output_width_17_num_1_ready),
  .push(output_width_17_num_1_fifo_in_valid),
  .rst_n(rst_n),
  .data_out(output_width_17_num_1_output_fifo_data_out),
  .empty(output_width_17_num_1_output_fifo_empty),
  .full(output_width_17_num_1_output_fifo_full)
);

reg_fifo_depth_2_w_17_afd_2 output_width_17_num_2_output_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(output_width_17_num_2_fifo_in),
  .flush(flush),
  .pop(MEM_output_width_17_num_2_ready),
  .push(output_width_17_num_2_fifo_in_valid),
  .rst_n(rst_n),
  .data_out(output_width_17_num_2_output_fifo_data_out),
  .empty(output_width_17_num_2_output_fifo_empty),
  .full(output_width_17_num_2_output_fifo_full)
);

sram_sp__0 memory_0 (
  .clk(gclk),
  .clk_en(memory_0_clk_en),
  .data_in_p0(memory_0_data_in_p0),
  .flush(flush),
  .read_addr_p0(memory_0_read_addr_p0),
  .read_enable_p0(memory_0_read_enable_p0),
  .write_addr_p0(memory_0_write_addr_p0),
  .write_enable_p0(memory_0_write_enable_p0),
  .data_out_p0(memory_0_data_out_p0)
);

storage_config_seq_2_64_16 config_seq (
  .clk(gclk),
  .clk_en(config_seq_clk_en),
  .config_addr_in(config_addr_in),
  .config_data_in(config_data_in_shrt),
  .config_en(config_en),
  .config_rd(config_read),
  .config_wr(config_write),
  .flush(flush),
  .rd_data_stg(config_seq_rd_data_stg),
  .rst_n(rst_n),
  .addr_out(config_seq_addr_out),
  .rd_data_out(config_data_out_shrt),
  .ren_out(config_seq_ren_out),
  .wen_out(config_seq_wen_out),
  .wr_data(config_seq_wr_data)
);

endmodule   // MemCore_inner

module MemCore_inner_W (
  input logic [31:0] CONFIG_SPACE_0,
  input logic [31:0] CONFIG_SPACE_1,
  input logic [31:0] CONFIG_SPACE_10,
  input logic [31:0] CONFIG_SPACE_11,
  input logic [31:0] CONFIG_SPACE_12,
  input logic [31:0] CONFIG_SPACE_13,
  input logic [31:0] CONFIG_SPACE_14,
  input logic [31:0] CONFIG_SPACE_15,
  input logic [31:0] CONFIG_SPACE_16,
  input logic [31:0] CONFIG_SPACE_17,
  input logic [31:0] CONFIG_SPACE_18,
  input logic [31:0] CONFIG_SPACE_19,
  input logic [31:0] CONFIG_SPACE_2,
  input logic [31:0] CONFIG_SPACE_20,
  input logic [31:0] CONFIG_SPACE_21,
  input logic [31:0] CONFIG_SPACE_22,
  input logic [31:0] CONFIG_SPACE_23,
  input logic [31:0] CONFIG_SPACE_24,
  input logic [31:0] CONFIG_SPACE_25,
  input logic [31:0] CONFIG_SPACE_26,
  input logic [31:0] CONFIG_SPACE_27,
  input logic [31:0] CONFIG_SPACE_28,
  input logic [31:0] CONFIG_SPACE_29,
  input logic [31:0] CONFIG_SPACE_3,
  input logic [31:0] CONFIG_SPACE_30,
  input logic [31:0] CONFIG_SPACE_31,
  input logic [31:0] CONFIG_SPACE_32,
  input logic [31:0] CONFIG_SPACE_33,
  input logic [31:0] CONFIG_SPACE_34,
  input logic [31:0] CONFIG_SPACE_35,
  input logic [31:0] CONFIG_SPACE_36,
  input logic [31:0] CONFIG_SPACE_37,
  input logic [31:0] CONFIG_SPACE_38,
  input logic [31:0] CONFIG_SPACE_39,
  input logic [31:0] CONFIG_SPACE_4,
  input logic [31:0] CONFIG_SPACE_40,
  input logic [31:0] CONFIG_SPACE_41,
  input logic [31:0] CONFIG_SPACE_42,
  input logic [31:0] CONFIG_SPACE_43,
  input logic [31:0] CONFIG_SPACE_44,
  input logic [18:0] CONFIG_SPACE_45,
  input logic [31:0] CONFIG_SPACE_5,
  input logic [31:0] CONFIG_SPACE_6,
  input logic [31:0] CONFIG_SPACE_7,
  input logic [31:0] CONFIG_SPACE_8,
  input logic [31:0] CONFIG_SPACE_9,
  input logic [0:0] [16:0] MEM_input_width_17_num_0,
  input logic MEM_input_width_17_num_0_valid,
  input logic [0:0] [16:0] MEM_input_width_17_num_1,
  input logic MEM_input_width_17_num_1_valid,
  input logic [0:0] [16:0] MEM_input_width_17_num_2,
  input logic MEM_input_width_17_num_2_valid,
  input logic [0:0] [16:0] MEM_input_width_17_num_3,
  input logic MEM_input_width_17_num_3_valid,
  input logic MEM_input_width_1_num_0,
  input logic MEM_input_width_1_num_1,
  input logic MEM_output_width_17_num_0_ready,
  input logic MEM_output_width_17_num_1_ready,
  input logic MEM_output_width_17_num_2_ready,
  input logic clk,
  input logic clk_en,
  input logic [7:0] config_addr_in,
  input logic [31:0] config_data_in,
  input logic [1:0] config_en,
  input logic config_read,
  input logic config_write,
  input logic flush,
  input logic [1:0] mode,
  input logic mode_excl,
  input logic rst_n,
  input logic tile_en,
  output logic MEM_input_width_17_num_0_ready,
  output logic MEM_input_width_17_num_1_ready,
  output logic MEM_input_width_17_num_2_ready,
  output logic MEM_input_width_17_num_3_ready,
  output logic [0:0] [16:0] MEM_output_width_17_num_0,
  output logic MEM_output_width_17_num_0_valid,
  output logic [0:0] [16:0] MEM_output_width_17_num_1,
  output logic MEM_output_width_17_num_1_valid,
  output logic [0:0] [16:0] MEM_output_width_17_num_2,
  output logic MEM_output_width_17_num_2_valid,
  output logic MEM_output_width_1_num_0,
  output logic MEM_output_width_1_num_1,
  output logic MEM_output_width_1_num_2,
  output logic [31:0] config_data_out_0,
  output logic [31:0] config_data_out_1
);

logic [1:0][31:0] MemCore_inner_config_data_out;
assign config_data_out_0 = MemCore_inner_config_data_out[0];
assign config_data_out_1 = MemCore_inner_config_data_out[1];
MemCore_inner MemCore_inner (
  .CONFIG_SPACE_0(CONFIG_SPACE_0),
  .CONFIG_SPACE_1(CONFIG_SPACE_1),
  .CONFIG_SPACE_10(CONFIG_SPACE_10),
  .CONFIG_SPACE_11(CONFIG_SPACE_11),
  .CONFIG_SPACE_12(CONFIG_SPACE_12),
  .CONFIG_SPACE_13(CONFIG_SPACE_13),
  .CONFIG_SPACE_14(CONFIG_SPACE_14),
  .CONFIG_SPACE_15(CONFIG_SPACE_15),
  .CONFIG_SPACE_16(CONFIG_SPACE_16),
  .CONFIG_SPACE_17(CONFIG_SPACE_17),
  .CONFIG_SPACE_18(CONFIG_SPACE_18),
  .CONFIG_SPACE_19(CONFIG_SPACE_19),
  .CONFIG_SPACE_2(CONFIG_SPACE_2),
  .CONFIG_SPACE_20(CONFIG_SPACE_20),
  .CONFIG_SPACE_21(CONFIG_SPACE_21),
  .CONFIG_SPACE_22(CONFIG_SPACE_22),
  .CONFIG_SPACE_23(CONFIG_SPACE_23),
  .CONFIG_SPACE_24(CONFIG_SPACE_24),
  .CONFIG_SPACE_25(CONFIG_SPACE_25),
  .CONFIG_SPACE_26(CONFIG_SPACE_26),
  .CONFIG_SPACE_27(CONFIG_SPACE_27),
  .CONFIG_SPACE_28(CONFIG_SPACE_28),
  .CONFIG_SPACE_29(CONFIG_SPACE_29),
  .CONFIG_SPACE_3(CONFIG_SPACE_3),
  .CONFIG_SPACE_30(CONFIG_SPACE_30),
  .CONFIG_SPACE_31(CONFIG_SPACE_31),
  .CONFIG_SPACE_32(CONFIG_SPACE_32),
  .CONFIG_SPACE_33(CONFIG_SPACE_33),
  .CONFIG_SPACE_34(CONFIG_SPACE_34),
  .CONFIG_SPACE_35(CONFIG_SPACE_35),
  .CONFIG_SPACE_36(CONFIG_SPACE_36),
  .CONFIG_SPACE_37(CONFIG_SPACE_37),
  .CONFIG_SPACE_38(CONFIG_SPACE_38),
  .CONFIG_SPACE_39(CONFIG_SPACE_39),
  .CONFIG_SPACE_4(CONFIG_SPACE_4),
  .CONFIG_SPACE_40(CONFIG_SPACE_40),
  .CONFIG_SPACE_41(CONFIG_SPACE_41),
  .CONFIG_SPACE_42(CONFIG_SPACE_42),
  .CONFIG_SPACE_43(CONFIG_SPACE_43),
  .CONFIG_SPACE_44(CONFIG_SPACE_44),
  .CONFIG_SPACE_45(CONFIG_SPACE_45),
  .CONFIG_SPACE_5(CONFIG_SPACE_5),
  .CONFIG_SPACE_6(CONFIG_SPACE_6),
  .CONFIG_SPACE_7(CONFIG_SPACE_7),
  .CONFIG_SPACE_8(CONFIG_SPACE_8),
  .CONFIG_SPACE_9(CONFIG_SPACE_9),
  .MEM_input_width_17_num_0(MEM_input_width_17_num_0),
  .MEM_input_width_17_num_0_valid(MEM_input_width_17_num_0_valid),
  .MEM_input_width_17_num_1(MEM_input_width_17_num_1),
  .MEM_input_width_17_num_1_valid(MEM_input_width_17_num_1_valid),
  .MEM_input_width_17_num_2(MEM_input_width_17_num_2),
  .MEM_input_width_17_num_2_valid(MEM_input_width_17_num_2_valid),
  .MEM_input_width_17_num_3(MEM_input_width_17_num_3),
  .MEM_input_width_17_num_3_valid(MEM_input_width_17_num_3_valid),
  .MEM_input_width_1_num_0(MEM_input_width_1_num_0),
  .MEM_input_width_1_num_1(MEM_input_width_1_num_1),
  .MEM_output_width_17_num_0_ready(MEM_output_width_17_num_0_ready),
  .MEM_output_width_17_num_1_ready(MEM_output_width_17_num_1_ready),
  .MEM_output_width_17_num_2_ready(MEM_output_width_17_num_2_ready),
  .clk(clk),
  .clk_en(clk_en),
  .config_addr_in(config_addr_in),
  .config_data_in(config_data_in),
  .config_en(config_en),
  .config_read(config_read),
  .config_write(config_write),
  .flush(flush),
  .mode(mode),
  .mode_excl(mode_excl),
  .rst_n(rst_n),
  .tile_en(tile_en),
  .MEM_input_width_17_num_0_ready(MEM_input_width_17_num_0_ready),
  .MEM_input_width_17_num_1_ready(MEM_input_width_17_num_1_ready),
  .MEM_input_width_17_num_2_ready(MEM_input_width_17_num_2_ready),
  .MEM_input_width_17_num_3_ready(MEM_input_width_17_num_3_ready),
  .MEM_output_width_17_num_0(MEM_output_width_17_num_0),
  .MEM_output_width_17_num_0_valid(MEM_output_width_17_num_0_valid),
  .MEM_output_width_17_num_1(MEM_output_width_17_num_1),
  .MEM_output_width_17_num_1_valid(MEM_output_width_17_num_1_valid),
  .MEM_output_width_17_num_2(MEM_output_width_17_num_2),
  .MEM_output_width_17_num_2_valid(MEM_output_width_17_num_2_valid),
  .MEM_output_width_1_num_0(MEM_output_width_1_num_0),
  .MEM_output_width_1_num_1(MEM_output_width_1_num_1),
  .MEM_output_width_1_num_2(MEM_output_width_1_num_2),
  .config_data_out(MemCore_inner_config_data_out)
);

endmodule   // MemCore_inner_W

module addr_gen_3_16 (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [1:0] mux_sel,
  input logic restart,
  input logic rst_n,
  input logic [15:0] starting_addr,
  input logic step,
  input logic [2:0] [15:0] strides,
  output logic [15:0] addr_out
);

logic [15:0] calc_addr;
logic [15:0] current_addr;
logic [15:0] strt_addr;
assign strt_addr = starting_addr;
assign addr_out = calc_addr;
assign calc_addr = current_addr;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    current_addr <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      current_addr <= strt_addr;
    end
    else if (step) begin
      if (restart) begin
        current_addr <= strt_addr;
      end
      else current_addr <= current_addr + strides[mux_sel];
    end
  end
end
endmodule   // addr_gen_3_16

module addr_gen_3_3 (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [1:0] mux_sel,
  input logic restart,
  input logic rst_n,
  input logic [2:0] starting_addr,
  input logic step,
  input logic [2:0] [2:0] strides,
  output logic [2:0] addr_out
);

logic [2:0] calc_addr;
logic [2:0] current_addr;
logic [2:0] strt_addr;
assign strt_addr = starting_addr;
assign addr_out = calc_addr;
assign calc_addr = current_addr;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    current_addr <= 3'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      current_addr <= strt_addr;
    end
    else if (step) begin
      if (restart) begin
        current_addr <= strt_addr;
      end
      else current_addr <= current_addr + strides[mux_sel];
    end
  end
end
endmodule   // addr_gen_3_3

module addr_gen_6_16 (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [2:0] mux_sel,
  input logic restart,
  input logic rst_n,
  input logic [15:0] starting_addr,
  input logic step,
  input logic [5:0] [15:0] strides,
  output logic [15:0] addr_out
);

logic [15:0] calc_addr;
logic [15:0] current_addr;
logic [15:0] strt_addr;
assign strt_addr = starting_addr;
assign addr_out = calc_addr;
assign calc_addr = current_addr;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    current_addr <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      current_addr <= strt_addr;
    end
    else if (step) begin
      if (restart) begin
        current_addr <= strt_addr;
      end
      else current_addr <= current_addr + strides[mux_sel];
    end
  end
end
endmodule   // addr_gen_6_16

module addr_gen_6_16_delay_addr_10 (
  input logic clk,
  input logic clk_en,
  input logic [9:0] delay,
  input logic flush,
  input logic [2:0] mux_sel,
  input logic restart,
  input logic rst_n,
  input logic [15:0] starting_addr,
  input logic step,
  input logic [5:0] [15:0] strides,
  output logic [15:0] addr_out,
  output logic [9:0] delay_out,
  output logic [15:0] delayed_addr_out
);

logic [15:0] calc_addr;
logic [15:0] current_addr;
logic [15:0] strt_addr;
assign delay_out = delay;
assign strt_addr = starting_addr;
assign addr_out = calc_addr;
assign calc_addr = current_addr;
assign delayed_addr_out = current_addr + 16'(delay);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    current_addr <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      current_addr <= strt_addr;
    end
    else if (step) begin
      if (restart) begin
        current_addr <= strt_addr;
      end
      else current_addr <= current_addr + strides[mux_sel];
    end
  end
end
endmodule   // addr_gen_6_16_delay_addr_10

module addr_gen_6_4 (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [2:0] mux_sel,
  input logic restart,
  input logic rst_n,
  input logic [3:0] starting_addr,
  input logic step,
  input logic [5:0] [3:0] strides,
  output logic [3:0] addr_out
);

logic [3:0] calc_addr;
logic [3:0] current_addr;
logic [3:0] strt_addr;
assign strt_addr = starting_addr;
assign addr_out = calc_addr;
assign calc_addr = current_addr;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    current_addr <= 4'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      current_addr <= strt_addr;
    end
    else if (step) begin
      if (restart) begin
        current_addr <= strt_addr;
      end
      else current_addr <= current_addr + strides[mux_sel];
    end
  end
end
endmodule   // addr_gen_6_4

module addr_gen_6_9 (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [2:0] mux_sel,
  input logic restart,
  input logic rst_n,
  input logic [8:0] starting_addr,
  input logic step,
  input logic [5:0] [8:0] strides,
  output logic [8:0] addr_out
);

logic [8:0] calc_addr;
logic [8:0] current_addr;
logic [8:0] strt_addr;
assign strt_addr = starting_addr;
assign addr_out = calc_addr;
assign calc_addr = current_addr;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    current_addr <= 9'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      current_addr <= strt_addr;
    end
    else if (step) begin
      if (restart) begin
        current_addr <= strt_addr;
      end
      else current_addr <= current_addr + strides[mux_sel];
    end
  end
end
endmodule   // addr_gen_6_9

module agg_sram_shared_addr_gen (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [1:0] mode,
  input logic rst_n,
  input logic [1:0] sram_read,
  input logic [1:0] [8:0] sram_read_addr,
  input logic [8:0] starting_addr,
  input logic step,
  output logic [8:0] addr_out
);

logic [3:0][8:0] addr_fifo;
logic [8:0] addr_fifo_in;
logic [8:0] addr_fifo_out;
logic addr_fifo_wr_en;
logic [8:0] lin_addr_cnter;
logic [1:0] rd_ptr;
logic [1:0] wr_ptr;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    lin_addr_cnter <= 9'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      lin_addr_cnter <= 9'h0;
    end
    else if (mode[1] == 1'h0) begin
      if (step) begin
        if (lin_addr_cnter == 9'h1FF) begin
          lin_addr_cnter <= 9'h0;
        end
        else lin_addr_cnter <= lin_addr_cnter + 9'h1;
      end
    end
  end
end
assign addr_fifo_wr_en = mode[0] ? sram_read[1]: sram_read[0];
assign addr_fifo_in = mode[0] ? sram_read_addr[1]: sram_read_addr[0];

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    wr_ptr <= 2'h0;
    rd_ptr <= 2'h0;
    addr_fifo <= 36'h0;
    addr_fifo_out <= 9'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      wr_ptr <= 2'h0;
      rd_ptr <= 2'h0;
      addr_fifo <= 36'h0;
      addr_fifo_out <= 9'h0;
    end
    else if (mode[1] == 1'h1) begin
      if (addr_fifo_wr_en) begin
        wr_ptr <= wr_ptr + 2'h1;
        addr_fifo[wr_ptr] <= addr_fifo_in;
      end
      if (step) begin
        rd_ptr <= rd_ptr + 2'h1;
      end
      addr_fifo_out <= addr_fifo[rd_ptr];
    end
  end
end
assign addr_out = mode[1] ? addr_fifo_out: lin_addr_cnter + starting_addr;
endmodule   // agg_sram_shared_addr_gen

module agg_sram_shared_sched_gen (
  input logic [7:0] agg_read_padding,
  input logic agg_write,
  input logic [1:0] agg_write_addr_l2b,
  input logic [2:0] agg_write_mux_sel,
  input logic agg_write_restart,
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [1:0] mode,
  input logic rst_n,
  input logic [1:0] sram_read_d,
  output logic valid_output
);

logic agg_write_4_r;
logic [7:0] pad_cnt;
logic pad_cnt_en;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    agg_write_4_r <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      agg_write_4_r <= 1'h0;
    end
    else if (mode[1] == 1'h0) begin
      agg_write_4_r <= agg_write & (&agg_write_addr_l2b);
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    pad_cnt_en <= 1'h0;
    pad_cnt <= 8'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      pad_cnt_en <= 1'h0;
      pad_cnt <= 8'h0;
    end
    else if ((mode[1] == 1'h0) & (agg_read_padding != 8'h0)) begin
      if (agg_write & ((agg_write_mux_sel != 3'h0) | agg_write_restart)) begin
        pad_cnt_en <= 1'h1;
      end
      else if (pad_cnt == agg_read_padding) begin
        pad_cnt_en <= 1'h0;
      end
      if (pad_cnt == agg_read_padding) begin
        pad_cnt <= 8'h0;
      end
      else if (pad_cnt_en | (agg_write & ((agg_write_mux_sel != 3'h0) | agg_write_restart))) begin
        pad_cnt <= pad_cnt + 8'h1;
      end
    end
  end
end
always_comb begin
  if (mode[1] == 1'h0) begin
    if (agg_read_padding != 8'h0) begin
      valid_output = (agg_read_padding == pad_cnt) | agg_write_4_r;
    end
    else valid_output = agg_write_4_r;
  end
  else valid_output = mode[0] ? sram_read_d[1]: sram_read_d[0];
end
endmodule   // agg_sram_shared_sched_gen

module arbiter_2_in_RR_algo (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [1:0] request_in,
  input logic resource_ready,
  input logic rst_n,
  output logic [1:0] grant_out
);

logic [1:0] grant_line;
logic [1:0] grant_line_ready;
logic [1:0] grant_out_consolation;
logic [1:0] grant_out_priority;
logic tmp_done;
logic tmp_out_first;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    grant_line <= 2'h1;
  end
  else if (clk_en) begin
    if (flush) begin
      grant_line <= 2'h1;
    end
    else grant_line <= {grant_line[0], grant_line[1]};
  end
end
assign grant_line_ready[0] = grant_line[0] & resource_ready;
assign grant_out_priority[0] = grant_line_ready[0] & request_in[0];
assign grant_line_ready[1] = grant_line[1] & resource_ready;
assign grant_out_priority[1] = grant_line_ready[1] & request_in[1];
always_comb begin
  tmp_done = 1'h0;
  tmp_out_first = 1'h0;
  if (~tmp_done) begin
    if (request_in[0]) begin
      tmp_out_first = 1'h0;
      tmp_done = 1'h1;
    end
  end
  if (~tmp_done) begin
    if (request_in[1]) begin
      tmp_out_first = 1'h1;
      tmp_done = 1'h1;
    end
  end
end
assign grant_out_consolation[0] = resource_ready & request_in[0] & (tmp_out_first == 1'h0);
assign grant_out[0] = (|grant_out_priority) ? grant_out_priority[0]: grant_out_consolation[0];
assign grant_out_consolation[1] = resource_ready & request_in[1] & (tmp_out_first == 1'h1);
assign grant_out[1] = (|grant_out_priority) ? grant_out_priority[1]: grant_out_consolation[1];
endmodule   // arbiter_2_in_RR_algo

module arbiter_4_in_RR_algo (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [3:0] request_in,
  input logic resource_ready,
  input logic rst_n,
  output logic [3:0] grant_out
);

logic [3:0] grant_line;
logic [3:0] grant_line_ready;
logic [3:0] grant_out_consolation;
logic [3:0] grant_out_priority;
logic tmp_done;
logic [1:0] tmp_out_first;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    grant_line <= 4'h1;
  end
  else if (clk_en) begin
    if (flush) begin
      grant_line <= 4'h1;
    end
    else grant_line <= {grant_line[2:0], grant_line[3]};
  end
end
assign grant_line_ready[0] = grant_line[0] & resource_ready;
assign grant_out_priority[0] = grant_line_ready[0] & request_in[0];
assign grant_line_ready[1] = grant_line[1] & resource_ready;
assign grant_out_priority[1] = grant_line_ready[1] & request_in[1];
assign grant_line_ready[2] = grant_line[2] & resource_ready;
assign grant_out_priority[2] = grant_line_ready[2] & request_in[2];
assign grant_line_ready[3] = grant_line[3] & resource_ready;
assign grant_out_priority[3] = grant_line_ready[3] & request_in[3];
always_comb begin
  tmp_done = 1'h0;
  tmp_out_first = 2'h0;
  if (~tmp_done) begin
    if (request_in[0]) begin
      tmp_out_first = 2'h0;
      tmp_done = 1'h1;
    end
  end
  if (~tmp_done) begin
    if (request_in[1]) begin
      tmp_out_first = 2'h1;
      tmp_done = 1'h1;
    end
  end
  if (~tmp_done) begin
    if (request_in[2]) begin
      tmp_out_first = 2'h2;
      tmp_done = 1'h1;
    end
  end
  if (~tmp_done) begin
    if (request_in[3]) begin
      tmp_out_first = 2'h3;
      tmp_done = 1'h1;
    end
  end
end
assign grant_out_consolation[0] = resource_ready & request_in[0] & (tmp_out_first == 2'h0);
assign grant_out[0] = (|grant_out_priority) ? grant_out_priority[0]: grant_out_consolation[0];
assign grant_out_consolation[1] = resource_ready & request_in[1] & (tmp_out_first == 2'h1);
assign grant_out[1] = (|grant_out_priority) ? grant_out_priority[1]: grant_out_consolation[1];
assign grant_out_consolation[2] = resource_ready & request_in[2] & (tmp_out_first == 2'h2);
assign grant_out[2] = (|grant_out_priority) ? grant_out_priority[2]: grant_out_consolation[2];
assign grant_out_consolation[3] = resource_ready & request_in[3] & (tmp_out_first == 2'h3);
assign grant_out[3] = (|grant_out_priority) ? grant_out_priority[3]: grant_out_consolation[3];
endmodule   // arbiter_4_in_RR_algo

module buffet_like_16 (
  input logic [1:0] [3:0] buffet_capacity_log,
  input logic clk,
  input logic clk_en,
  input logic [3:0] [15:0] data_from_mem,
  input logic flush,
  input logic [0:0] [16:0] rd_ID,
  input logic rd_ID_valid,
  input logic [0:0] [16:0] rd_addr,
  input logic rd_addr_valid,
  input logic [0:0] [16:0] rd_op,
  input logic rd_op_valid,
  input logic rd_rsp_data_ready,
  input logic rst_n,
  input logic tile_en,
  input logic [0:0] [16:0] wr_ID,
  input logic wr_ID_valid,
  input logic [0:0] [16:0] wr_addr,
  input logic wr_addr_valid,
  input logic [0:0] [16:0] wr_data,
  input logic wr_data_valid,
  output logic [8:0] addr_to_mem,
  output logic [3:0] [15:0] data_to_mem,
  output logic rd_ID_ready,
  output logic rd_addr_ready,
  output logic rd_op_ready,
  output logic [0:0] [16:0] rd_rsp_data,
  output logic rd_rsp_data_valid,
  output logic ren_to_mem,
  output logic wen_to_mem,
  output logic wr_ID_ready,
  output logic wr_addr_ready,
  output logic wr_data_ready
);

typedef enum logic {
  RD_START_0 = 1'h0
} read_fsm_0_state;
typedef enum logic {
  RD_START_1 = 1'h0
} read_fsm_1_state;
typedef enum logic[1:0] {
  MODIFY_0 = 2'h0,
  WRITING_0 = 2'h1,
  WR_START_0 = 2'h2
} write_fsm_0_state;
typedef enum logic[1:0] {
  MODIFY_1 = 2'h0,
  WRITING_1 = 2'h1,
  WR_START_1 = 2'h2
} write_fsm_1_state;
logic PREVIOUS_WR_OP;
logic [15:0] addr_to_mem_local;
logic any_sram_lock;
logic [3:0] base_rr;
logic [1:0][15:0] blk_base;
logic [1:0][15:0] blk_bounds;
logic [0:0][31:0] blk_fifo_0_data_in;
logic [0:0][31:0] blk_fifo_0_data_out;
logic blk_fifo_0_empty;
logic blk_fifo_0_full;
logic [0:0][31:0] blk_fifo_1_data_in;
logic [0:0][31:0] blk_fifo_1_data_out;
logic blk_fifo_1_empty;
logic blk_fifo_1_full;
logic [1:0] blk_full;
logic [1:0] blk_valid;
logic [1:0][15:0] buffet_base;
logic [1:0][15:0] buffet_capacity;
logic [1:0][15:0] buffet_capacity_mask;
logic [15:0] cached_read_word_addr_0;
logic [15:0] cached_read_word_addr_1;
logic [15:0] chosen_read_0;
logic [15:0] chosen_read_1;
logic clr_cached_read_0;
logic clr_cached_read_1;
logic clr_write_wide_word_0;
logic clr_write_wide_word_1;
logic [15:0] curr_base_0;
logic [15:0] curr_base_1;
logic [15:0] curr_base_pre_0;
logic [15:0] curr_base_pre_1;
logic [15:0] curr_bounds_0;
logic [15:0] curr_bounds_1;
logic [1:0][15:0] curr_capacity_pre;
logic [15:0] decode_ret_size_request_full_blk_bounds;
logic decode_sel_done_size_request_full_blk_bounds;
logic [1:0] en_curr_base;
logic [1:0] en_curr_bounds;
logic first_base_set_0_sticky;
logic first_base_set_0_was_high;
logic first_base_set_1_sticky;
logic first_base_set_1_was_high;
logic gclk;
logic joined_in_fifo;
logic [15:0] last_read_ID;
logic [1:0] last_read_addr;
logic [15:0] last_read_addr_wide;
logic [3:0] mem_acq;
logic [2:0] num_bits_valid_mask_0_sum;
logic [2:0] num_bits_valid_mask_1_sum;
logic [1:0] pop_blk;
logic pop_in_fifos;
logic [1:0] pop_in_full;
logic [1:0] push_blk;
logic rd_ID_fifo_empty;
logic rd_ID_fifo_full;
logic [15:0] rd_ID_fifo_out_data;
logic rd_ID_fifo_pop;
logic rd_ID_fifo_valid;
logic rd_addr_fifo_empty;
logic rd_addr_fifo_full;
logic [15:0] rd_addr_fifo_out_addr;
logic rd_addr_fifo_pop;
logic rd_addr_fifo_valid;
logic rd_op_fifo_empty;
logic rd_op_fifo_full;
logic [15:0] rd_op_fifo_out_op;
logic rd_op_fifo_pop;
logic rd_op_fifo_valid;
logic rd_rsp_fifo_almost_full;
logic [0:0][16:0] rd_rsp_fifo_data_out;
logic rd_rsp_fifo_empty;
logic rd_rsp_fifo_full;
logic [16:0] rd_rsp_fifo_in_data;
logic rd_rsp_fifo_push;
logic [15:0] read_ID_d1;
logic read_d1;
logic read_from_sram_write_side_0;
logic read_from_sram_write_side_1;
read_fsm_0_state read_fsm_0_current_state;
read_fsm_0_state read_fsm_0_next_state;
read_fsm_1_state read_fsm_1_current_state;
read_fsm_1_state read_fsm_1_next_state;
logic read_joined;
logic read_pop;
logic [1:0] read_pop_full;
logic [3:0][15:0] read_wide_word_0;
logic [3:0][15:0] read_wide_word_1;
logic read_wide_word_valid_sticky_0_sticky;
logic read_wide_word_valid_sticky_0_was_high;
logic read_wide_word_valid_sticky_1_sticky;
logic read_wide_word_valid_sticky_1_was_high;
logic [1:0] ren_full;
logic ren_full_delayed_0;
logic ren_full_delayed_1;
logic rr_arbiter_resource_ready;
logic set_cached_read_0;
logic set_cached_read_1;
logic set_read_word_addr_0;
logic set_read_word_addr_1;
logic set_wide_word_addr_0;
logic set_wide_word_addr_1;
logic set_write_wide_word_0;
logic set_write_wide_word_1;
logic [1:0] size_request_full;
logic sram_lock_0;
logic sram_lock_1;
logic [15:0] tmp_addr_0;
logic [15:0] tmp_addr_1;
logic [15:0] tmp_rd_base;
logic [15:0] tmp_wr_base;
logic use_cached_read_0;
logic use_cached_read_1;
logic valid_from_mem;
logic [1:0] wen_full;
logic wr_ID_fifo_empty;
logic wr_ID_fifo_full;
logic [15:0] wr_ID_fifo_out_data;
logic wr_ID_fifo_pop;
logic wr_ID_fifo_valid;
logic wr_addr_fifo_empty;
logic wr_addr_fifo_full;
logic [15:0] wr_addr_fifo_out_data;
logic wr_addr_fifo_pop;
logic wr_addr_fifo_valid;
logic [0:0][16:0] wr_data_fifo_data_out;
logic wr_data_fifo_empty;
logic wr_data_fifo_full;
logic [15:0] wr_data_fifo_out_data;
logic wr_data_fifo_out_op;
logic wr_data_fifo_pop;
logic wr_data_fifo_valid;
write_fsm_0_state write_fsm_0_current_state;
write_fsm_0_state write_fsm_0_next_state;
write_fsm_1_state write_fsm_1_current_state;
write_fsm_1_state write_fsm_1_next_state;
logic write_full_word_0;
logic write_full_word_1;
logic write_to_sram_0;
logic write_to_sram_1;
logic [3:0][15:0] write_wide_word_comb_in_0;
logic [3:0][15:0] write_wide_word_comb_in_1;
logic [3:0][15:0] write_wide_word_comb_out_0;
logic [3:0][15:0] write_wide_word_comb_out_1;
logic [3:0] write_wide_word_mask_comb_0;
logic [3:0] write_wide_word_mask_comb_1;
logic [3:0] write_wide_word_mask_reg_in_0;
logic [3:0] write_wide_word_mask_reg_in_1;
logic [3:0] write_wide_word_mask_reg_out_0;
logic [3:0] write_wide_word_mask_reg_out_1;
logic [3:0] write_wide_word_mask_reg_strg_0;
logic [3:0] write_wide_word_mask_reg_strg_1;
logic [3:0][15:0] write_wide_word_modified_0;
logic [3:0][15:0] write_wide_word_modified_1;
logic [3:0][15:0] write_wide_word_reg_0;
logic [3:0][15:0] write_wide_word_reg_1;
logic [15:0] write_word_addr_reg_0;
logic [15:0] write_word_addr_reg_1;
logic write_word_addr_valid_sticky_0_sticky;
logic write_word_addr_valid_sticky_0_was_high;
logic write_word_addr_valid_sticky_1_sticky;
logic write_word_addr_valid_sticky_1_was_high;
assign gclk = clk & tile_en;
assign buffet_capacity_mask[0][0] = (buffet_capacity_log[0] > 4'h0) & (buffet_capacity_log[0] != 4'h0);
assign buffet_capacity_mask[0][1] = (buffet_capacity_log[0] > 4'h1) & (buffet_capacity_log[0] != 4'h0);
assign buffet_capacity_mask[0][2] = (buffet_capacity_log[0] > 4'h2) & (buffet_capacity_log[0] != 4'h0);
assign buffet_capacity_mask[0][3] = (buffet_capacity_log[0] > 4'h3) & (buffet_capacity_log[0] != 4'h0);
assign buffet_capacity_mask[0][4] = (buffet_capacity_log[0] > 4'h4) & (buffet_capacity_log[0] != 4'h0);
assign buffet_capacity_mask[0][5] = (buffet_capacity_log[0] > 4'h5) & (buffet_capacity_log[0] != 4'h0);
assign buffet_capacity_mask[0][6] = (buffet_capacity_log[0] > 4'h6) & (buffet_capacity_log[0] != 4'h0);
assign buffet_capacity_mask[0][7] = (buffet_capacity_log[0] > 4'h7) & (buffet_capacity_log[0] != 4'h0);
assign buffet_capacity_mask[0][8] = (buffet_capacity_log[0] > 4'h8) & (buffet_capacity_log[0] != 4'h0);
assign buffet_capacity_mask[0][9] = (buffet_capacity_log[0] > 4'h9) & (buffet_capacity_log[0] != 4'h0);
assign buffet_capacity_mask[0][10] = (buffet_capacity_log[0] > 4'hA) & (buffet_capacity_log[0] != 4'h0);
assign buffet_capacity_mask[0][11] = (buffet_capacity_log[0] > 4'hB) & (buffet_capacity_log[0] != 4'h0);
assign buffet_capacity_mask[0][12] = (buffet_capacity_log[0] > 4'hC) & (buffet_capacity_log[0] != 4'h0);
assign buffet_capacity_mask[0][13] = (buffet_capacity_log[0] > 4'hD) & (buffet_capacity_log[0] != 4'h0);
assign buffet_capacity_mask[0][14] = (buffet_capacity_log[0] > 4'hE) & (buffet_capacity_log[0] != 4'h0);
assign buffet_capacity_mask[0][15] = (buffet_capacity_log[0] > 4'hF) & (buffet_capacity_log[0] != 4'h0);
assign buffet_capacity_mask[1][0] = (buffet_capacity_log[1] > 4'h0) & (buffet_capacity_log[1] != 4'h0);
assign buffet_capacity_mask[1][1] = (buffet_capacity_log[1] > 4'h1) & (buffet_capacity_log[1] != 4'h0);
assign buffet_capacity_mask[1][2] = (buffet_capacity_log[1] > 4'h2) & (buffet_capacity_log[1] != 4'h0);
assign buffet_capacity_mask[1][3] = (buffet_capacity_log[1] > 4'h3) & (buffet_capacity_log[1] != 4'h0);
assign buffet_capacity_mask[1][4] = (buffet_capacity_log[1] > 4'h4) & (buffet_capacity_log[1] != 4'h0);
assign buffet_capacity_mask[1][5] = (buffet_capacity_log[1] > 4'h5) & (buffet_capacity_log[1] != 4'h0);
assign buffet_capacity_mask[1][6] = (buffet_capacity_log[1] > 4'h6) & (buffet_capacity_log[1] != 4'h0);
assign buffet_capacity_mask[1][7] = (buffet_capacity_log[1] > 4'h7) & (buffet_capacity_log[1] != 4'h0);
assign buffet_capacity_mask[1][8] = (buffet_capacity_log[1] > 4'h8) & (buffet_capacity_log[1] != 4'h0);
assign buffet_capacity_mask[1][9] = (buffet_capacity_log[1] > 4'h9) & (buffet_capacity_log[1] != 4'h0);
assign buffet_capacity_mask[1][10] = (buffet_capacity_log[1] > 4'hA) & (buffet_capacity_log[1] != 4'h0);
assign buffet_capacity_mask[1][11] = (buffet_capacity_log[1] > 4'hB) & (buffet_capacity_log[1] != 4'h0);
assign buffet_capacity_mask[1][12] = (buffet_capacity_log[1] > 4'hC) & (buffet_capacity_log[1] != 4'h0);
assign buffet_capacity_mask[1][13] = (buffet_capacity_log[1] > 4'hD) & (buffet_capacity_log[1] != 4'h0);
assign buffet_capacity_mask[1][14] = (buffet_capacity_log[1] > 4'hE) & (buffet_capacity_log[1] != 4'h0);
assign buffet_capacity_mask[1][15] = (buffet_capacity_log[1] > 4'hF) & (buffet_capacity_log[1] != 4'h0);
assign buffet_capacity[0] = (buffet_capacity_log[0] == 4'h0) ? 16'h0: 16'h1 << 16'(buffet_capacity_log[0] +
    4'h2);
assign buffet_capacity[1] = (buffet_capacity_log[1] == 4'h0) ? 16'h0: 16'h1 << 16'(buffet_capacity_log[1] +
    4'h2);
assign buffet_base[0] = 16'h0;
assign buffet_base[1] = 16'h100;
assign {wr_data_fifo_out_op, wr_data_fifo_out_data} = wr_data_fifo_data_out;
assign wr_data_ready = ~wr_data_fifo_full;
assign wr_data_fifo_valid = ~wr_data_fifo_empty;
assign wr_addr_ready = ~wr_addr_fifo_full;
assign wr_addr_fifo_valid = ~wr_addr_fifo_empty;
assign wr_ID_ready = ~wr_ID_fifo_full;
assign wr_ID_fifo_valid = ~wr_ID_fifo_empty;
assign rd_op_ready = ~rd_op_fifo_full;
assign rd_op_fifo_valid = ~rd_op_fifo_empty;
assign rd_addr_ready = ~rd_addr_fifo_full;
assign rd_addr_fifo_valid = ~rd_addr_fifo_empty;
assign rd_ID_ready = ~rd_ID_fifo_full;
assign rd_ID_fifo_valid = ~rd_ID_fifo_empty;
assign read_joined = rd_ID_fifo_valid & rd_op_fifo_valid & rd_addr_fifo_valid;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    curr_bounds_0 <= 16'hFFFF;
  end
  else if (clk_en) begin
    if (flush) begin
      curr_bounds_0 <= 16'hFFFF;
    end
    else if (1'h0) begin
      curr_bounds_0 <= 16'h0;
    end
    else if (en_curr_bounds[0]) begin
      curr_bounds_0 <= wr_addr_fifo_out_data;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    curr_bounds_1 <= 16'hFFFF;
  end
  else if (clk_en) begin
    if (flush) begin
      curr_bounds_1 <= 16'hFFFF;
    end
    else if (1'h0) begin
      curr_bounds_1 <= 16'h0;
    end
    else if (en_curr_bounds[1]) begin
      curr_bounds_1 <= wr_addr_fifo_out_data;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    first_base_set_0_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      first_base_set_0_was_high <= 1'h0;
    end
    else if (1'h0) begin
      first_base_set_0_was_high <= 1'h0;
    end
    else if (en_curr_base[0]) begin
      first_base_set_0_was_high <= 1'h1;
    end
  end
end
assign first_base_set_0_sticky = first_base_set_0_was_high;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    first_base_set_1_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      first_base_set_1_was_high <= 1'h0;
    end
    else if (1'h0) begin
      first_base_set_1_was_high <= 1'h0;
    end
    else if (en_curr_base[1]) begin
      first_base_set_1_was_high <= 1'h1;
    end
  end
end
assign first_base_set_1_sticky = first_base_set_1_was_high;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    curr_base_0 <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      curr_base_0 <= 16'h0;
    end
    else if (1'h0) begin
      curr_base_0 <= 16'h0;
    end
    else if (en_curr_base[0]) begin
      curr_base_0 <= curr_base_pre_0;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    curr_base_1 <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      curr_base_1 <= 16'h0;
    end
    else if (1'h0) begin
      curr_base_1 <= 16'h0;
    end
    else if (en_curr_base[1]) begin
      curr_base_1 <= curr_base_pre_1;
    end
  end
end
assign curr_base_pre_0 = first_base_set_0_sticky ? (curr_bounds_0 >> 16'h2) + 16'h1 + curr_base_0: 16'h0;
assign curr_base_pre_1 = first_base_set_1_sticky ? (curr_bounds_1 >> 16'h2) + 16'h1 + curr_base_1: 16'h0;
assign addr_to_mem = addr_to_mem_local[8:0];
assign tmp_addr_0 = ((16'(wr_addr_fifo_out_data[15:2]) + curr_base_0) & buffet_capacity_mask[0]) +
    buffet_base[0];
assign tmp_addr_1 = ((16'(wr_addr_fifo_out_data[15:2]) + curr_base_1) & buffet_capacity_mask[1]) +
    buffet_base[1];

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    write_word_addr_reg_0 <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      write_word_addr_reg_0 <= 16'h0;
    end
    else if (1'h0) begin
      write_word_addr_reg_0 <= 16'h0;
    end
    else if (set_wide_word_addr_0) begin
      write_word_addr_reg_0 <= tmp_addr_0;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    write_word_addr_reg_1 <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      write_word_addr_reg_1 <= 16'h0;
    end
    else if (1'h0) begin
      write_word_addr_reg_1 <= 16'h0;
    end
    else if (set_wide_word_addr_1) begin
      write_word_addr_reg_1 <= tmp_addr_1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    write_word_addr_valid_sticky_0_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      write_word_addr_valid_sticky_0_was_high <= 1'h0;
    end
    else if (1'h0) begin
      write_word_addr_valid_sticky_0_was_high <= 1'h0;
    end
    else if (set_wide_word_addr_0) begin
      write_word_addr_valid_sticky_0_was_high <= 1'h1;
    end
  end
end
assign write_word_addr_valid_sticky_0_sticky = write_word_addr_valid_sticky_0_was_high;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    write_word_addr_valid_sticky_1_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      write_word_addr_valid_sticky_1_was_high <= 1'h0;
    end
    else if (1'h0) begin
      write_word_addr_valid_sticky_1_was_high <= 1'h0;
    end
    else if (set_wide_word_addr_1) begin
      write_word_addr_valid_sticky_1_was_high <= 1'h1;
    end
  end
end
assign write_word_addr_valid_sticky_1_sticky = write_word_addr_valid_sticky_1_was_high;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    write_wide_word_mask_reg_strg_0 <= 4'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      write_wide_word_mask_reg_strg_0 <= 4'h0;
    end
    else if (1'h0) begin
      write_wide_word_mask_reg_strg_0 <= 4'h0;
    end
    else if (set_write_wide_word_0 | clr_write_wide_word_0) begin
      write_wide_word_mask_reg_strg_0 <= write_wide_word_mask_reg_in_0;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    write_wide_word_mask_reg_strg_1 <= 4'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      write_wide_word_mask_reg_strg_1 <= 4'h0;
    end
    else if (1'h0) begin
      write_wide_word_mask_reg_strg_1 <= 4'h0;
    end
    else if (set_write_wide_word_1 | clr_write_wide_word_1) begin
      write_wide_word_mask_reg_strg_1 <= write_wide_word_mask_reg_in_1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    write_wide_word_reg_0 <= 64'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      write_wide_word_reg_0 <= 64'h0;
    end
    else if (1'h0) begin
      write_wide_word_reg_0 <= 64'h0;
    end
    else if (set_write_wide_word_0 | clr_write_wide_word_0) begin
      write_wide_word_reg_0 <= write_wide_word_comb_in_0;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    write_wide_word_reg_1 <= 64'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      write_wide_word_reg_1 <= 64'h0;
    end
    else if (1'h0) begin
      write_wide_word_reg_1 <= 64'h0;
    end
    else if (set_write_wide_word_1 | clr_write_wide_word_1) begin
      write_wide_word_reg_1 <= write_wide_word_comb_in_1;
    end
  end
end
assign write_wide_word_comb_out_0[0] = write_wide_word_mask_reg_out_0[0] ? write_wide_word_reg_0[0]:
    wr_data_fifo_out_data;
assign write_wide_word_comb_out_0[1] = write_wide_word_mask_reg_out_0[1] ? write_wide_word_reg_0[1]:
    wr_data_fifo_out_data;
assign write_wide_word_comb_out_0[2] = write_wide_word_mask_reg_out_0[2] ? write_wide_word_reg_0[2]:
    wr_data_fifo_out_data;
assign write_wide_word_comb_out_0[3] = write_wide_word_mask_reg_out_0[3] ? write_wide_word_reg_0[3]:
    wr_data_fifo_out_data;
assign write_wide_word_comb_out_1[0] = write_wide_word_mask_reg_out_1[0] ? write_wide_word_reg_1[0]:
    wr_data_fifo_out_data;
assign write_wide_word_comb_out_1[1] = write_wide_word_mask_reg_out_1[1] ? write_wide_word_reg_1[1]:
    wr_data_fifo_out_data;
assign write_wide_word_comb_out_1[2] = write_wide_word_mask_reg_out_1[2] ? write_wide_word_reg_1[2]:
    wr_data_fifo_out_data;
assign write_wide_word_comb_out_1[3] = write_wide_word_mask_reg_out_1[3] ? write_wide_word_reg_1[3]:
    wr_data_fifo_out_data;
assign write_wide_word_comb_in_0[0] = (write_wide_word_mask_reg_out_0[0] & (~clr_write_wide_word_0)) ?
    write_wide_word_reg_0[0]: wr_data_fifo_out_data;
assign write_wide_word_comb_in_0[1] = (write_wide_word_mask_reg_out_0[1] & (~clr_write_wide_word_0)) ?
    write_wide_word_reg_0[1]: wr_data_fifo_out_data;
assign write_wide_word_comb_in_0[2] = (write_wide_word_mask_reg_out_0[2] & (~clr_write_wide_word_0)) ?
    write_wide_word_reg_0[2]: wr_data_fifo_out_data;
assign write_wide_word_comb_in_0[3] = (write_wide_word_mask_reg_out_0[3] & (~clr_write_wide_word_0)) ?
    write_wide_word_reg_0[3]: wr_data_fifo_out_data;
assign write_wide_word_comb_in_1[0] = (write_wide_word_mask_reg_out_1[0] & (~clr_write_wide_word_1)) ?
    write_wide_word_reg_1[0]: wr_data_fifo_out_data;
assign write_wide_word_comb_in_1[1] = (write_wide_word_mask_reg_out_1[1] & (~clr_write_wide_word_1)) ?
    write_wide_word_reg_1[1]: wr_data_fifo_out_data;
assign write_wide_word_comb_in_1[2] = (write_wide_word_mask_reg_out_1[2] & (~clr_write_wide_word_1)) ?
    write_wide_word_reg_1[2]: wr_data_fifo_out_data;
assign write_wide_word_comb_in_1[3] = (write_wide_word_mask_reg_out_1[3] & (~clr_write_wide_word_1)) ?
    write_wide_word_reg_1[3]: wr_data_fifo_out_data;
assign write_wide_word_modified_0[0] = write_wide_word_mask_reg_out_0[0] ? write_wide_word_reg_0[0]: data_from_mem[0];
assign write_wide_word_modified_0[1] = write_wide_word_mask_reg_out_0[1] ? write_wide_word_reg_0[1]: data_from_mem[1];
assign write_wide_word_modified_0[2] = write_wide_word_mask_reg_out_0[2] ? write_wide_word_reg_0[2]: data_from_mem[2];
assign write_wide_word_modified_0[3] = write_wide_word_mask_reg_out_0[3] ? write_wide_word_reg_0[3]: data_from_mem[3];
assign write_wide_word_modified_1[0] = write_wide_word_mask_reg_out_1[0] ? write_wide_word_reg_1[0]: data_from_mem[0];
assign write_wide_word_modified_1[1] = write_wide_word_mask_reg_out_1[1] ? write_wide_word_reg_1[1]: data_from_mem[1];
assign write_wide_word_modified_1[2] = write_wide_word_mask_reg_out_1[2] ? write_wide_word_reg_1[2]: data_from_mem[2];
assign write_wide_word_modified_1[3] = write_wide_word_mask_reg_out_1[3] ? write_wide_word_reg_1[3]: data_from_mem[3];
assign write_wide_word_mask_reg_out_0 = write_wide_word_mask_reg_strg_0;
assign write_wide_word_mask_reg_out_1 = write_wide_word_mask_reg_strg_1;
assign write_wide_word_mask_comb_0 = write_wide_word_mask_reg_out_0 | 4'(2'(((tmp_addr_0 == write_word_addr_reg_0) &
    joined_in_fifo & (1'h1 == wr_data_fifo_out_op) & (16'h0 == wr_ID_fifo_out_data))
    ? 1'h1: 1'h0) << wr_addr_fifo_out_data[1:0]);
assign write_wide_word_mask_comb_1 = write_wide_word_mask_reg_out_1 | 4'(2'(((tmp_addr_1 == write_word_addr_reg_1) &
    joined_in_fifo & (1'h1 == wr_data_fifo_out_op) & (16'h1 == wr_ID_fifo_out_data))
    ? 1'h1: 1'h0) << wr_addr_fifo_out_data[1:0]);
assign write_wide_word_mask_reg_in_0 = (clr_write_wide_word_0 ? 4'h0: write_wide_word_mask_reg_out_0) |
    (((((clr_write_wide_word_0 & (tmp_addr_0 != write_word_addr_reg_0)) |
    ((tmp_addr_0 == write_word_addr_reg_0) & ((~write_full_word_0) |
    (write_full_word_0 & (~mem_acq[0]))))) & (1'h1 == wr_data_fifo_out_op) & (16'h0
    == wr_ID_fifo_out_data)) ? {3'h0, joined_in_fifo}: 4'h0) <<
    4'(wr_addr_fifo_out_data[1:0]));
assign write_wide_word_mask_reg_in_1 = (clr_write_wide_word_1 ? 4'h0: write_wide_word_mask_reg_out_1) |
    (((((clr_write_wide_word_1 & (tmp_addr_1 != write_word_addr_reg_1)) |
    ((tmp_addr_1 == write_word_addr_reg_1) & ((~write_full_word_1) |
    (write_full_word_1 & (~mem_acq[2]))))) & (1'h1 == wr_data_fifo_out_op) & (16'h1
    == wr_ID_fifo_out_data)) ? {3'h0, joined_in_fifo}: 4'h0) <<
    4'(wr_addr_fifo_out_data[1:0]));
always_comb begin
  num_bits_valid_mask_0_sum = 3'h0;
  num_bits_valid_mask_0_sum = num_bits_valid_mask_0_sum + 3'(write_wide_word_mask_comb_0[0]);
  num_bits_valid_mask_0_sum = num_bits_valid_mask_0_sum + 3'(write_wide_word_mask_comb_0[1]);
  num_bits_valid_mask_0_sum = num_bits_valid_mask_0_sum + 3'(write_wide_word_mask_comb_0[2]);
  num_bits_valid_mask_0_sum = num_bits_valid_mask_0_sum + 3'(write_wide_word_mask_comb_0[3]);
end
always_comb begin
  num_bits_valid_mask_1_sum = 3'h0;
  num_bits_valid_mask_1_sum = num_bits_valid_mask_1_sum + 3'(write_wide_word_mask_comb_1[0]);
  num_bits_valid_mask_1_sum = num_bits_valid_mask_1_sum + 3'(write_wide_word_mask_comb_1[1]);
  num_bits_valid_mask_1_sum = num_bits_valid_mask_1_sum + 3'(write_wide_word_mask_comb_1[2]);
  num_bits_valid_mask_1_sum = num_bits_valid_mask_1_sum + 3'(write_wide_word_mask_comb_1[3]);
end
assign write_full_word_0 = 3'h4 == num_bits_valid_mask_0_sum;
assign write_full_word_1 = 3'h4 == num_bits_valid_mask_1_sum;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    read_wide_word_0 <= 64'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      read_wide_word_0 <= 64'h0;
    end
    else if (1'h0) begin
      read_wide_word_0 <= 64'h0;
    end
    else if (set_cached_read_0) begin
      read_wide_word_0 <= data_from_mem;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    read_wide_word_1 <= 64'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      read_wide_word_1 <= 64'h0;
    end
    else if (1'h0) begin
      read_wide_word_1 <= 64'h0;
    end
    else if (set_cached_read_1) begin
      read_wide_word_1 <= data_from_mem;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    read_wide_word_valid_sticky_0_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      read_wide_word_valid_sticky_0_was_high <= 1'h0;
    end
    else if (clr_cached_read_0) begin
      read_wide_word_valid_sticky_0_was_high <= 1'h0;
    end
    else if (set_cached_read_0) begin
      read_wide_word_valid_sticky_0_was_high <= 1'h1;
    end
  end
end
assign read_wide_word_valid_sticky_0_sticky = set_cached_read_0 | read_wide_word_valid_sticky_0_was_high;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    read_wide_word_valid_sticky_1_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      read_wide_word_valid_sticky_1_was_high <= 1'h0;
    end
    else if (clr_cached_read_1) begin
      read_wide_word_valid_sticky_1_was_high <= 1'h0;
    end
    else if (set_cached_read_1) begin
      read_wide_word_valid_sticky_1_was_high <= 1'h1;
    end
  end
end
assign read_wide_word_valid_sticky_1_sticky = set_cached_read_1 | read_wide_word_valid_sticky_1_was_high;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    last_read_addr <= 2'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      last_read_addr <= 2'h0;
    end
    else if (1'h0) begin
      last_read_addr <= 2'h0;
    end
    else if (ren_to_mem) begin
      last_read_addr <= rd_addr_fifo_out_addr[1:0];
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    last_read_addr_wide <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      last_read_addr_wide <= 16'h0;
    end
    else if (1'h0) begin
      last_read_addr_wide <= 16'h0;
    end
    else if (ren_to_mem) begin
      last_read_addr_wide <= addr_to_mem_local;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    last_read_ID <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      last_read_ID <= 16'h0;
    end
    else if (1'h0) begin
      last_read_ID <= 16'h0;
    end
    else if (ren_to_mem) begin
      last_read_ID <= rd_ID_fifo_out_data;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    cached_read_word_addr_0 <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      cached_read_word_addr_0 <= 16'h0;
    end
    else if (1'h0) begin
      cached_read_word_addr_0 <= 16'h0;
    end
    else if (set_read_word_addr_0) begin
      cached_read_word_addr_0 <= addr_to_mem_local;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    cached_read_word_addr_1 <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      cached_read_word_addr_1 <= 16'h0;
    end
    else if (1'h0) begin
      cached_read_word_addr_1 <= 16'h0;
    end
    else if (set_read_word_addr_1) begin
      cached_read_word_addr_1 <= addr_to_mem_local;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    ren_full_delayed_0 <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      ren_full_delayed_0 <= 1'h0;
    end
    else if (1'h0) begin
      ren_full_delayed_0 <= 1'h0;
    end
    else if (1'h1) begin
      ren_full_delayed_0 <= ren_full[0];
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    ren_full_delayed_1 <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      ren_full_delayed_1 <= 1'h0;
    end
    else if (1'h0) begin
      ren_full_delayed_1 <= 1'h0;
    end
    else if (1'h1) begin
      ren_full_delayed_1 <= ren_full[1];
    end
  end
end
assign use_cached_read_0 = read_wide_word_valid_sticky_0_sticky & ((valid_from_mem & ren_full_delayed_0) ?
    (16'h0 == last_read_ID) & (last_read_addr_wide == cached_read_word_addr_0):
    (16'h0 == rd_ID_fifo_out_data) & ((((16'(rd_addr_fifo_out_addr[15:2]) +
    blk_base[0]) & buffet_capacity_mask[0]) + buffet_base[0]) ==
    cached_read_word_addr_0) & (16'h1 == rd_op_fifo_out_op) & (~valid_from_mem) &
    read_joined);
assign use_cached_read_1 = read_wide_word_valid_sticky_1_sticky & ((valid_from_mem & ren_full_delayed_1) ?
    (16'h1 == last_read_ID) & (last_read_addr_wide == cached_read_word_addr_1):
    (16'h1 == rd_ID_fifo_out_data) & ((((16'(rd_addr_fifo_out_addr[15:2]) +
    blk_base[1]) & buffet_capacity_mask[1]) + buffet_base[1]) ==
    cached_read_word_addr_1) & (16'h1 == rd_op_fifo_out_op) & (~valid_from_mem) &
    read_joined);
assign chosen_read_0 = (use_cached_read_0 & read_wide_word_valid_sticky_0_sticky & (~valid_from_mem)) ?
    read_wide_word_0[rd_addr_fifo_out_addr[1:0]]: data_from_mem[last_read_addr[1:0]];
assign chosen_read_1 = (use_cached_read_1 & read_wide_word_valid_sticky_1_sticky & (~valid_from_mem)) ?
    read_wide_word_1[rd_addr_fifo_out_addr[1:0]]: data_from_mem[last_read_addr[1:0]];
assign any_sram_lock = |{sram_lock_0, sram_lock_1};

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    read_d1 <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      read_d1 <= 1'h0;
    end
    else if (1'h0) begin
      read_d1 <= 1'h0;
    end
    else if (1'h1) begin
      read_d1 <= |{mem_acq[1], mem_acq[3]};
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    read_ID_d1 <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      read_ID_d1 <= 16'h0;
    end
    else if (1'h0) begin
      read_ID_d1 <= 16'h0;
    end
    else if (ren_to_mem) begin
      read_ID_d1 <= rd_ID_fifo_out_data;
    end
  end
end
assign valid_from_mem = read_d1;
assign rd_rsp_data[0] = rd_rsp_fifo_data_out;
assign rd_rsp_data_valid = ~rd_rsp_fifo_empty;
always_comb begin
  decode_sel_done_size_request_full_blk_bounds = 1'h0;
  decode_ret_size_request_full_blk_bounds = 16'h0;
  if ((~decode_sel_done_size_request_full_blk_bounds) & size_request_full[0]) begin
    decode_ret_size_request_full_blk_bounds = blk_bounds[0];
    decode_sel_done_size_request_full_blk_bounds = 1'h1;
  end
  if ((~decode_sel_done_size_request_full_blk_bounds) & size_request_full[1]) begin
    decode_ret_size_request_full_blk_bounds = blk_bounds[1];
    decode_sel_done_size_request_full_blk_bounds = 1'h1;
  end
end
assign rd_rsp_fifo_in_data[15:0] = (use_cached_read_0 & read_wide_word_valid_sticky_0_sticky) ? chosen_read_0:
    (use_cached_read_1 & read_wide_word_valid_sticky_1_sticky) ? chosen_read_1:
    decode_ret_size_request_full_blk_bounds + 16'h1;
assign rd_rsp_fifo_in_data[16] = use_cached_read_0 ? 1'h0: 1'h1;
assign rd_rsp_fifo_push = valid_from_mem | (|{use_cached_read_0, use_cached_read_1}) |
    (|size_request_full);
assign joined_in_fifo = wr_data_fifo_valid & wr_addr_fifo_valid & wr_ID_fifo_valid;
assign {wr_addr_fifo_pop, wr_data_fifo_pop, wr_ID_fifo_pop} = {pop_in_fifos, pop_in_fifos, pop_in_fifos};
assign pop_in_fifos = |pop_in_full;
assign {rd_ID_fifo_pop, rd_op_fifo_pop, rd_addr_fifo_pop} = {read_pop, read_pop, read_pop};
assign read_pop = |read_pop_full;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    curr_capacity_pre[0] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      curr_capacity_pre[0] <= 16'h0;
    end
    else if (push_blk[0] || pop_blk[0]) begin
      curr_capacity_pre[0] <= (curr_capacity_pre[0] + (push_blk[0] ? blk_bounds[0]: 16'h0)) - (pop_blk[0] ?
          blk_bounds[0]: 16'h0);
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    curr_capacity_pre[1] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      curr_capacity_pre[1] <= 16'h0;
    end
    else if (push_blk[1] || pop_blk[1]) begin
      curr_capacity_pre[1] <= (curr_capacity_pre[1] + (push_blk[1] ? blk_bounds[1]: 16'h0)) - (pop_blk[1] ?
          blk_bounds[1]: 16'h0);
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    PREVIOUS_WR_OP <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      PREVIOUS_WR_OP <= 1'h0;
    end
    else if (1'h0) begin
      PREVIOUS_WR_OP <= 1'h0;
    end
    else if (1'h1) begin
      PREVIOUS_WR_OP <= wr_data_fifo_out_op;
    end
  end
end
assign blk_fifo_0_data_in = {curr_base_0, curr_bounds_0};
assign {blk_base[0], blk_bounds[0]} = blk_fifo_0_data_out;
assign blk_full[0] = blk_fifo_0_full;
assign blk_valid[0] = ~blk_fifo_0_empty;
assign blk_fifo_1_data_in = {curr_base_1, curr_bounds_1};
assign {blk_base[1], blk_bounds[1]} = blk_fifo_1_data_out;
assign blk_full[1] = blk_fifo_1_full;
assign blk_valid[1] = ~blk_fifo_1_empty;

always_ff @(posedge clk, negedge rst_n) begin
  if (!rst_n) begin
    read_fsm_0_current_state <= RD_START_0;
  end
  else if (clk_en) begin
    if (flush) begin
      read_fsm_0_current_state <= RD_START_0;
    end
    else read_fsm_0_current_state <= read_fsm_0_next_state;
  end
end
always_comb begin
  read_fsm_0_next_state = read_fsm_0_current_state;
  unique case (read_fsm_0_current_state)
    RD_START_0: read_fsm_0_next_state = RD_START_0;
    default: begin end
  endcase
end
always_comb begin
  unique case (read_fsm_0_current_state)
    RD_START_0: begin :read_fsm_0_RD_START_0_Output
        pop_blk[0] = (rd_op_fifo_out_op == 16'h0) & read_joined & (16'h0 == rd_ID_fifo_out_data);
        ren_full[0] = (rd_op_fifo_out_op == 16'h1) & (~use_cached_read_0) & read_joined &
            (~rd_rsp_fifo_almost_full) & blk_valid[0] & (((16'(rd_addr_fifo_out_addr[15:2])
            + blk_base[0] + buffet_base[0]) != cached_read_word_addr_0) |
            (~read_wide_word_valid_sticky_0_sticky)) & (16'h0 == rd_ID_fifo_out_data);
        read_pop_full[0] = ((rd_op_fifo_out_op == 16'h2) ? (~valid_from_mem) & blk_valid[0]:
            (rd_op_fifo_out_op == 16'h1) ? (mem_acq[1] | (use_cached_read_0 &
            (~valid_from_mem))) & (~rd_rsp_fifo_full): 1'h1) & read_joined & (16'h0 ==
            rd_ID_fifo_out_data);
        size_request_full[0] = blk_valid[0] & (rd_op_fifo_out_op == 16'h2) & read_joined & (16'h0 ==
            rd_ID_fifo_out_data);
        set_cached_read_0 = valid_from_mem & (16'h0 == read_ID_d1);
        clr_cached_read_0 = (rd_op_fifo_out_op == 16'h0) & read_joined & (16'h0 == rd_ID_fifo_out_data);
        set_read_word_addr_0 = ren_full[0] & mem_acq[1] & (addr_to_mem_local != cached_read_word_addr_0) &
            (16'h0 == rd_ID_fifo_out_data);
      end :read_fsm_0_RD_START_0_Output
    default: begin end
  endcase
end

always_ff @(posedge clk, negedge rst_n) begin
  if (!rst_n) begin
    read_fsm_1_current_state <= RD_START_1;
  end
  else if (clk_en) begin
    if (flush) begin
      read_fsm_1_current_state <= RD_START_1;
    end
    else read_fsm_1_current_state <= read_fsm_1_next_state;
  end
end
always_comb begin
  read_fsm_1_next_state = read_fsm_1_current_state;
  unique case (read_fsm_1_current_state)
    RD_START_1: read_fsm_1_next_state = RD_START_1;
    default: begin end
  endcase
end
always_comb begin
  unique case (read_fsm_1_current_state)
    RD_START_1: begin :read_fsm_1_RD_START_1_Output
        pop_blk[1] = (rd_op_fifo_out_op == 16'h0) & read_joined & (16'h1 == rd_ID_fifo_out_data);
        ren_full[1] = (rd_op_fifo_out_op == 16'h1) & (~use_cached_read_1) & read_joined &
            (~rd_rsp_fifo_almost_full) & blk_valid[1] & (((16'(rd_addr_fifo_out_addr[15:2])
            + blk_base[1] + buffet_base[1]) != cached_read_word_addr_1) |
            (~read_wide_word_valid_sticky_1_sticky)) & (16'h1 == rd_ID_fifo_out_data);
        read_pop_full[1] = ((rd_op_fifo_out_op == 16'h2) ? (~valid_from_mem) & blk_valid[1]:
            (rd_op_fifo_out_op == 16'h1) ? (mem_acq[3] | (use_cached_read_1 &
            (~valid_from_mem))) & (~rd_rsp_fifo_full): 1'h1) & read_joined & (16'h1 ==
            rd_ID_fifo_out_data);
        size_request_full[1] = blk_valid[1] & (rd_op_fifo_out_op == 16'h2) & read_joined & (16'h1 ==
            rd_ID_fifo_out_data);
        set_cached_read_1 = valid_from_mem & (16'h1 == read_ID_d1);
        clr_cached_read_1 = (rd_op_fifo_out_op == 16'h0) & read_joined & (16'h1 == rd_ID_fifo_out_data);
        set_read_word_addr_1 = ren_full[1] & mem_acq[3] & (addr_to_mem_local != cached_read_word_addr_1) &
            (16'h1 == rd_ID_fifo_out_data);
      end :read_fsm_1_RD_START_1_Output
    default: begin end
  endcase
end

always_ff @(posedge clk, negedge rst_n) begin
  if (!rst_n) begin
    write_fsm_0_current_state <= WR_START_0;
  end
  else if (clk_en) begin
    if (flush) begin
      write_fsm_0_current_state <= WR_START_0;
    end
    else write_fsm_0_current_state <= write_fsm_0_next_state;
  end
end
always_comb begin
  write_fsm_0_next_state = write_fsm_0_current_state;
  unique case (write_fsm_0_current_state)
    MODIFY_0: begin
        if (1'h1 == PREVIOUS_WR_OP) begin
          write_fsm_0_next_state = WRITING_0;
        end
        else if ((1'h0 == PREVIOUS_WR_OP) & (~blk_full[0])) begin
          write_fsm_0_next_state = WR_START_0;
        end
        else write_fsm_0_next_state = MODIFY_0;
      end
    WRITING_0: begin
        if (joined_in_fifo & (wr_data_fifo_out_op == 1'h0) & (~blk_full[0]) & ((write_full_word_0 & mem_acq[0]) | (num_bits_valid_mask_0_sum == 3'h0)) & (16'h0 == wr_ID_fifo_out_data)) begin
          write_fsm_0_next_state = WR_START_0;
        end
        else if (joined_in_fifo & (16'h0 == wr_ID_fifo_out_data) & mem_acq[0] & ((1'h0 == wr_data_fifo_out_op) | ((tmp_addr_0 != write_word_addr_reg_0) & write_word_addr_valid_sticky_0_sticky & (1'h1 == wr_data_fifo_out_op))) & (num_bits_valid_mask_0_sum > 3'h0) & (~write_full_word_0)) begin
          write_fsm_0_next_state = MODIFY_0;
        end
        else write_fsm_0_next_state = WRITING_0;
      end
    WR_START_0: begin
        if (joined_in_fifo & (wr_data_fifo_out_op == 1'h0) & (16'h0 == wr_ID_fifo_out_data) & tile_en) begin
          write_fsm_0_next_state = WRITING_0;
        end
        else write_fsm_0_next_state = WR_START_0;
      end
    default: write_fsm_0_next_state = write_fsm_0_current_state;
  endcase
end
always_comb begin
  unique case (write_fsm_0_current_state)
    MODIFY_0: begin :write_fsm_0_MODIFY_0_Output
        push_blk[0] = (1'h0 == PREVIOUS_WR_OP) & (~blk_full[0]);
        en_curr_base[0] = (1'h0 == PREVIOUS_WR_OP) & (~blk_full[0]);
        en_curr_bounds[0] = 1'h0;
        wen_full[0] = ~blk_full[0];
        pop_in_full[0] = ~blk_full[0];
        set_write_wide_word_0 = 1'h0;
        clr_write_wide_word_0 = ~blk_full[0];
        write_to_sram_0 = ~blk_full[0];
        read_from_sram_write_side_0 = 1'h0;
        set_wide_word_addr_0 = 1'h0;
        sram_lock_0 = ~blk_full[0];
      end :write_fsm_0_MODIFY_0_Output
    WRITING_0: begin :write_fsm_0_WRITING_0_Output
        push_blk[0] = joined_in_fifo & (wr_data_fifo_out_op == 1'h0) & (~blk_full[0]) &
            ((write_full_word_0 & mem_acq[0]) | (num_bits_valid_mask_0_sum == 3'h0)) &
            (16'h0 == wr_ID_fifo_out_data);
        en_curr_base[0] = joined_in_fifo & (wr_data_fifo_out_op == 1'h0) & (~blk_full[0]) &
            ((write_full_word_0 & mem_acq[0]) | (num_bits_valid_mask_0_sum == 3'h0)) &
            (16'h0 == wr_ID_fifo_out_data);
        set_write_wide_word_0 = (tmp_addr_0 == write_word_addr_reg_0) & write_word_addr_valid_sticky_0_sticky &
            joined_in_fifo & (wr_data_fifo_out_op == 1'h1) & (16'h0 == wr_ID_fifo_out_data);
        en_curr_bounds[0] = (mem_acq[0] | set_write_wide_word_0) & joined_in_fifo & (wr_data_fifo_out_op ==
            1'h1) & (16'h0 == wr_ID_fifo_out_data);
        wen_full[0] = joined_in_fifo & (wr_data_fifo_out_op == 1'h1) & ((buffet_capacity[0] -
            curr_capacity_pre[0]) > wr_addr_fifo_out_data) & (16'h0 == wr_ID_fifo_out_data);
        clr_write_wide_word_0 = ((tmp_addr_0 != write_word_addr_reg_0) |
            (~write_word_addr_valid_sticky_0_sticky) | ((tmp_addr_0 ==
            write_word_addr_reg_0) & write_word_addr_valid_sticky_0_sticky &
            write_full_word_0)) & joined_in_fifo & (wr_data_fifo_out_op == 1'h1) &
            mem_acq[0] & (16'h0 == wr_ID_fifo_out_data);
        write_to_sram_0 = write_full_word_0 & joined_in_fifo & ((buffet_capacity[0] -
            curr_capacity_pre[0]) > wr_addr_fifo_out_data) & (16'h0 == wr_ID_fifo_out_data);
        set_wide_word_addr_0 = ((tmp_addr_0 != write_word_addr_reg_0) |
            (~write_word_addr_valid_sticky_0_sticky)) & joined_in_fifo &
            (wr_data_fifo_out_op == 1'h1) & (16'h0 == wr_ID_fifo_out_data);
        sram_lock_0 = 1'h0;
        read_from_sram_write_side_0 = joined_in_fifo & (16'h0 == wr_ID_fifo_out_data) & (~any_sram_lock) &
            ((buffet_capacity[0] - curr_capacity_pre[0]) > wr_addr_fifo_out_data) & ((1'h0
            == wr_data_fifo_out_op) | ((tmp_addr_0 != write_word_addr_reg_0) &
            write_word_addr_valid_sticky_0_sticky & (1'h1 == wr_data_fifo_out_op))) &
            (num_bits_valid_mask_0_sum > 3'h0) & (~write_full_word_0);
        pop_in_full[0] = ((mem_acq[0] | set_write_wide_word_0) & joined_in_fifo & (wr_data_fifo_out_op ==
            1'h1) & ((buffet_capacity[0] - curr_capacity_pre[0]) > wr_addr_fifo_out_data) &
            (16'h0 == wr_ID_fifo_out_data)) | (joined_in_fifo & (wr_data_fifo_out_op ==
            1'h0) & (~blk_full[0]) & ((write_full_word_0 & mem_acq[0]) |
            (num_bits_valid_mask_0_sum == 3'h0)) & (16'h0 == wr_ID_fifo_out_data));
      end :write_fsm_0_WRITING_0_Output
    WR_START_0: begin :write_fsm_0_WR_START_0_Output
        push_blk[0] = 1'h0;
        en_curr_base[0] = 1'h0;
        en_curr_bounds[0] = 1'h0;
        wen_full[0] = 1'h0;
        pop_in_full[0] = (wr_data_fifo_out_op == 1'h0) & (16'h0 == wr_ID_fifo_out_data);
        set_write_wide_word_0 = 1'h0;
        clr_write_wide_word_0 = 1'h0;
        write_to_sram_0 = 1'h0;
        set_wide_word_addr_0 = 1'h0;
        sram_lock_0 = 1'h0;
        read_from_sram_write_side_0 = 1'h0;
      end :write_fsm_0_WR_START_0_Output
    default: begin :write_fsm_0_default_Output
        push_blk[0] = 1'h0;
        en_curr_base[0] = 1'h0;
        en_curr_bounds[0] = 1'h0;
        wen_full[0] = 1'h0;
        pop_in_full[0] = (wr_data_fifo_out_op == 1'h0) & (16'h0 == wr_ID_fifo_out_data);
        set_write_wide_word_0 = 1'h0;
        clr_write_wide_word_0 = 1'h0;
        write_to_sram_0 = 1'h0;
        set_wide_word_addr_0 = 1'h0;
        sram_lock_0 = 1'h0;
        read_from_sram_write_side_0 = 1'h0;
      end :write_fsm_0_default_Output
  endcase
end

always_ff @(posedge clk, negedge rst_n) begin
  if (!rst_n) begin
    write_fsm_1_current_state <= WR_START_1;
  end
  else if (clk_en) begin
    if (flush) begin
      write_fsm_1_current_state <= WR_START_1;
    end
    else write_fsm_1_current_state <= write_fsm_1_next_state;
  end
end
always_comb begin
  write_fsm_1_next_state = write_fsm_1_current_state;
  unique case (write_fsm_1_current_state)
    MODIFY_1: begin
        if (1'h1 == PREVIOUS_WR_OP) begin
          write_fsm_1_next_state = WRITING_1;
        end
        else if ((1'h0 == PREVIOUS_WR_OP) & (~blk_full[1])) begin
          write_fsm_1_next_state = WR_START_1;
        end
        else write_fsm_1_next_state = MODIFY_1;
      end
    WRITING_1: begin
        if (joined_in_fifo & (wr_data_fifo_out_op == 1'h0) & (~blk_full[1]) & ((write_full_word_1 & mem_acq[2]) | (num_bits_valid_mask_1_sum == 3'h0)) & (16'h1 == wr_ID_fifo_out_data)) begin
          write_fsm_1_next_state = WR_START_1;
        end
        else if (joined_in_fifo & (16'h1 == wr_ID_fifo_out_data) & mem_acq[2] & ((1'h0 == wr_data_fifo_out_op) | ((tmp_addr_1 != write_word_addr_reg_1) & write_word_addr_valid_sticky_1_sticky & (1'h1 == wr_data_fifo_out_op))) & (num_bits_valid_mask_1_sum > 3'h0) & (~write_full_word_1)) begin
          write_fsm_1_next_state = MODIFY_1;
        end
        else write_fsm_1_next_state = WRITING_1;
      end
    WR_START_1: begin
        if (joined_in_fifo & (wr_data_fifo_out_op == 1'h0) & (16'h1 == wr_ID_fifo_out_data) & tile_en) begin
          write_fsm_1_next_state = WRITING_1;
        end
        else write_fsm_1_next_state = WR_START_1;
      end
    default: write_fsm_1_next_state = write_fsm_1_current_state;
  endcase
end
always_comb begin
  unique case (write_fsm_1_current_state)
    MODIFY_1: begin :write_fsm_1_MODIFY_1_Output
        push_blk[1] = (1'h0 == PREVIOUS_WR_OP) & (~blk_full[1]);
        en_curr_base[1] = (1'h0 == PREVIOUS_WR_OP) & (~blk_full[1]);
        en_curr_bounds[1] = 1'h0;
        wen_full[1] = ~blk_full[1];
        pop_in_full[1] = ~blk_full[1];
        set_write_wide_word_1 = 1'h0;
        clr_write_wide_word_1 = ~blk_full[1];
        write_to_sram_1 = ~blk_full[1];
        read_from_sram_write_side_1 = 1'h0;
        set_wide_word_addr_1 = 1'h0;
        sram_lock_1 = ~blk_full[1];
      end :write_fsm_1_MODIFY_1_Output
    WRITING_1: begin :write_fsm_1_WRITING_1_Output
        push_blk[1] = joined_in_fifo & (wr_data_fifo_out_op == 1'h0) & (~blk_full[1]) &
            ((write_full_word_1 & mem_acq[2]) | (num_bits_valid_mask_1_sum == 3'h0)) &
            (16'h1 == wr_ID_fifo_out_data);
        en_curr_base[1] = joined_in_fifo & (wr_data_fifo_out_op == 1'h0) & (~blk_full[1]) &
            ((write_full_word_1 & mem_acq[2]) | (num_bits_valid_mask_1_sum == 3'h0)) &
            (16'h1 == wr_ID_fifo_out_data);
        set_write_wide_word_1 = (tmp_addr_1 == write_word_addr_reg_1) & write_word_addr_valid_sticky_1_sticky &
            joined_in_fifo & (wr_data_fifo_out_op == 1'h1) & (16'h1 == wr_ID_fifo_out_data);
        en_curr_bounds[1] = (mem_acq[2] | set_write_wide_word_1) & joined_in_fifo & (wr_data_fifo_out_op ==
            1'h1) & (16'h1 == wr_ID_fifo_out_data);
        wen_full[1] = joined_in_fifo & (wr_data_fifo_out_op == 1'h1) & ((buffet_capacity[1] -
            curr_capacity_pre[1]) > wr_addr_fifo_out_data) & (16'h1 == wr_ID_fifo_out_data);
        clr_write_wide_word_1 = ((tmp_addr_1 != write_word_addr_reg_1) |
            (~write_word_addr_valid_sticky_1_sticky) | ((tmp_addr_1 ==
            write_word_addr_reg_1) & write_word_addr_valid_sticky_1_sticky &
            write_full_word_1)) & joined_in_fifo & (wr_data_fifo_out_op == 1'h1) &
            mem_acq[2] & (16'h1 == wr_ID_fifo_out_data);
        write_to_sram_1 = write_full_word_1 & joined_in_fifo & ((buffet_capacity[1] -
            curr_capacity_pre[1]) > wr_addr_fifo_out_data) & (16'h1 == wr_ID_fifo_out_data);
        set_wide_word_addr_1 = ((tmp_addr_1 != write_word_addr_reg_1) |
            (~write_word_addr_valid_sticky_1_sticky)) & joined_in_fifo &
            (wr_data_fifo_out_op == 1'h1) & (16'h1 == wr_ID_fifo_out_data);
        sram_lock_1 = 1'h0;
        read_from_sram_write_side_1 = joined_in_fifo & (16'h1 == wr_ID_fifo_out_data) & (~any_sram_lock) &
            ((buffet_capacity[1] - curr_capacity_pre[1]) > wr_addr_fifo_out_data) & ((1'h0
            == wr_data_fifo_out_op) | ((tmp_addr_1 != write_word_addr_reg_1) &
            write_word_addr_valid_sticky_1_sticky & (1'h1 == wr_data_fifo_out_op))) &
            (num_bits_valid_mask_1_sum > 3'h0) & (~write_full_word_1);
        pop_in_full[1] = ((mem_acq[2] | set_write_wide_word_1) & joined_in_fifo & (wr_data_fifo_out_op ==
            1'h1) & ((buffet_capacity[1] - curr_capacity_pre[1]) > wr_addr_fifo_out_data) &
            (16'h1 == wr_ID_fifo_out_data)) | (joined_in_fifo & (wr_data_fifo_out_op ==
            1'h0) & (~blk_full[1]) & ((write_full_word_1 & mem_acq[2]) |
            (num_bits_valid_mask_1_sum == 3'h0)) & (16'h1 == wr_ID_fifo_out_data));
      end :write_fsm_1_WRITING_1_Output
    WR_START_1: begin :write_fsm_1_WR_START_1_Output
        push_blk[1] = 1'h0;
        en_curr_base[1] = 1'h0;
        en_curr_bounds[1] = 1'h0;
        wen_full[1] = 1'h0;
        pop_in_full[1] = (wr_data_fifo_out_op == 1'h0) & (16'h1 == wr_ID_fifo_out_data);
        set_write_wide_word_1 = 1'h0;
        clr_write_wide_word_1 = 1'h0;
        write_to_sram_1 = 1'h0;
        set_wide_word_addr_1 = 1'h0;
        sram_lock_1 = 1'h0;
        read_from_sram_write_side_1 = 1'h0;
      end :write_fsm_1_WR_START_1_Output
    default: begin :write_fsm_1_default_Output
        push_blk[1] = 1'h0;
        en_curr_base[1] = 1'h0;
        en_curr_bounds[1] = 1'h0;
        wen_full[1] = 1'h0;
        pop_in_full[1] = (wr_data_fifo_out_op == 1'h0) & (16'h1 == wr_ID_fifo_out_data);
        set_write_wide_word_1 = 1'h0;
        clr_write_wide_word_1 = 1'h0;
        write_to_sram_1 = 1'h0;
        set_wide_word_addr_1 = 1'h0;
        sram_lock_1 = 1'h0;
        read_from_sram_write_side_1 = 1'h0;
      end :write_fsm_1_default_Output
  endcase
end
assign base_rr = {ren_full[1], write_to_sram_1 | read_from_sram_write_side_1, {ren_full[0],
    write_to_sram_0 | read_from_sram_write_side_0}};
assign rr_arbiter_resource_ready = ~any_sram_lock;
assign ren_to_mem = (|{mem_acq[1] & ren_full[0], mem_acq[3] & ren_full[1]}) |
    (|{read_from_sram_write_side_0, read_from_sram_write_side_1});
assign wen_to_mem = |({mem_acq[0] & write_to_sram_0, mem_acq[2] & write_to_sram_1} | {sram_lock_0,
    sram_lock_1});
assign tmp_wr_base = (mem_acq[2] & write_to_sram_1) ? curr_base_1 + buffet_base[1]: (mem_acq[0] &
    write_to_sram_0) ? curr_base_0 + buffet_base[0]: 16'h0;
assign tmp_rd_base = (mem_acq[3] & ren_full[1]) ? blk_base[1] + buffet_base[1]: (mem_acq[1] &
    ren_full[0]) ? blk_base[0] + buffet_base[0]: 16'h0;
assign data_to_mem = (mem_acq[0] & write_to_sram_0) ? write_wide_word_comb_out_0: (mem_acq[2] &
    write_to_sram_1) ? write_wide_word_comb_out_1: sram_lock_0 ?
    write_wide_word_modified_0: sram_lock_1 ? write_wide_word_modified_1: 64'h0;
assign addr_to_mem_local = (wen_to_mem | mem_acq[0] | mem_acq[2]) ? (mem_acq[0] | sram_lock_0) ?
    write_word_addr_reg_0: write_word_addr_reg_1: (mem_acq[1] & ren_full[0]) ?
    ((16'(rd_addr_fifo_out_addr[15:2]) + blk_base[0]) & buffet_capacity_mask[0]) +
    buffet_base[0]: ((16'(rd_addr_fifo_out_addr[15:2]) + blk_base[1]) &
    buffet_capacity_mask[1]) + buffet_base[1];
reg_fifo_depth_2_w_17_afd_2 wr_data_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(wr_data),
  .flush(flush),
  .pop(wr_data_fifo_pop),
  .push(wr_data_valid),
  .rst_n(rst_n),
  .data_out(wr_data_fifo_data_out),
  .empty(wr_data_fifo_empty),
  .full(wr_data_fifo_full)
);

reg_fifo_depth_2_w_16_afd_2 wr_addr_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(wr_addr[0][15:0]),
  .flush(flush),
  .pop(wr_addr_fifo_pop),
  .push(wr_addr_valid),
  .rst_n(rst_n),
  .data_out(wr_addr_fifo_out_data),
  .empty(wr_addr_fifo_empty),
  .full(wr_addr_fifo_full)
);

reg_fifo_depth_2_w_16_afd_2 wr_ID_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(wr_ID[0][15:0]),
  .flush(flush),
  .pop(wr_ID_fifo_pop),
  .push(wr_ID_valid),
  .rst_n(rst_n),
  .data_out(wr_ID_fifo_out_data),
  .empty(wr_ID_fifo_empty),
  .full(wr_ID_fifo_full)
);

reg_fifo_depth_2_w_16_afd_2 rd_op_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(rd_op[0][15:0]),
  .flush(flush),
  .pop(rd_op_fifo_pop),
  .push(rd_op_valid),
  .rst_n(rst_n),
  .data_out(rd_op_fifo_out_op),
  .empty(rd_op_fifo_empty),
  .full(rd_op_fifo_full)
);

reg_fifo_depth_2_w_16_afd_2 rd_addr_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(rd_addr[0][15:0]),
  .flush(flush),
  .pop(rd_addr_fifo_pop),
  .push(rd_addr_valid),
  .rst_n(rst_n),
  .data_out(rd_addr_fifo_out_addr),
  .empty(rd_addr_fifo_empty),
  .full(rd_addr_fifo_full)
);

reg_fifo_depth_2_w_16_afd_2 rd_ID_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(rd_ID[0][15:0]),
  .flush(flush),
  .pop(rd_ID_fifo_pop),
  .push(rd_ID_valid),
  .rst_n(rst_n),
  .data_out(rd_ID_fifo_out_data),
  .empty(rd_ID_fifo_empty),
  .full(rd_ID_fifo_full)
);

reg_fifo_depth_2_w_17_afd_1 rd_rsp_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(rd_rsp_fifo_in_data),
  .flush(flush),
  .pop(rd_rsp_data_ready),
  .push(rd_rsp_fifo_push),
  .rst_n(rst_n),
  .almost_full(rd_rsp_fifo_almost_full),
  .data_out(rd_rsp_fifo_data_out),
  .empty(rd_rsp_fifo_empty),
  .full(rd_rsp_fifo_full)
);

reg_fifo_depth_2_w_32_afd_2 blk_fifo_0 (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(blk_fifo_0_data_in),
  .flush(flush),
  .pop(pop_blk[0]),
  .push(push_blk[0]),
  .rst_n(rst_n),
  .data_out(blk_fifo_0_data_out),
  .empty(blk_fifo_0_empty),
  .full(blk_fifo_0_full)
);

reg_fifo_depth_2_w_32_afd_2 blk_fifo_1 (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(blk_fifo_1_data_in),
  .flush(flush),
  .pop(pop_blk[1]),
  .push(push_blk[1]),
  .rst_n(rst_n),
  .data_out(blk_fifo_1_data_out),
  .empty(blk_fifo_1_empty),
  .full(blk_fifo_1_full)
);

arbiter_4_in_RR_algo rr_arbiter (
  .clk(gclk),
  .clk_en(clk_en),
  .flush(flush),
  .request_in(base_rr),
  .resource_ready(rr_arbiter_resource_ready),
  .rst_n(rst_n),
  .grant_out(mem_acq)
);

endmodule   // buffet_like_16

module fiber_access_16 (
  input logic [1:0] [3:0] buffet_buffet_capacity_log,
  input logic [3:0] [15:0] buffet_data_from_mem_lifted,
  input logic buffet_tile_en,
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic read_scanner_block_mode,
  input logic read_scanner_block_rd_out_ready,
  input logic read_scanner_coord_out_ready,
  input logic read_scanner_dense,
  input logic [15:0] read_scanner_dim_size,
  input logic read_scanner_do_repeat,
  input logic [15:0] read_scanner_inner_dim_offset,
  input logic read_scanner_lookup,
  input logic read_scanner_pos_out_ready,
  input logic [15:0] read_scanner_repeat_factor,
  input logic read_scanner_repeat_outer_inner_n,
  input logic read_scanner_root,
  input logic read_scanner_spacc_mode,
  input logic [15:0] read_scanner_stop_lvl,
  input logic read_scanner_tile_en,
  input logic [16:0] read_scanner_us_pos_in,
  input logic read_scanner_us_pos_in_valid,
  input logic rst_n,
  input logic tile_en,
  input logic [16:0] write_scanner_addr_in,
  input logic write_scanner_addr_in_valid,
  input logic write_scanner_block_mode,
  input logic [16:0] write_scanner_block_wr_in,
  input logic write_scanner_block_wr_in_valid,
  input logic write_scanner_compressed,
  input logic [16:0] write_scanner_data_in,
  input logic write_scanner_data_in_valid,
  input logic write_scanner_init_blank,
  input logic write_scanner_lowest_level,
  input logic write_scanner_spacc_mode,
  input logic [15:0] write_scanner_stop_lvl,
  input logic write_scanner_tile_en,
  output logic [8:0] buffet_addr_to_mem_lifted,
  output logic [3:0] [15:0] buffet_data_to_mem_lifted,
  output logic buffet_ren_to_mem_lifted,
  output logic buffet_wen_to_mem_lifted,
  output logic [16:0] read_scanner_block_rd_out,
  output logic read_scanner_block_rd_out_valid,
  output logic [16:0] read_scanner_coord_out,
  output logic read_scanner_coord_out_valid,
  output logic [16:0] read_scanner_pos_out,
  output logic read_scanner_pos_out_valid,
  output logic read_scanner_us_pos_in_ready,
  output logic write_scanner_addr_in_ready,
  output logic write_scanner_block_wr_in_ready,
  output logic write_scanner_data_in_ready
);

logic [0:0][16:0] buffet_rd_ID;
logic buffet_rd_ID_ready;
logic buffet_rd_ID_valid;
logic [0:0][16:0] buffet_rd_addr;
logic buffet_rd_addr_ready;
logic buffet_rd_addr_valid;
logic [0:0][16:0] buffet_rd_op;
logic buffet_rd_op_ready;
logic buffet_rd_op_valid;
logic [0:0][16:0] buffet_rd_rsp_data;
logic buffet_rd_rsp_data_ready;
logic buffet_rd_rsp_data_valid;
logic [0:0][16:0] buffet_wr_ID;
logic buffet_wr_ID_ready;
logic buffet_wr_ID_valid;
logic [0:0][16:0] buffet_wr_addr;
logic buffet_wr_addr_ready;
logic buffet_wr_addr_valid;
logic [0:0][16:0] buffet_wr_data;
logic buffet_wr_data_ready;
logic buffet_wr_data_valid;
logic gclk;
assign gclk = clk & tile_en;
buffet_like_16 buffet (
  .buffet_capacity_log(buffet_buffet_capacity_log),
  .clk(gclk),
  .clk_en(clk_en),
  .data_from_mem(buffet_data_from_mem_lifted),
  .flush(flush),
  .rd_ID(buffet_rd_ID),
  .rd_ID_valid(buffet_rd_ID_valid),
  .rd_addr(buffet_rd_addr),
  .rd_addr_valid(buffet_rd_addr_valid),
  .rd_op(buffet_rd_op),
  .rd_op_valid(buffet_rd_op_valid),
  .rd_rsp_data_ready(buffet_rd_rsp_data_ready),
  .rst_n(rst_n),
  .tile_en(buffet_tile_en),
  .wr_ID(buffet_wr_ID),
  .wr_ID_valid(buffet_wr_ID_valid),
  .wr_addr(buffet_wr_addr),
  .wr_addr_valid(buffet_wr_addr_valid),
  .wr_data(buffet_wr_data),
  .wr_data_valid(buffet_wr_data_valid),
  .addr_to_mem(buffet_addr_to_mem_lifted),
  .data_to_mem(buffet_data_to_mem_lifted),
  .rd_ID_ready(buffet_rd_ID_ready),
  .rd_addr_ready(buffet_rd_addr_ready),
  .rd_op_ready(buffet_rd_op_ready),
  .rd_rsp_data(buffet_rd_rsp_data),
  .rd_rsp_data_valid(buffet_rd_rsp_data_valid),
  .ren_to_mem(buffet_ren_to_mem_lifted),
  .wen_to_mem(buffet_wen_to_mem_lifted),
  .wr_ID_ready(buffet_wr_ID_ready),
  .wr_addr_ready(buffet_wr_addr_ready),
  .wr_data_ready(buffet_wr_data_ready)
);

write_scanner write_scanner (
  .ID_out_ready(buffet_wr_ID_ready),
  .addr_in(write_scanner_addr_in),
  .addr_in_valid(write_scanner_addr_in_valid),
  .addr_out_ready(buffet_wr_addr_ready),
  .block_mode(write_scanner_block_mode),
  .block_wr_in(write_scanner_block_wr_in),
  .block_wr_in_valid(write_scanner_block_wr_in_valid),
  .clk(gclk),
  .clk_en(clk_en),
  .compressed(write_scanner_compressed),
  .data_in(write_scanner_data_in),
  .data_in_valid(write_scanner_data_in_valid),
  .data_out_ready(buffet_wr_data_ready),
  .flush(flush),
  .init_blank(write_scanner_init_blank),
  .lowest_level(write_scanner_lowest_level),
  .rst_n(rst_n),
  .spacc_mode(write_scanner_spacc_mode),
  .stop_lvl(write_scanner_stop_lvl),
  .tile_en(write_scanner_tile_en),
  .ID_out(buffet_wr_ID),
  .ID_out_valid(buffet_wr_ID_valid),
  .addr_in_ready(write_scanner_addr_in_ready),
  .addr_out(buffet_wr_addr),
  .addr_out_valid(buffet_wr_addr_valid),
  .block_wr_in_ready(write_scanner_block_wr_in_ready),
  .data_in_ready(write_scanner_data_in_ready),
  .data_out(buffet_wr_data),
  .data_out_valid(buffet_wr_data_valid)
);

scanner_pipe read_scanner (
  .ID_out_ready(buffet_rd_ID_ready),
  .addr_out_ready(buffet_rd_addr_ready),
  .block_mode(read_scanner_block_mode),
  .block_rd_out_ready(read_scanner_block_rd_out_ready),
  .clk(gclk),
  .clk_en(clk_en),
  .coord_out_ready(read_scanner_coord_out_ready),
  .dense(read_scanner_dense),
  .dim_size(read_scanner_dim_size),
  .do_repeat(read_scanner_do_repeat),
  .flush(flush),
  .inner_dim_offset(read_scanner_inner_dim_offset),
  .lookup(read_scanner_lookup),
  .op_out_ready(buffet_rd_op_ready),
  .pos_out_ready(read_scanner_pos_out_ready),
  .rd_rsp_data_in(buffet_rd_rsp_data),
  .rd_rsp_data_in_valid(buffet_rd_rsp_data_valid),
  .repeat_factor(read_scanner_repeat_factor),
  .repeat_outer_inner_n(read_scanner_repeat_outer_inner_n),
  .root(read_scanner_root),
  .rst_n(rst_n),
  .spacc_mode(read_scanner_spacc_mode),
  .stop_lvl(read_scanner_stop_lvl),
  .tile_en(read_scanner_tile_en),
  .us_pos_in(read_scanner_us_pos_in),
  .us_pos_in_valid(read_scanner_us_pos_in_valid),
  .ID_out(buffet_rd_ID),
  .ID_out_valid(buffet_rd_ID_valid),
  .addr_out(buffet_rd_addr),
  .addr_out_valid(buffet_rd_addr_valid),
  .block_rd_out(read_scanner_block_rd_out),
  .block_rd_out_valid(read_scanner_block_rd_out_valid),
  .coord_out(read_scanner_coord_out),
  .coord_out_valid(read_scanner_coord_out_valid),
  .op_out(buffet_rd_op),
  .op_out_valid(buffet_rd_op_valid),
  .pos_out(read_scanner_pos_out),
  .pos_out_valid(read_scanner_pos_out_valid),
  .rd_rsp_data_in_ready(buffet_rd_rsp_data_ready),
  .us_pos_in_ready(read_scanner_us_pos_in_ready)
);

endmodule   // fiber_access_16

module fiber_access_16_flat (
  input logic clk,
  input logic clk_en,
  input logic [3:0] fiber_access_16_inst_buffet_buffet_capacity_log_0,
  input logic [3:0] fiber_access_16_inst_buffet_buffet_capacity_log_1,
  input logic [3:0] [15:0] fiber_access_16_inst_buffet_data_from_mem_lifted_lifted,
  input logic fiber_access_16_inst_buffet_tile_en,
  input logic fiber_access_16_inst_read_scanner_block_mode,
  input logic fiber_access_16_inst_read_scanner_dense,
  input logic [15:0] fiber_access_16_inst_read_scanner_dim_size,
  input logic fiber_access_16_inst_read_scanner_do_repeat,
  input logic [15:0] fiber_access_16_inst_read_scanner_inner_dim_offset,
  input logic fiber_access_16_inst_read_scanner_lookup,
  input logic [15:0] fiber_access_16_inst_read_scanner_repeat_factor,
  input logic fiber_access_16_inst_read_scanner_repeat_outer_inner_n,
  input logic fiber_access_16_inst_read_scanner_root,
  input logic fiber_access_16_inst_read_scanner_spacc_mode,
  input logic [15:0] fiber_access_16_inst_read_scanner_stop_lvl,
  input logic fiber_access_16_inst_read_scanner_tile_en,
  input logic fiber_access_16_inst_tile_en,
  input logic fiber_access_16_inst_write_scanner_block_mode,
  input logic fiber_access_16_inst_write_scanner_compressed,
  input logic fiber_access_16_inst_write_scanner_init_blank,
  input logic fiber_access_16_inst_write_scanner_lowest_level,
  input logic fiber_access_16_inst_write_scanner_spacc_mode,
  input logic [15:0] fiber_access_16_inst_write_scanner_stop_lvl,
  input logic fiber_access_16_inst_write_scanner_tile_en,
  input logic flush,
  input logic read_scanner_block_rd_out_ready_f_,
  input logic read_scanner_coord_out_ready_f_,
  input logic read_scanner_pos_out_ready_f_,
  input logic [0:0] [16:0] read_scanner_us_pos_in_f_,
  input logic read_scanner_us_pos_in_valid_f_,
  input logic rst_n,
  input logic [0:0] [16:0] write_scanner_addr_in_f_,
  input logic write_scanner_addr_in_valid_f_,
  input logic [0:0] [16:0] write_scanner_block_wr_in_f_,
  input logic write_scanner_block_wr_in_valid_f_,
  input logic [0:0] [16:0] write_scanner_data_in_f_,
  input logic write_scanner_data_in_valid_f_,
  output logic [8:0] fiber_access_16_inst_buffet_addr_to_mem_lifted_lifted,
  output logic [3:0] [15:0] fiber_access_16_inst_buffet_data_to_mem_lifted_lifted,
  output logic fiber_access_16_inst_buffet_ren_to_mem_lifted_lifted,
  output logic fiber_access_16_inst_buffet_wen_to_mem_lifted_lifted,
  output logic [0:0] [16:0] read_scanner_block_rd_out_f_,
  output logic read_scanner_block_rd_out_valid_f_,
  output logic [0:0] [16:0] read_scanner_coord_out_f_,
  output logic read_scanner_coord_out_valid_f_,
  output logic [0:0] [16:0] read_scanner_pos_out_f_,
  output logic read_scanner_pos_out_valid_f_,
  output logic read_scanner_us_pos_in_ready_f_,
  output logic write_scanner_addr_in_ready_f_,
  output logic write_scanner_block_wr_in_ready_f_,
  output logic write_scanner_data_in_ready_f_
);

logic [1:0][3:0] fiber_access_16_inst_buffet_buffet_capacity_log;
assign fiber_access_16_inst_buffet_buffet_capacity_log[0] = fiber_access_16_inst_buffet_buffet_capacity_log_0;
assign fiber_access_16_inst_buffet_buffet_capacity_log[1] = fiber_access_16_inst_buffet_buffet_capacity_log_1;
fiber_access_16 fiber_access_16_inst (
  .buffet_buffet_capacity_log(fiber_access_16_inst_buffet_buffet_capacity_log),
  .buffet_data_from_mem_lifted(fiber_access_16_inst_buffet_data_from_mem_lifted_lifted),
  .buffet_tile_en(fiber_access_16_inst_buffet_tile_en),
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .read_scanner_block_mode(fiber_access_16_inst_read_scanner_block_mode),
  .read_scanner_block_rd_out_ready(read_scanner_block_rd_out_ready_f_),
  .read_scanner_coord_out_ready(read_scanner_coord_out_ready_f_),
  .read_scanner_dense(fiber_access_16_inst_read_scanner_dense),
  .read_scanner_dim_size(fiber_access_16_inst_read_scanner_dim_size),
  .read_scanner_do_repeat(fiber_access_16_inst_read_scanner_do_repeat),
  .read_scanner_inner_dim_offset(fiber_access_16_inst_read_scanner_inner_dim_offset),
  .read_scanner_lookup(fiber_access_16_inst_read_scanner_lookup),
  .read_scanner_pos_out_ready(read_scanner_pos_out_ready_f_),
  .read_scanner_repeat_factor(fiber_access_16_inst_read_scanner_repeat_factor),
  .read_scanner_repeat_outer_inner_n(fiber_access_16_inst_read_scanner_repeat_outer_inner_n),
  .read_scanner_root(fiber_access_16_inst_read_scanner_root),
  .read_scanner_spacc_mode(fiber_access_16_inst_read_scanner_spacc_mode),
  .read_scanner_stop_lvl(fiber_access_16_inst_read_scanner_stop_lvl),
  .read_scanner_tile_en(fiber_access_16_inst_read_scanner_tile_en),
  .read_scanner_us_pos_in(read_scanner_us_pos_in_f_),
  .read_scanner_us_pos_in_valid(read_scanner_us_pos_in_valid_f_),
  .rst_n(rst_n),
  .tile_en(fiber_access_16_inst_tile_en),
  .write_scanner_addr_in(write_scanner_addr_in_f_),
  .write_scanner_addr_in_valid(write_scanner_addr_in_valid_f_),
  .write_scanner_block_mode(fiber_access_16_inst_write_scanner_block_mode),
  .write_scanner_block_wr_in(write_scanner_block_wr_in_f_),
  .write_scanner_block_wr_in_valid(write_scanner_block_wr_in_valid_f_),
  .write_scanner_compressed(fiber_access_16_inst_write_scanner_compressed),
  .write_scanner_data_in(write_scanner_data_in_f_),
  .write_scanner_data_in_valid(write_scanner_data_in_valid_f_),
  .write_scanner_init_blank(fiber_access_16_inst_write_scanner_init_blank),
  .write_scanner_lowest_level(fiber_access_16_inst_write_scanner_lowest_level),
  .write_scanner_spacc_mode(fiber_access_16_inst_write_scanner_spacc_mode),
  .write_scanner_stop_lvl(fiber_access_16_inst_write_scanner_stop_lvl),
  .write_scanner_tile_en(fiber_access_16_inst_write_scanner_tile_en),
  .buffet_addr_to_mem_lifted(fiber_access_16_inst_buffet_addr_to_mem_lifted_lifted),
  .buffet_data_to_mem_lifted(fiber_access_16_inst_buffet_data_to_mem_lifted_lifted),
  .buffet_ren_to_mem_lifted(fiber_access_16_inst_buffet_ren_to_mem_lifted_lifted),
  .buffet_wen_to_mem_lifted(fiber_access_16_inst_buffet_wen_to_mem_lifted_lifted),
  .read_scanner_block_rd_out(read_scanner_block_rd_out_f_),
  .read_scanner_block_rd_out_valid(read_scanner_block_rd_out_valid_f_),
  .read_scanner_coord_out(read_scanner_coord_out_f_),
  .read_scanner_coord_out_valid(read_scanner_coord_out_valid_f_),
  .read_scanner_pos_out(read_scanner_pos_out_f_),
  .read_scanner_pos_out_valid(read_scanner_pos_out_valid_f_),
  .read_scanner_us_pos_in_ready(read_scanner_us_pos_in_ready_f_),
  .write_scanner_addr_in_ready(write_scanner_addr_in_ready_f_),
  .write_scanner_block_wr_in_ready(write_scanner_block_wr_in_ready_f_),
  .write_scanner_data_in_ready(write_scanner_data_in_ready_f_)
);

endmodule   // fiber_access_16_flat

module for_loop_3_11 #(
  parameter CONFIG_WIDTH = 5'hB,
  parameter ITERATOR_SUPPORT = 3'h3,
  parameter ITERATOR_SUPPORT2 = 2'h2
)
(
  input logic clk,
  input logic clk_en,
  input logic [2:0] dimensionality,
  input logic flush,
  input logic [2:0] [10:0] ranges,
  input logic rst_n,
  input logic step,
  output logic [1:0] mux_sel_out,
  output logic restart
);

logic [2:0] clear;
logic [2:0][10:0] dim_counter;
logic done;
logic [2:0] inc;
logic [10:0] inced_cnt;
logic [2:0] max_value;
logic maxed_value;
logic [1:0] mux_sel;
assign mux_sel_out = mux_sel;
assign inced_cnt = dim_counter[mux_sel] + 11'h1;
assign maxed_value = (dim_counter[mux_sel] == ranges[mux_sel]) & inc[mux_sel];
always_comb begin
  mux_sel = 2'h0;
  done = 1'h0;
  if (~done) begin
    if ((~max_value[0]) & (dimensionality > 3'h0)) begin
      mux_sel = 2'h0;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[1]) & (dimensionality > 3'h1)) begin
      mux_sel = 2'h1;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[2]) & (dimensionality > 3'h2)) begin
      mux_sel = 2'h2;
      done = 1'h1;
    end
  end
end
always_comb begin
  clear[0] = 1'h0;
  if (((mux_sel > 2'h0) | (~done)) & step) begin
    clear[0] = 1'h1;
  end
end
always_comb begin
  inc[0] = 1'h0;
  if ((5'h0 == 5'h0) & step & (dimensionality > 3'h0)) begin
    inc[0] = 1'h1;
  end
  else if ((mux_sel == 2'h0) & step & (dimensionality > 3'h0)) begin
    inc[0] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[0] <= 11'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[0] <= 11'h0;
    end
    else if (clear[0]) begin
      dim_counter[0] <= 11'h0;
    end
    else if (inc[0]) begin
      dim_counter[0] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[0] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[0] <= 1'h0;
    end
    else if (clear[0]) begin
      max_value[0] <= 1'h0;
    end
    else if (inc[0]) begin
      max_value[0] <= maxed_value;
    end
  end
end
always_comb begin
  clear[1] = 1'h0;
  if (((mux_sel > 2'h1) | (~done)) & step) begin
    clear[1] = 1'h1;
  end
end
always_comb begin
  inc[1] = 1'h0;
  if ((5'h1 == 5'h0) & step & (dimensionality > 3'h1)) begin
    inc[1] = 1'h1;
  end
  else if ((mux_sel == 2'h1) & step & (dimensionality > 3'h1)) begin
    inc[1] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[1] <= 11'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[1] <= 11'h0;
    end
    else if (clear[1]) begin
      dim_counter[1] <= 11'h0;
    end
    else if (inc[1]) begin
      dim_counter[1] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[1] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[1] <= 1'h0;
    end
    else if (clear[1]) begin
      max_value[1] <= 1'h0;
    end
    else if (inc[1]) begin
      max_value[1] <= maxed_value;
    end
  end
end
always_comb begin
  clear[2] = 1'h0;
  if (((mux_sel > 2'h2) | (~done)) & step) begin
    clear[2] = 1'h1;
  end
end
always_comb begin
  inc[2] = 1'h0;
  if ((5'h2 == 5'h0) & step & (dimensionality > 3'h2)) begin
    inc[2] = 1'h1;
  end
  else if ((mux_sel == 2'h2) & step & (dimensionality > 3'h2)) begin
    inc[2] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[2] <= 11'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[2] <= 11'h0;
    end
    else if (clear[2]) begin
      dim_counter[2] <= 11'h0;
    end
    else if (inc[2]) begin
      dim_counter[2] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[2] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[2] <= 1'h0;
    end
    else if (clear[2]) begin
      max_value[2] <= 1'h0;
    end
    else if (inc[2]) begin
      max_value[2] <= maxed_value;
    end
  end
end
assign restart = step & (~done);
endmodule   // for_loop_3_11

module for_loop_6_11 #(
  parameter CONFIG_WIDTH = 5'hB,
  parameter ITERATOR_SUPPORT = 4'h6,
  parameter ITERATOR_SUPPORT2 = 2'h2
)
(
  input logic clk,
  input logic clk_en,
  input logic [3:0] dimensionality,
  input logic flush,
  input logic [5:0] [10:0] ranges,
  input logic rst_n,
  input logic step,
  output logic [2:0] mux_sel_out,
  output logic restart
);

logic [5:0] clear;
logic [5:0][10:0] dim_counter;
logic done;
logic [5:0] inc;
logic [10:0] inced_cnt;
logic [5:0] max_value;
logic maxed_value;
logic [2:0] mux_sel;
assign mux_sel_out = mux_sel;
assign inced_cnt = dim_counter[mux_sel] + 11'h1;
assign maxed_value = (dim_counter[mux_sel] == ranges[mux_sel]) & inc[mux_sel];
always_comb begin
  mux_sel = 3'h0;
  done = 1'h0;
  if (~done) begin
    if ((~max_value[0]) & (dimensionality > 4'h0)) begin
      mux_sel = 3'h0;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[1]) & (dimensionality > 4'h1)) begin
      mux_sel = 3'h1;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[2]) & (dimensionality > 4'h2)) begin
      mux_sel = 3'h2;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[3]) & (dimensionality > 4'h3)) begin
      mux_sel = 3'h3;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[4]) & (dimensionality > 4'h4)) begin
      mux_sel = 3'h4;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[5]) & (dimensionality > 4'h5)) begin
      mux_sel = 3'h5;
      done = 1'h1;
    end
  end
end
always_comb begin
  clear[0] = 1'h0;
  if (((mux_sel > 3'h0) | (~done)) & step) begin
    clear[0] = 1'h1;
  end
end
always_comb begin
  inc[0] = 1'h0;
  if ((5'h0 == 5'h0) & step & (dimensionality > 4'h0)) begin
    inc[0] = 1'h1;
  end
  else if ((mux_sel == 3'h0) & step & (dimensionality > 4'h0)) begin
    inc[0] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[0] <= 11'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[0] <= 11'h0;
    end
    else if (clear[0]) begin
      dim_counter[0] <= 11'h0;
    end
    else if (inc[0]) begin
      dim_counter[0] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[0] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[0] <= 1'h0;
    end
    else if (clear[0]) begin
      max_value[0] <= 1'h0;
    end
    else if (inc[0]) begin
      max_value[0] <= maxed_value;
    end
  end
end
always_comb begin
  clear[1] = 1'h0;
  if (((mux_sel > 3'h1) | (~done)) & step) begin
    clear[1] = 1'h1;
  end
end
always_comb begin
  inc[1] = 1'h0;
  if ((5'h1 == 5'h0) & step & (dimensionality > 4'h1)) begin
    inc[1] = 1'h1;
  end
  else if ((mux_sel == 3'h1) & step & (dimensionality > 4'h1)) begin
    inc[1] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[1] <= 11'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[1] <= 11'h0;
    end
    else if (clear[1]) begin
      dim_counter[1] <= 11'h0;
    end
    else if (inc[1]) begin
      dim_counter[1] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[1] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[1] <= 1'h0;
    end
    else if (clear[1]) begin
      max_value[1] <= 1'h0;
    end
    else if (inc[1]) begin
      max_value[1] <= maxed_value;
    end
  end
end
always_comb begin
  clear[2] = 1'h0;
  if (((mux_sel > 3'h2) | (~done)) & step) begin
    clear[2] = 1'h1;
  end
end
always_comb begin
  inc[2] = 1'h0;
  if ((5'h2 == 5'h0) & step & (dimensionality > 4'h2)) begin
    inc[2] = 1'h1;
  end
  else if ((mux_sel == 3'h2) & step & (dimensionality > 4'h2)) begin
    inc[2] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[2] <= 11'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[2] <= 11'h0;
    end
    else if (clear[2]) begin
      dim_counter[2] <= 11'h0;
    end
    else if (inc[2]) begin
      dim_counter[2] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[2] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[2] <= 1'h0;
    end
    else if (clear[2]) begin
      max_value[2] <= 1'h0;
    end
    else if (inc[2]) begin
      max_value[2] <= maxed_value;
    end
  end
end
always_comb begin
  clear[3] = 1'h0;
  if (((mux_sel > 3'h3) | (~done)) & step) begin
    clear[3] = 1'h1;
  end
end
always_comb begin
  inc[3] = 1'h0;
  if ((5'h3 == 5'h0) & step & (dimensionality > 4'h3)) begin
    inc[3] = 1'h1;
  end
  else if ((mux_sel == 3'h3) & step & (dimensionality > 4'h3)) begin
    inc[3] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[3] <= 11'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[3] <= 11'h0;
    end
    else if (clear[3]) begin
      dim_counter[3] <= 11'h0;
    end
    else if (inc[3]) begin
      dim_counter[3] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[3] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[3] <= 1'h0;
    end
    else if (clear[3]) begin
      max_value[3] <= 1'h0;
    end
    else if (inc[3]) begin
      max_value[3] <= maxed_value;
    end
  end
end
always_comb begin
  clear[4] = 1'h0;
  if (((mux_sel > 3'h4) | (~done)) & step) begin
    clear[4] = 1'h1;
  end
end
always_comb begin
  inc[4] = 1'h0;
  if ((5'h4 == 5'h0) & step & (dimensionality > 4'h4)) begin
    inc[4] = 1'h1;
  end
  else if ((mux_sel == 3'h4) & step & (dimensionality > 4'h4)) begin
    inc[4] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[4] <= 11'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[4] <= 11'h0;
    end
    else if (clear[4]) begin
      dim_counter[4] <= 11'h0;
    end
    else if (inc[4]) begin
      dim_counter[4] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[4] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[4] <= 1'h0;
    end
    else if (clear[4]) begin
      max_value[4] <= 1'h0;
    end
    else if (inc[4]) begin
      max_value[4] <= maxed_value;
    end
  end
end
always_comb begin
  clear[5] = 1'h0;
  if (((mux_sel > 3'h5) | (~done)) & step) begin
    clear[5] = 1'h1;
  end
end
always_comb begin
  inc[5] = 1'h0;
  if ((5'h5 == 5'h0) & step & (dimensionality > 4'h5)) begin
    inc[5] = 1'h1;
  end
  else if ((mux_sel == 3'h5) & step & (dimensionality > 4'h5)) begin
    inc[5] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[5] <= 11'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[5] <= 11'h0;
    end
    else if (clear[5]) begin
      dim_counter[5] <= 11'h0;
    end
    else if (inc[5]) begin
      dim_counter[5] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[5] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[5] <= 1'h0;
    end
    else if (clear[5]) begin
      max_value[5] <= 1'h0;
    end
    else if (inc[5]) begin
      max_value[5] <= maxed_value;
    end
  end
end
assign restart = step & (~done);
endmodule   // for_loop_6_11

module reg_fifo_depth_0_w_16_afd_2 (
  input logic clk,
  input logic clk_en,
  input logic [0:0] [15:0] data_in,
  input logic flush,
  input logic pop,
  input logic push,
  input logic rst_n,
  output logic almost_full,
  output logic [0:0] [15:0] data_out,
  output logic empty,
  output logic full,
  output logic valid
);

assign data_out = data_in;
assign valid = push;
assign empty = ~push;
assign full = ~pop;
assign almost_full = ~pop;
endmodule   // reg_fifo_depth_0_w_16_afd_2

module reg_fifo_depth_2_w_16_afd_2 (
  input logic clk,
  input logic clk_en,
  input logic [0:0] [15:0] data_in,
  input logic flush,
  input logic pop,
  input logic push,
  input logic rst_n,
  output logic almost_full,
  output logic [0:0] [15:0] data_out,
  output logic empty,
  output logic full,
  output logic valid
);

logic [1:0] num_items;
logic passthru;
logic rd_ptr;
logic read;
logic [1:0][0:0][15:0] reg_array;
logic wr_ptr;
logic write;
assign full = num_items == 2'h2;
assign almost_full = num_items >= 2'h0;
assign empty = num_items == 2'h0;
assign read = pop & (~passthru) & (~empty);
assign passthru = 1'h0;
assign write = push & (~passthru) & (~full);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_items <= 2'h0;
  end
  else if (flush) begin
    num_items <= 2'h0;
  end
  else if (clk_en) begin
    if (write & (~read)) begin
      num_items <= num_items + 2'h1;
    end
    else if ((~write) & read) begin
      num_items <= num_items - 2'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    reg_array <= 32'h0;
  end
  else if (flush) begin
    reg_array <= 32'h0;
  end
  else if (clk_en) begin
    if (write) begin
      reg_array[wr_ptr] <= data_in;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    wr_ptr <= 1'h0;
  end
  else if (flush) begin
    wr_ptr <= 1'h0;
  end
  else if (clk_en) begin
    if (write) begin
      if (wr_ptr == 1'h1) begin
        wr_ptr <= 1'h0;
      end
      else wr_ptr <= wr_ptr + 1'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    rd_ptr <= 1'h0;
  end
  else if (flush) begin
    rd_ptr <= 1'h0;
  end
  else if (clk_en) begin
    if (read) begin
      rd_ptr <= rd_ptr + 1'h1;
    end
  end
end
always_comb begin
  if (passthru) begin
    data_out = data_in;
  end
  else data_out = reg_array[rd_ptr];
end
always_comb begin
  valid = (~empty) | passthru;
end
endmodule   // reg_fifo_depth_2_w_16_afd_2

module reg_fifo_depth_2_w_17_afd_1 (
  input logic clk,
  input logic clk_en,
  input logic [0:0] [16:0] data_in,
  input logic flush,
  input logic pop,
  input logic push,
  input logic rst_n,
  output logic almost_full,
  output logic [0:0] [16:0] data_out,
  output logic empty,
  output logic full,
  output logic valid
);

logic [1:0] num_items;
logic passthru;
logic rd_ptr;
logic read;
logic [1:0][0:0][16:0] reg_array;
logic wr_ptr;
logic write;
assign full = num_items == 2'h2;
assign almost_full = num_items >= 2'h1;
assign empty = num_items == 2'h0;
assign read = pop & (~passthru) & (~empty);
assign passthru = 1'h0;
assign write = push & (~passthru) & (~full);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_items <= 2'h0;
  end
  else if (flush) begin
    num_items <= 2'h0;
  end
  else if (clk_en) begin
    if (write & (~read)) begin
      num_items <= num_items + 2'h1;
    end
    else if ((~write) & read) begin
      num_items <= num_items - 2'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    reg_array <= 34'h0;
  end
  else if (flush) begin
    reg_array <= 34'h0;
  end
  else if (clk_en) begin
    if (write) begin
      reg_array[wr_ptr] <= data_in;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    wr_ptr <= 1'h0;
  end
  else if (flush) begin
    wr_ptr <= 1'h0;
  end
  else if (clk_en) begin
    if (write) begin
      if (wr_ptr == 1'h1) begin
        wr_ptr <= 1'h0;
      end
      else wr_ptr <= wr_ptr + 1'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    rd_ptr <= 1'h0;
  end
  else if (flush) begin
    rd_ptr <= 1'h0;
  end
  else if (clk_en) begin
    if (read) begin
      rd_ptr <= rd_ptr + 1'h1;
    end
  end
end
always_comb begin
  if (passthru) begin
    data_out = data_in;
  end
  else data_out = reg_array[rd_ptr];
end
always_comb begin
  valid = (~empty) | passthru;
end
endmodule   // reg_fifo_depth_2_w_17_afd_1

module reg_fifo_depth_2_w_32_afd_2 (
  input logic clk,
  input logic clk_en,
  input logic [0:0] [31:0] data_in,
  input logic flush,
  input logic pop,
  input logic push,
  input logic rst_n,
  output logic almost_full,
  output logic [0:0] [31:0] data_out,
  output logic empty,
  output logic full,
  output logic valid
);

logic [1:0] num_items;
logic passthru;
logic rd_ptr;
logic read;
logic [1:0][0:0][31:0] reg_array;
logic wr_ptr;
logic write;
assign full = num_items == 2'h2;
assign almost_full = num_items >= 2'h0;
assign empty = num_items == 2'h0;
assign read = pop & (~passthru) & (~empty);
assign passthru = 1'h0;
assign write = push & (~passthru) & (~full);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_items <= 2'h0;
  end
  else if (flush) begin
    num_items <= 2'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (clk_en) begin
        if (write & (~read)) begin
          num_items <= num_items + 2'h1;
        end
        else if ((~write) & read) begin
          num_items <= num_items - 2'h1;
        end
      end
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    reg_array <= 64'h0;
  end
  else if (flush) begin
    reg_array <= 64'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (clk_en) begin
        if (write) begin
          reg_array[wr_ptr] <= data_in;
        end
      end
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    wr_ptr <= 1'h0;
  end
  else if (flush) begin
    wr_ptr <= 1'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (clk_en) begin
        if (write) begin
          if (wr_ptr == 1'h1) begin
            wr_ptr <= 1'h0;
          end
          else wr_ptr <= wr_ptr + 1'h1;
        end
      end
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    rd_ptr <= 1'h0;
  end
  else if (flush) begin
    rd_ptr <= 1'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (clk_en) begin
        if (read) begin
          rd_ptr <= rd_ptr + 1'h1;
        end
      end
    end
  end
end
always_comb begin
  if (passthru) begin
    data_out = data_in;
  end
  else data_out = reg_array[rd_ptr];
end
always_comb begin
  valid = (~empty) | passthru;
end
endmodule   // reg_fifo_depth_2_w_32_afd_2

module reservation_fifo_depth_8_w_17_num_per_1 (
  input logic clk,
  input logic clk_en,
  input logic [16:0] data_in_0,
  input logic [16:0] fill_data_in,
  input logic flush,
  input logic pop,
  input logic push_alloc,
  input logic push_fill,
  input logic push_reserve,
  input logic rst_n,
  output logic [16:0] data_out_0,
  output logic empty,
  output logic full,
  output logic valid
);

logic clr_item_ptr;
logic clr_read_ptr;
logic clr_write_ptr;
logic [0:0][16:0] data_in_packed;
logic [0:0][16:0] data_out;
logic enable_reserve_ptr;
logic inc_item_ptr;
logic inc_read_ptr;
logic inc_reserve_count;
logic inc_write_ptr;
logic item_ptr;
logic jump_next_0;
logic [2:0] next_0_valid;
logic [2:0] next_0_valid_d1;
logic [2:0] next_0_valid_high;
logic next_0_valid_high_done;
logic next_0_valid_high_found;
logic [2:0] next_0_valid_low;
logic next_0_valid_low_done;
logic next_0_valid_low_found;
logic [3:0] num_items;
logic read;
logic [2:0] read_ptr_addr;
logic [7:0][0:0][16:0] reg_array;
logic [15:0] reserve_count;
logic [2:0] reserve_ptr_val;
logic [7:0] valid_mask;
logic write_alloc;
logic write_fill;
logic [2:0] write_ptr_addr;
logic write_reserve;
logic write_reserve_final;
assign data_in_packed[0] = data_in_0;
assign data_out_0 = data_out[0];
assign item_ptr = 1'h0;
assign inc_item_ptr = push_reserve;
assign clr_item_ptr = push_reserve & (item_ptr == 1'h0);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    read_ptr_addr <= 3'h0;
  end
  else if (flush) begin
    read_ptr_addr <= 3'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (clr_read_ptr) begin
        read_ptr_addr <= 3'h0;
      end
      else if (inc_read_ptr) begin
        read_ptr_addr <= read_ptr_addr + 3'h1;
      end
    end
  end
end
assign inc_read_ptr = read;
assign clr_read_ptr = 1'h0;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    write_ptr_addr <= 3'h0;
  end
  else if (flush) begin
    write_ptr_addr <= 3'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (clr_write_ptr) begin
        write_ptr_addr <= 3'h0;
      end
      else if (inc_write_ptr) begin
        write_ptr_addr <= write_ptr_addr + 3'h1;
      end
    end
  end
end
assign inc_write_ptr = write_alloc | write_fill;
assign clr_write_ptr = 1'h0;
assign jump_next_0 = next_0_valid_high_found | next_0_valid_low_found;
assign enable_reserve_ptr = write_reserve_final | (write_fill & (reserve_ptr_val == write_ptr_addr));

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    next_0_valid_d1 <= 3'h0;
  end
  else if (flush) begin
    next_0_valid_d1 <= 3'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (1'h0) begin
        next_0_valid_d1 <= 3'h0;
      end
      else if (enable_reserve_ptr) begin
        next_0_valid_d1 <= next_0_valid;
      end
    end
  end
end
assign reserve_ptr_val = next_0_valid_d1;
assign next_0_valid = (write_fill & ((next_0_valid_d1 == write_ptr_addr) | ((~next_0_valid_high_found)
    & (~next_0_valid_low_found)) | (next_0_valid_high_found ? next_0_valid_high ==
    write_ptr_addr: next_0_valid_low == write_ptr_addr))) ? write_ptr_addr + 3'h1:
    ((~next_0_valid_high_found) & (~next_0_valid_low_found)) ? write_ptr_addr:
    next_0_valid_high_found ? next_0_valid_high: next_0_valid_low;
assign full = num_items == 4'h8;
assign empty = num_items == 4'h0;
assign write_fill = push_fill & push_alloc & (~full);
assign write_alloc = push_alloc & (~full);
assign write_reserve = inc_item_ptr;
assign write_reserve_final = clr_item_ptr;
assign read = pop & valid_mask[read_ptr_addr];

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_items <= 4'h0;
  end
  else if (flush) begin
    num_items <= 4'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (write_alloc & (~read)) begin
        num_items <= num_items + 4'h1;
      end
      else if ((~write_alloc) & read) begin
        num_items <= num_items - 4'h1;
      end
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    reg_array <= 136'h0;
  end
  else if (flush) begin
    reg_array <= 136'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (write_fill) begin
        reg_array[write_ptr_addr] <= fill_data_in;
      end
      if (write_reserve) begin
        reg_array[next_0_valid_d1] <= data_in_packed;
      end
    end
  end
end
always_comb begin
  data_out = reg_array[read_ptr_addr];
end
always_comb begin
  valid = valid_mask[read_ptr_addr];
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    valid_mask <= 8'h0;
  end
  else if (flush) begin
    valid_mask <= 8'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (write_fill) begin
        valid_mask[write_ptr_addr] <= 1'h1;
      end
      if (write_reserve_final) begin
        valid_mask[next_0_valid_d1] <= 1'h1;
      end
      if (read) begin
        valid_mask[read_ptr_addr] <= 1'h0;
      end
    end
  end
end
always_comb begin
  next_0_valid_high_found = 1'h0;
  next_0_valid_high = 3'h0;
  next_0_valid_high_done = 1'h0;
  if (~next_0_valid_high_done) begin
    if (next_0_valid_d1 < 3'h0) begin
      if (valid_mask[0] == 1'h0) begin
        next_0_valid_high_found = 1'h1;
        next_0_valid_high = 3'h0;
        next_0_valid_high_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_high_done) begin
    if (next_0_valid_d1 < 3'h1) begin
      if (valid_mask[1] == 1'h0) begin
        next_0_valid_high_found = 1'h1;
        next_0_valid_high = 3'h1;
        next_0_valid_high_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_high_done) begin
    if (next_0_valid_d1 < 3'h2) begin
      if (valid_mask[2] == 1'h0) begin
        next_0_valid_high_found = 1'h1;
        next_0_valid_high = 3'h2;
        next_0_valid_high_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_high_done) begin
    if (next_0_valid_d1 < 3'h3) begin
      if (valid_mask[3] == 1'h0) begin
        next_0_valid_high_found = 1'h1;
        next_0_valid_high = 3'h3;
        next_0_valid_high_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_high_done) begin
    if (next_0_valid_d1 < 3'h4) begin
      if (valid_mask[4] == 1'h0) begin
        next_0_valid_high_found = 1'h1;
        next_0_valid_high = 3'h4;
        next_0_valid_high_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_high_done) begin
    if (next_0_valid_d1 < 3'h5) begin
      if (valid_mask[5] == 1'h0) begin
        next_0_valid_high_found = 1'h1;
        next_0_valid_high = 3'h5;
        next_0_valid_high_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_high_done) begin
    if (next_0_valid_d1 < 3'h6) begin
      if (valid_mask[6] == 1'h0) begin
        next_0_valid_high_found = 1'h1;
        next_0_valid_high = 3'h6;
        next_0_valid_high_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_high_done) begin
    if (next_0_valid_d1 < 3'h7) begin
      if (valid_mask[7] == 1'h0) begin
        next_0_valid_high_found = 1'h1;
        next_0_valid_high = 3'h7;
        next_0_valid_high_done = 1'h1;
      end
    end
  end
end
always_comb begin
  next_0_valid_low_found = 1'h0;
  next_0_valid_low = 3'h0;
  next_0_valid_low_done = 1'h0;
  if (~next_0_valid_low_done) begin
    if (next_0_valid_d1 > 3'h0) begin
      if (valid_mask[0] == 1'h0) begin
        next_0_valid_low_found = 1'h1;
        next_0_valid_low = 3'h0;
        next_0_valid_low_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_low_done) begin
    if (next_0_valid_d1 > 3'h1) begin
      if (valid_mask[1] == 1'h0) begin
        next_0_valid_low_found = 1'h1;
        next_0_valid_low = 3'h1;
        next_0_valid_low_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_low_done) begin
    if (next_0_valid_d1 > 3'h2) begin
      if (valid_mask[2] == 1'h0) begin
        next_0_valid_low_found = 1'h1;
        next_0_valid_low = 3'h2;
        next_0_valid_low_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_low_done) begin
    if (next_0_valid_d1 > 3'h3) begin
      if (valid_mask[3] == 1'h0) begin
        next_0_valid_low_found = 1'h1;
        next_0_valid_low = 3'h3;
        next_0_valid_low_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_low_done) begin
    if (next_0_valid_d1 > 3'h4) begin
      if (valid_mask[4] == 1'h0) begin
        next_0_valid_low_found = 1'h1;
        next_0_valid_low = 3'h4;
        next_0_valid_low_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_low_done) begin
    if (next_0_valid_d1 > 3'h5) begin
      if (valid_mask[5] == 1'h0) begin
        next_0_valid_low_found = 1'h1;
        next_0_valid_low = 3'h5;
        next_0_valid_low_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_low_done) begin
    if (next_0_valid_d1 > 3'h6) begin
      if (valid_mask[6] == 1'h0) begin
        next_0_valid_low_found = 1'h1;
        next_0_valid_low = 3'h6;
        next_0_valid_low_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_low_done) begin
    if (next_0_valid_d1 > 3'h7) begin
      if (valid_mask[7] == 1'h0) begin
        next_0_valid_low_found = 1'h1;
        next_0_valid_low = 3'h7;
        next_0_valid_low_done = 1'h1;
      end
    end
  end
end
assign inc_reserve_count = write_alloc & (~write_fill);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    reserve_count <= 16'h0;
  end
  else if (flush) begin
    reserve_count <= 16'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (inc_reserve_count) begin
        reserve_count <= reserve_count + 16'h1;
      end
    end
  end
end
endmodule   // reservation_fifo_depth_8_w_17_num_per_1

module reservation_fifo_depth_8_w_17_num_per_2 (
  input logic clk,
  input logic clk_en,
  input logic [16:0] data_in_0,
  input logic [16:0] data_in_1,
  input logic [16:0] fill_data_in,
  input logic flush,
  input logic pop,
  input logic push_alloc,
  input logic push_fill,
  input logic push_reserve,
  input logic rst_n,
  output logic [16:0] data_out_0,
  output logic [16:0] data_out_1,
  output logic empty,
  output logic full,
  output logic valid
);

logic clr_item_ptr;
logic clr_read_ptr;
logic clr_write_ptr;
logic [1:0][16:0] data_in_packed;
logic [1:0][16:0] data_out;
logic enable_reserve_ptr;
logic inc_item_ptr;
logic inc_read_ptr;
logic inc_reserve_count;
logic inc_write_ptr;
logic item_ptr_addr;
logic jump_next_0;
logic [2:0] next_0_valid;
logic [2:0] next_0_valid_d1;
logic [2:0] next_0_valid_high;
logic next_0_valid_high_done;
logic next_0_valid_high_found;
logic [2:0] next_0_valid_low;
logic next_0_valid_low_done;
logic next_0_valid_low_found;
logic [3:0] num_items;
logic read;
logic [2:0] read_ptr_addr;
logic [7:0][1:0][16:0] reg_array;
logic [15:0] reserve_count;
logic [2:0] reserve_ptr_val;
logic [7:0] valid_mask;
logic write_alloc;
logic write_fill;
logic [2:0] write_ptr_addr;
logic write_reserve;
logic write_reserve_final;
assign data_in_packed[0] = data_in_0;
assign data_in_packed[1] = data_in_1;
assign data_out_0 = data_out[0];
assign data_out_1 = data_out[1];

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    item_ptr_addr <= 1'h0;
  end
  else if (flush) begin
    item_ptr_addr <= 1'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (clr_item_ptr) begin
        item_ptr_addr <= 1'h0;
      end
      else if (inc_item_ptr) begin
        item_ptr_addr <= item_ptr_addr + 1'h1;
      end
    end
  end
end
assign inc_item_ptr = push_reserve;
assign clr_item_ptr = push_reserve & (item_ptr_addr == 1'h1);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    read_ptr_addr <= 3'h0;
  end
  else if (flush) begin
    read_ptr_addr <= 3'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (clr_read_ptr) begin
        read_ptr_addr <= 3'h0;
      end
      else if (inc_read_ptr) begin
        read_ptr_addr <= read_ptr_addr + 3'h1;
      end
    end
  end
end
assign inc_read_ptr = read;
assign clr_read_ptr = 1'h0;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    write_ptr_addr <= 3'h0;
  end
  else if (flush) begin
    write_ptr_addr <= 3'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (clr_write_ptr) begin
        write_ptr_addr <= 3'h0;
      end
      else if (inc_write_ptr) begin
        write_ptr_addr <= write_ptr_addr + 3'h1;
      end
    end
  end
end
assign inc_write_ptr = write_alloc | write_fill;
assign clr_write_ptr = 1'h0;
assign jump_next_0 = next_0_valid_high_found | next_0_valid_low_found;
assign enable_reserve_ptr = write_reserve_final | (write_fill & (reserve_ptr_val == write_ptr_addr));

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    next_0_valid_d1 <= 3'h0;
  end
  else if (flush) begin
    next_0_valid_d1 <= 3'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (1'h0) begin
        next_0_valid_d1 <= 3'h0;
      end
      else if (enable_reserve_ptr) begin
        next_0_valid_d1 <= next_0_valid;
      end
    end
  end
end
assign reserve_ptr_val = next_0_valid_d1;
assign next_0_valid = (write_fill & ((next_0_valid_d1 == write_ptr_addr) | ((~next_0_valid_high_found)
    & (~next_0_valid_low_found)) | (next_0_valid_high_found ? next_0_valid_high ==
    write_ptr_addr: next_0_valid_low == write_ptr_addr))) ? write_ptr_addr + 3'h1:
    ((~next_0_valid_high_found) & (~next_0_valid_low_found)) ? write_ptr_addr:
    next_0_valid_high_found ? next_0_valid_high: next_0_valid_low;
assign full = num_items == 4'h8;
assign empty = num_items == 4'h0;
assign write_fill = push_fill & push_alloc & (~full);
assign write_alloc = push_alloc & (~full);
assign write_reserve = inc_item_ptr;
assign write_reserve_final = clr_item_ptr;
assign read = pop & valid_mask[read_ptr_addr];

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_items <= 4'h0;
  end
  else if (flush) begin
    num_items <= 4'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (write_alloc & (~read)) begin
        num_items <= num_items + 4'h1;
      end
      else if ((~write_alloc) & read) begin
        num_items <= num_items - 4'h1;
      end
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    reg_array <= 272'h0;
  end
  else if (flush) begin
    reg_array <= 272'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (write_fill) begin
        reg_array[write_ptr_addr][0] <= fill_data_in;
      end
      if (write_reserve) begin
        reg_array[next_0_valid_d1][item_ptr_addr] <= data_in_packed[item_ptr_addr];
      end
    end
  end
end
always_comb begin
  data_out = reg_array[read_ptr_addr];
end
always_comb begin
  valid = valid_mask[read_ptr_addr];
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    valid_mask <= 8'h0;
  end
  else if (flush) begin
    valid_mask <= 8'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (write_fill) begin
        valid_mask[write_ptr_addr] <= 1'h1;
      end
      if (write_reserve_final) begin
        valid_mask[next_0_valid_d1] <= 1'h1;
      end
      if (read) begin
        valid_mask[read_ptr_addr] <= 1'h0;
      end
    end
  end
end
always_comb begin
  next_0_valid_high_found = 1'h0;
  next_0_valid_high = 3'h0;
  next_0_valid_high_done = 1'h0;
  if (~next_0_valid_high_done) begin
    if (next_0_valid_d1 < 3'h0) begin
      if (valid_mask[0] == 1'h0) begin
        next_0_valid_high_found = 1'h1;
        next_0_valid_high = 3'h0;
        next_0_valid_high_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_high_done) begin
    if (next_0_valid_d1 < 3'h1) begin
      if (valid_mask[1] == 1'h0) begin
        next_0_valid_high_found = 1'h1;
        next_0_valid_high = 3'h1;
        next_0_valid_high_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_high_done) begin
    if (next_0_valid_d1 < 3'h2) begin
      if (valid_mask[2] == 1'h0) begin
        next_0_valid_high_found = 1'h1;
        next_0_valid_high = 3'h2;
        next_0_valid_high_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_high_done) begin
    if (next_0_valid_d1 < 3'h3) begin
      if (valid_mask[3] == 1'h0) begin
        next_0_valid_high_found = 1'h1;
        next_0_valid_high = 3'h3;
        next_0_valid_high_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_high_done) begin
    if (next_0_valid_d1 < 3'h4) begin
      if (valid_mask[4] == 1'h0) begin
        next_0_valid_high_found = 1'h1;
        next_0_valid_high = 3'h4;
        next_0_valid_high_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_high_done) begin
    if (next_0_valid_d1 < 3'h5) begin
      if (valid_mask[5] == 1'h0) begin
        next_0_valid_high_found = 1'h1;
        next_0_valid_high = 3'h5;
        next_0_valid_high_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_high_done) begin
    if (next_0_valid_d1 < 3'h6) begin
      if (valid_mask[6] == 1'h0) begin
        next_0_valid_high_found = 1'h1;
        next_0_valid_high = 3'h6;
        next_0_valid_high_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_high_done) begin
    if (next_0_valid_d1 < 3'h7) begin
      if (valid_mask[7] == 1'h0) begin
        next_0_valid_high_found = 1'h1;
        next_0_valid_high = 3'h7;
        next_0_valid_high_done = 1'h1;
      end
    end
  end
end
always_comb begin
  next_0_valid_low_found = 1'h0;
  next_0_valid_low = 3'h0;
  next_0_valid_low_done = 1'h0;
  if (~next_0_valid_low_done) begin
    if (next_0_valid_d1 > 3'h0) begin
      if (valid_mask[0] == 1'h0) begin
        next_0_valid_low_found = 1'h1;
        next_0_valid_low = 3'h0;
        next_0_valid_low_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_low_done) begin
    if (next_0_valid_d1 > 3'h1) begin
      if (valid_mask[1] == 1'h0) begin
        next_0_valid_low_found = 1'h1;
        next_0_valid_low = 3'h1;
        next_0_valid_low_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_low_done) begin
    if (next_0_valid_d1 > 3'h2) begin
      if (valid_mask[2] == 1'h0) begin
        next_0_valid_low_found = 1'h1;
        next_0_valid_low = 3'h2;
        next_0_valid_low_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_low_done) begin
    if (next_0_valid_d1 > 3'h3) begin
      if (valid_mask[3] == 1'h0) begin
        next_0_valid_low_found = 1'h1;
        next_0_valid_low = 3'h3;
        next_0_valid_low_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_low_done) begin
    if (next_0_valid_d1 > 3'h4) begin
      if (valid_mask[4] == 1'h0) begin
        next_0_valid_low_found = 1'h1;
        next_0_valid_low = 3'h4;
        next_0_valid_low_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_low_done) begin
    if (next_0_valid_d1 > 3'h5) begin
      if (valid_mask[5] == 1'h0) begin
        next_0_valid_low_found = 1'h1;
        next_0_valid_low = 3'h5;
        next_0_valid_low_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_low_done) begin
    if (next_0_valid_d1 > 3'h6) begin
      if (valid_mask[6] == 1'h0) begin
        next_0_valid_low_found = 1'h1;
        next_0_valid_low = 3'h6;
        next_0_valid_low_done = 1'h1;
      end
    end
  end
  if (~next_0_valid_low_done) begin
    if (next_0_valid_d1 > 3'h7) begin
      if (valid_mask[7] == 1'h0) begin
        next_0_valid_low_found = 1'h1;
        next_0_valid_low = 3'h7;
        next_0_valid_low_done = 1'h1;
      end
    end
  end
end
assign inc_reserve_count = write_alloc & (~write_fill);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    reserve_count <= 16'h0;
  end
  else if (flush) begin
    reserve_count <= 16'h0;
  end
  else if (clk_en) begin
    if (clk_en) begin
      if (inc_reserve_count) begin
        reserve_count <= reserve_count + 16'h1;
      end
    end
  end
end
endmodule   // reservation_fifo_depth_8_w_17_num_per_2

module scanner_pipe (
  input logic ID_out_ready,
  input logic addr_out_ready,
  input logic block_mode,
  input logic block_rd_out_ready,
  input logic clk,
  input logic clk_en,
  input logic coord_out_ready,
  input logic dense,
  input logic [15:0] dim_size,
  input logic do_repeat,
  input logic flush,
  input logic [15:0] inner_dim_offset,
  input logic lookup,
  input logic op_out_ready,
  input logic pos_out_ready,
  input logic [0:0] [16:0] rd_rsp_data_in,
  input logic rd_rsp_data_in_valid,
  input logic [15:0] repeat_factor,
  input logic repeat_outer_inner_n,
  input logic root,
  input logic rst_n,
  input logic spacc_mode,
  input logic [15:0] stop_lvl,
  input logic tile_en,
  input logic [16:0] us_pos_in,
  input logic us_pos_in_valid,
  output logic [0:0] [16:0] ID_out,
  output logic ID_out_valid,
  output logic [0:0] [16:0] addr_out,
  output logic addr_out_valid,
  output logic [16:0] block_rd_out,
  output logic block_rd_out_valid,
  output logic [16:0] coord_out,
  output logic coord_out_valid,
  output logic [0:0] [16:0] op_out,
  output logic op_out_valid,
  output logic [16:0] pos_out,
  output logic pos_out_valid,
  output logic rd_rsp_data_in_ready,
  output logic us_pos_in_ready
);

typedef enum logic[3:0] {
  BLOCK_1_RD = 4'h0,
  BLOCK_1_SIZE_REC = 4'h1,
  BLOCK_1_SIZE_REQ = 4'h2,
  BLOCK_2_RD = 4'h3,
  BLOCK_2_SIZE_REC = 4'h4,
  BLOCK_2_SIZE_REQ = 4'h5,
  DENSE_STRM = 4'h6,
  DONE_CRD = 4'h7,
  FREE_CRD = 4'h8,
  FREE_CRD2 = 4'h9,
  PASS_DONE_CRD = 4'hA,
  READOUT_SYNC_LOCK = 4'hB,
  SEQ_STRM = 4'hC,
  START_CRD = 4'hD
} scan_seq_crd_state;
typedef enum logic[3:0] {
  DONE_SEG = 4'h0,
  FREE_SEG = 4'h1,
  INJECT_0 = 4'h2,
  INJECT_DONE = 4'h3,
  INJECT_ROUTING = 4'h4,
  LOOKUP = 4'h5,
  PASS_DONE_SEG = 4'h6,
  PASS_STOP_SEG = 4'h7,
  READ = 4'h8,
  READ_ALT = 4'h9,
  START_SEG = 4'hA
} scan_seq_seg_state;
logic [0:0][16:0] ID_out_fifo_data_in;
logic ID_out_fifo_empty;
logic ID_out_fifo_full;
logic ID_out_fifo_push;
logic [0:0][15:0] ID_out_to_fifo;
logic [15:0] READS_MADE;
logic [15:0] READS_REC_CRD_READ;
logic [0:0][16:0] addr_out_fifo_data_in;
logic addr_out_fifo_empty;
logic addr_out_fifo_full;
logic addr_out_fifo_push;
logic [0:0][15:0] addr_out_to_fifo;
logic [1:0] base_rr;
logic block_rd_fifo_empty;
logic block_rd_fifo_full;
logic block_rd_fifo_push;
logic clr_fiber_addr;
logic clr_final_pushed_done;
logic clr_pop_infifo_sticky;
logic clr_pushed_done_crd;
logic clr_pushed_done_seg;
logic clr_readout_loop_crd;
logic clr_readout_loop_seg;
logic clr_rep;
logic clr_req_made_crd;
logic clr_req_made_seg;
logic clr_req_rec_crd;
logic clr_req_rec_seg;
logic clr_seen_root_eos;
logic clr_used_data;
logic [16:0] coord_fifo_in_packed;
logic [16:0] coord_fifo_out_packed;
logic coordinate_fifo_empty;
logic coordinate_fifo_full;
logic coordinate_fifo_push;
logic [0:0][15:0] crd_ID_out_to_fifo;
logic [0:0][15:0] crd_addr_out_to_fifo;
logic crd_grant_push;
logic crd_in_done_state;
logic [0:0][15:0] crd_op_out_to_fifo;
logic [16:0] crd_out_to_fifo;
logic crd_pop_infifo;
logic crd_rd_rsp_fifo_pop;
logic crd_req_push;
logic [16:0] crd_res_fifo_data_in_0;
logic [16:0] crd_res_fifo_data_out;
logic [16:0] crd_res_fifo_fill_data_in;
logic crd_res_fifo_full;
logic crd_res_fifo_pop;
logic crd_res_fifo_push_alloc;
logic crd_res_fifo_push_alloc_0;
logic crd_res_fifo_push_fill;
logic crd_res_fifo_push_fill_0;
logic crd_res_fifo_push_reserve_0;
logic crd_res_fifo_valid;
logic crd_stop_lvl_geq;
logic done_in;
logic en_reg_data_in;
logic eos_in;
logic [15:0] fiber_addr;
logic [15:0] fiber_addr_pre;
logic [15:0] fiber_addr_pre_d1;
logic [15:0] fiber_addr_pre_d1_d1;
logic fifo_full;
logic [1:0] fifo_full_pre;
logic [16:0] fifo_out_us_packed;
logic fifo_us_full;
logic [16:0] fifo_us_in_packed;
logic final_pushed_done_sticky_sticky;
logic final_pushed_done_sticky_was_high;
logic gclk;
logic go_to_readout_sticky_sticky;
logic go_to_readout_sticky_was_high;
logic inc_fiber_addr;
logic inc_rep;
logic inc_req_made_crd;
logic inc_req_made_seg;
logic inc_req_rec_crd;
logic inc_req_rec_seg;
logic inc_requests_REC_CRD_READ;
logic inc_requests_made_CRDDD_READ;
logic infifo_eos_in;
logic [15:0] infifo_pos_in;
logic infifo_valid_in;
logic [0:0][16:0] input_fifo_data_out;
logic input_fifo_empty;
logic iter_finish_sticky;
logic iter_finish_was_high;
logic last_stop_done;
logic [16:0] last_stop_token;
logic last_valid_accepting;
logic maybe_in;
logic [15:0] next_seq_addr;
logic [15:0] next_seq_length;
logic no_outfifo_full;
logic [15:0] num_reps;
logic [15:0] num_req_made_crd;
logic [15:0] num_req_made_seg;
logic [15:0] num_req_rec_crd;
logic [15:0] num_req_rec_seg;
logic [0:0][16:0] op_out_fifo_data_in;
logic op_out_fifo_empty;
logic op_out_fifo_full;
logic op_out_fifo_push;
logic [0:0][15:0] op_out_to_fifo;
logic [15:0] payload_ptr;
logic pop_infifo;
logic pop_infifo_sticky_sticky;
logic pop_infifo_sticky_was_high;
logic [15:0] pos_addr;
logic pos_fifo_empty;
logic pos_fifo_full;
logic [16:0] pos_fifo_in_packed;
logic [16:0] pos_fifo_out_packed;
logic pos_out_fifo_push;
logic [16:0] pos_out_to_fifo;
logic [15:0] ptr_in;
logic [15:0] ptr_in_d1;
logic ptr_reg_en;
logic pushed_done_sticky_sticky;
logic pushed_done_sticky_was_high;
logic rd_rsp_fifo_empty;
logic rd_rsp_fifo_full;
logic [16:0] rd_rsp_fifo_out_data;
logic [16:0] rd_rsp_fifo_out_data_d1;
logic rd_rsp_fifo_valid;
logic readout_dst_crd;
logic readout_dst_seg;
logic readout_loop_sticky_sticky;
logic readout_loop_sticky_was_high;
logic rep_finish_sticky;
logic rep_finish_was_high;
logic [1:0] rr_arbiter_grant_out;
scan_seq_crd_state scan_seq_crd_current_state;
scan_seq_crd_state scan_seq_crd_next_state;
scan_seq_seg_state scan_seq_seg_current_state;
scan_seq_seg_state scan_seq_seg_next_state;
logic seen_root_eos_sticky;
logic seen_root_eos_was_high;
logic [0:0][15:0] seg_ID_out_to_fifo;
logic [0:0][15:0] seg_addr_out_to_fifo;
logic seg_grant_push;
logic seg_in_done_state;
logic seg_in_start_state;
logic [0:0][15:0] seg_op_out_to_fifo;
logic seg_pop_infifo;
logic seg_rd_rsp_fifo_pop;
logic seg_req_push;
logic [16:0] seg_res_fifo_data_out_0;
logic [16:0] seg_res_fifo_data_out_1;
logic seg_res_fifo_done_out;
logic [16:0] seg_res_fifo_fill_data_in;
logic seg_res_fifo_full;
logic seg_res_fifo_pop;
logic seg_res_fifo_pop_0;
logic seg_res_fifo_push_alloc;
logic seg_res_fifo_push_alloc_0;
logic seg_res_fifo_push_fill;
logic seg_res_fifo_push_fill_0;
logic seg_res_fifo_push_reserve_0;
logic seg_res_fifo_valid;
logic seg_stop_lvl_geq;
logic seg_stop_lvl_geq_p1;
logic [15:0] seq_addr;
logic [15:0] seq_length;
logic [15:0] seq_length_ptr_math;
logic set_final_pushed_done;
logic set_pushed_done_crd;
logic set_pushed_done_seg;
logic set_readout_loop_crd;
logic set_readout_loop_seg;
logic update_seq_state;
logic [15:0] us_fifo_inject_data;
logic us_fifo_inject_eos;
logic us_fifo_inject_push;
logic us_fifo_push;
logic use_data_sticky_sticky;
logic use_data_sticky_was_high;
logic [15:0] valid_cnt;
logic valid_inc;
logic valid_rst;
assign gclk = clk & tile_en;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    fiber_addr_pre <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      fiber_addr_pre <= 16'h0;
    end
    else if (clr_fiber_addr) begin
      fiber_addr_pre <= 16'h0;
    end
    else if (inc_fiber_addr) begin
      fiber_addr_pre <= fiber_addr_pre + 16'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_reps <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      num_reps <= 16'h0;
    end
    else if (clr_rep) begin
      num_reps <= 16'h0;
    end
    else if (inc_rep) begin
      num_reps <= num_reps + 16'h1;
    end
  end
end
assign us_fifo_push = root ? us_fifo_inject_push: us_pos_in_valid;
assign fifo_us_in_packed[16] = root ? us_fifo_inject_eos: us_pos_in[16];
assign fifo_us_in_packed[15:0] = root ? us_fifo_inject_data: us_pos_in[15:0];
assign infifo_eos_in = fifo_out_us_packed[16];
assign infifo_pos_in = fifo_out_us_packed[15:0];
assign pop_infifo = seg_pop_infifo | crd_pop_infifo;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    pop_infifo_sticky_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      pop_infifo_sticky_was_high <= 1'h0;
    end
    else if (clr_pop_infifo_sticky) begin
      pop_infifo_sticky_was_high <= 1'h0;
    end
    else if (pop_infifo) begin
      pop_infifo_sticky_was_high <= 1'h1;
    end
  end
end
assign pop_infifo_sticky_sticky = pop_infifo_sticky_was_high;
assign fifo_out_us_packed = input_fifo_data_out;
assign us_pos_in_ready = ~fifo_us_full;
assign infifo_valid_in = ~input_fifo_empty;
assign rd_rsp_data_in_ready = ~rd_rsp_fifo_full;
assign rd_rsp_fifo_valid = ~rd_rsp_fifo_empty;
assign base_rr = {crd_req_push, seg_req_push};
assign {crd_grant_push, seg_grant_push} = rr_arbiter_grant_out;
assign addr_out_to_fifo = crd_grant_push ? crd_addr_out_to_fifo: seg_addr_out_to_fifo;
assign op_out_to_fifo = crd_grant_push ? crd_op_out_to_fifo: seg_op_out_to_fifo;
assign ID_out_to_fifo = crd_grant_push ? crd_ID_out_to_fifo: seg_ID_out_to_fifo;
assign addr_out_fifo_push = seg_grant_push | crd_grant_push;
assign addr_out_fifo_data_in = {1'h0, addr_out_to_fifo};
assign addr_out_valid = ~addr_out_fifo_empty;
assign op_out_fifo_push = seg_grant_push | crd_grant_push;
assign op_out_fifo_data_in = {1'h0, op_out_to_fifo};
assign op_out_valid = ~op_out_fifo_empty;
assign ID_out_fifo_push = seg_grant_push | crd_grant_push;
assign ID_out_fifo_data_in = {1'h0, ID_out_to_fifo};
assign ID_out_valid = ~ID_out_fifo_empty;
assign no_outfifo_full = ~(ID_out_fifo_full | op_out_fifo_full | addr_out_fifo_full);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    pushed_done_sticky_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      pushed_done_sticky_was_high <= 1'h0;
    end
    else if (clr_pushed_done_seg | clr_pushed_done_crd) begin
      pushed_done_sticky_was_high <= 1'h0;
    end
    else if (set_pushed_done_seg | set_pushed_done_crd) begin
      pushed_done_sticky_was_high <= 1'h1;
    end
  end
end
assign pushed_done_sticky_sticky = pushed_done_sticky_was_high;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    readout_loop_sticky_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      readout_loop_sticky_was_high <= 1'h0;
    end
    else if (clr_readout_loop_seg | clr_readout_loop_crd) begin
      readout_loop_sticky_was_high <= 1'h0;
    end
    else if (set_readout_loop_seg | set_readout_loop_crd) begin
      readout_loop_sticky_was_high <= 1'h1;
    end
  end
end
assign readout_loop_sticky_sticky = readout_loop_sticky_was_high;
assign seg_res_fifo_push_alloc_0 = seg_res_fifo_push_alloc & (~lookup);
assign seg_res_fifo_push_reserve_0 = rd_rsp_fifo_valid & (rd_rsp_fifo_out_data[16] == 1'h0) & (~block_mode) &
    (~lookup);
assign seg_res_fifo_push_fill_0 = seg_res_fifo_push_fill & (~lookup);
assign seg_res_fifo_pop_0 = seg_res_fifo_pop & (~lookup);
assign crd_res_fifo_data_in_0 = {1'h0, rd_rsp_fifo_out_data[15:0]};
assign crd_res_fifo_fill_data_in = lookup ? seg_res_fifo_fill_data_in: dense ? crd_out_to_fifo:
    seg_res_fifo_data_out_0;
assign crd_res_fifo_push_alloc_0 = lookup ? seg_res_fifo_push_alloc: crd_res_fifo_push_alloc;
assign crd_res_fifo_push_reserve_0 = rd_rsp_fifo_valid & ((rd_rsp_fifo_out_data[16] == 1'h1) | block_mode | lookup);
assign crd_res_fifo_push_fill_0 = lookup ? seg_res_fifo_push_fill: crd_res_fifo_push_fill;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    last_stop_token <= 17'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      last_stop_token <= 17'h0;
    end
    else if (1'h0) begin
      last_stop_token <= 17'h0;
    end
    else if (seg_in_start_state ? 1'h0: seg_res_fifo_push_fill & seg_res_fifo_push_alloc & (lookup ? ~crd_res_fifo_full: ~seg_res_fifo_full) & seg_res_fifo_fill_data_in[16] & (seg_res_fifo_fill_data_in[9:8] == 2'h0)) begin
      last_stop_token <= seg_in_start_state ? input_fifo_data_out + 17'h1: seg_res_fifo_fill_data_in;
    end
  end
end
assign last_stop_done = last_stop_token[15:0] == (stop_lvl + 16'h2);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    use_data_sticky_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      use_data_sticky_was_high <= 1'h0;
    end
    else if (clr_used_data) begin
      use_data_sticky_was_high <= 1'h0;
    end
    else if (infifo_valid_in & (~infifo_eos_in)) begin
      use_data_sticky_was_high <= 1'h1;
    end
  end
end
assign use_data_sticky_sticky = use_data_sticky_was_high;
assign clr_used_data = readout_loop_sticky_sticky & spacc_mode;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    valid_cnt <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      valid_cnt <= 16'h0;
    end
    else if (valid_rst) begin
      valid_cnt <= 16'h0;
    end
    else if (valid_inc) begin
      valid_cnt <= valid_cnt + 16'h1;
    end
  end
end
assign ptr_in = rd_rsp_fifo_out_data[15:0];

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    ptr_in_d1 <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      ptr_in_d1 <= 16'h0;
    end
    else if (1'h0) begin
      ptr_in_d1 <= 16'h0;
    end
    else if (ptr_reg_en) begin
      ptr_in_d1 <= ptr_in;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    fiber_addr_pre_d1 <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      fiber_addr_pre_d1 <= 16'h0;
    end
    else if (1'h0) begin
      fiber_addr_pre_d1 <= 16'h0;
    end
    else if (1'h1) begin
      fiber_addr_pre_d1 <= fiber_addr_pre;
    end
  end
end
assign seq_length_ptr_math = seg_res_fifo_data_out_1 - seg_res_fifo_data_out_0[15:0];
assign pos_addr = root ? 16'h0: infifo_pos_in;
assign next_seq_addr = ptr_in_d1 + inner_dim_offset;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    seq_length <= 16'h0;
    seq_addr <= 16'h0;
    payload_ptr <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      seq_length <= 16'h0;
      seq_addr <= 16'h0;
      payload_ptr <= 16'h0;
    end
    else if (update_seq_state) begin
      seq_length <= next_seq_length;
      seq_addr <= next_seq_addr;
      payload_ptr <= ptr_in_d1;
    end
  end
end
assign fiber_addr = fiber_addr_pre + seq_addr;
assign fifo_full = |fifo_full_pre;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    iter_finish_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      iter_finish_was_high <= 1'h0;
    end
    else if (clr_fiber_addr) begin
      iter_finish_was_high <= 1'h0;
    end
    else if (last_valid_accepting) begin
      iter_finish_was_high <= 1'h1;
    end
  end
end
assign iter_finish_sticky = last_valid_accepting | iter_finish_was_high;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    rep_finish_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      rep_finish_was_high <= 1'h0;
    end
    else if (clr_rep) begin
      rep_finish_was_high <= 1'h0;
    end
    else if (((repeat_factor - 16'h1) == num_reps) & inc_rep) begin
      rep_finish_was_high <= 1'h1;
    end
  end
end
assign rep_finish_sticky = (((repeat_factor - 16'h1) == num_reps) & inc_rep) | rep_finish_was_high;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    seen_root_eos_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      seen_root_eos_was_high <= 1'h0;
    end
    else if (clr_seen_root_eos) begin
      seen_root_eos_was_high <= 1'h0;
    end
    else if (infifo_eos_in & (infifo_pos_in == 16'h0)) begin
      seen_root_eos_was_high <= 1'h1;
    end
  end
end
assign seen_root_eos_sticky = (infifo_eos_in & (infifo_pos_in == 16'h0)) | seen_root_eos_was_high;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    rd_rsp_fifo_out_data_d1 <= 17'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      rd_rsp_fifo_out_data_d1 <= 17'h0;
    end
    else if (1'h0) begin
      rd_rsp_fifo_out_data_d1 <= 17'h0;
    end
    else if (en_reg_data_in) begin
      rd_rsp_fifo_out_data_d1 <= rd_rsp_fifo_out_data;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    fiber_addr_pre_d1_d1 <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      fiber_addr_pre_d1_d1 <= 16'h0;
    end
    else if (1'h0) begin
      fiber_addr_pre_d1_d1 <= 16'h0;
    end
    else if (en_reg_data_in) begin
      fiber_addr_pre_d1_d1 <= fiber_addr_pre_d1;
    end
  end
end
assign done_in = infifo_eos_in & infifo_valid_in & (infifo_pos_in[9:8] == 2'h1);
assign eos_in = infifo_eos_in & infifo_valid_in & (infifo_pos_in[9:8] == 2'h0);
assign maybe_in = infifo_eos_in & infifo_valid_in & (infifo_pos_in[9:8] == 2'h2);
assign seg_stop_lvl_geq = seg_res_fifo_fill_data_in[16] & (seg_res_fifo_fill_data_in[9:8] == 2'h0) &
    (seg_res_fifo_fill_data_in[7:0] >= stop_lvl[7:0]);
assign seg_stop_lvl_geq_p1 = seg_res_fifo_fill_data_in[16] & (seg_res_fifo_fill_data_in[9:8] == 2'h0) &
    (seg_res_fifo_fill_data_in[7:0] >= (stop_lvl[7:0] + 8'h1));

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    go_to_readout_sticky_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      go_to_readout_sticky_was_high <= 1'h0;
    end
    else if (clr_readout_loop_seg) begin
      go_to_readout_sticky_was_high <= 1'h0;
    end
    else if (seg_stop_lvl_geq_p1 & seg_res_fifo_push_alloc & seg_res_fifo_push_fill) begin
      go_to_readout_sticky_was_high <= 1'h1;
    end
  end
end
assign go_to_readout_sticky_sticky = (seg_stop_lvl_geq_p1 & seg_res_fifo_push_alloc & seg_res_fifo_push_fill) |
    go_to_readout_sticky_was_high;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_req_made_seg <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      num_req_made_seg <= 16'h0;
    end
    else if (clr_req_made_seg) begin
      num_req_made_seg <= 16'h0;
    end
    else if (inc_req_made_seg) begin
      num_req_made_seg <= num_req_made_seg + 16'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_req_rec_seg <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      num_req_rec_seg <= 16'h0;
    end
    else if (clr_req_rec_seg) begin
      num_req_rec_seg <= 16'h0;
    end
    else if (inc_req_rec_seg) begin
      num_req_rec_seg <= num_req_rec_seg + 16'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_req_made_crd <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      num_req_made_crd <= 16'h0;
    end
    else if (clr_req_made_crd) begin
      num_req_made_crd <= 16'h0;
    end
    else if (inc_req_made_crd) begin
      num_req_made_crd <= num_req_made_crd + 16'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_req_rec_crd <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      num_req_rec_crd <= 16'h0;
    end
    else if (clr_req_rec_crd) begin
      num_req_rec_crd <= 16'h0;
    end
    else if (inc_req_rec_crd) begin
      num_req_rec_crd <= num_req_rec_crd + 16'h1;
    end
  end
end
assign seg_res_fifo_done_out = seg_res_fifo_valid & seg_res_fifo_data_out_0[16] & (seg_res_fifo_data_out_0[9:8]
    == 2'h1);
assign crd_stop_lvl_geq = seg_res_fifo_valid & seg_res_fifo_data_out_0[16] & (seg_res_fifo_data_out_0[9:8]
    == 2'h0) & (seg_res_fifo_data_out_0[7:0] >= stop_lvl[7:0]);
assign readout_dst_crd = readout_loop_sticky_sticky;
assign readout_dst_seg = readout_loop_sticky_sticky;
assign inc_requests_made_CRDDD_READ = crd_grant_push;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    READS_MADE <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      READS_MADE <= 16'h0;
    end
    else if (inc_requests_made_CRDDD_READ) begin
      READS_MADE <= READS_MADE + 16'h1;
    end
  end
end
assign inc_requests_REC_CRD_READ = rd_rsp_fifo_valid & (rd_rsp_fifo_out_data[16] == 1'h1);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    READS_REC_CRD_READ <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      READS_REC_CRD_READ <= 16'h0;
    end
    else if (inc_requests_REC_CRD_READ) begin
      READS_REC_CRD_READ <= READS_REC_CRD_READ + 16'h1;
    end
  end
end
assign coord_fifo_in_packed = crd_res_fifo_data_out;
assign coord_out[16] = coord_fifo_out_packed[16];
assign coord_out[15:0] = coord_fifo_out_packed[15:0];

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    final_pushed_done_sticky_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      final_pushed_done_sticky_was_high <= 1'h0;
    end
    else if (clr_final_pushed_done) begin
      final_pushed_done_sticky_was_high <= 1'h0;
    end
    else if (set_final_pushed_done) begin
      final_pushed_done_sticky_was_high <= 1'h1;
    end
  end
end
assign final_pushed_done_sticky_sticky = final_pushed_done_sticky_was_high;
assign set_final_pushed_done = crd_res_fifo_valid & (~block_mode) & crd_res_fifo_data_out[16] &
    crd_res_fifo_valid & (crd_res_fifo_data_out[9:8] == 2'h3) & spacc_mode &
    crd_res_fifo_data_out[0];
assign clr_final_pushed_done = crd_res_fifo_valid & (~block_mode) & crd_res_fifo_data_out[16] &
    crd_res_fifo_valid & (crd_res_fifo_data_out[9:8] == 2'h3) & spacc_mode &
    (~crd_res_fifo_data_out[0]);
assign coordinate_fifo_push = crd_res_fifo_valid & (~block_mode) & (~(spacc_mode &
    final_pushed_done_sticky_sticky)) & (~(crd_res_fifo_data_out[16] &
    crd_res_fifo_valid & (crd_res_fifo_data_out[9:8] == 2'h3)));
assign coord_out_valid = ~coordinate_fifo_empty;
assign fifo_full_pre[0] = coordinate_fifo_full;
assign crd_res_fifo_pop = block_mode ? ~block_rd_fifo_full: spacc_mode ? (crd_res_fifo_data_out[16] &
    crd_res_fifo_valid & (crd_res_fifo_data_out[9:8] == 2'h3)) ? 1'h1:
    final_pushed_done_sticky_sticky ? ~block_rd_fifo_full: ~coordinate_fifo_full:
    ~coordinate_fifo_full;
assign pos_fifo_in_packed = pos_out_to_fifo;
assign pos_out[16] = pos_fifo_out_packed[16];
assign pos_out[15:0] = pos_fifo_out_packed[15:0];
assign pos_out_valid = ~pos_fifo_empty;
assign fifo_full_pre[1] = pos_fifo_full;
assign block_rd_fifo_push = crd_res_fifo_valid & (block_mode | (spacc_mode &
    final_pushed_done_sticky_sticky)) & (~(crd_res_fifo_data_out[16] &
    crd_res_fifo_valid & (crd_res_fifo_data_out[9:8] == 2'h3)));
assign block_rd_out_valid = ~block_rd_fifo_empty;

always_ff @(posedge clk, negedge rst_n) begin
  if (!rst_n) begin
    scan_seq_crd_current_state <= START_CRD;
  end
  else if (clk_en) begin
    if (flush) begin
      scan_seq_crd_current_state <= START_CRD;
    end
    else scan_seq_crd_current_state <= scan_seq_crd_next_state;
  end
end
always_comb begin
  scan_seq_crd_next_state = scan_seq_crd_current_state;
  unique case (scan_seq_crd_current_state)
    BLOCK_1_RD: begin
        if ((num_req_rec_crd == ptr_in_d1) & (~lookup)) begin
          scan_seq_crd_next_state = BLOCK_2_SIZE_REQ;
        end
        else if ((num_req_rec_crd == ptr_in_d1) & lookup) begin
          scan_seq_crd_next_state = FREE_CRD;
        end
        else scan_seq_crd_next_state = BLOCK_1_RD;
      end
    BLOCK_1_SIZE_REC: begin
        if (rd_rsp_fifo_valid) begin
          scan_seq_crd_next_state = BLOCK_1_RD;
        end
        else scan_seq_crd_next_state = BLOCK_1_SIZE_REC;
      end
    BLOCK_1_SIZE_REQ: begin
        if (crd_grant_push) begin
          scan_seq_crd_next_state = BLOCK_1_SIZE_REC;
        end
        else scan_seq_crd_next_state = BLOCK_1_SIZE_REQ;
      end
    BLOCK_2_RD: begin
        if (num_req_rec_crd == ptr_in_d1) begin
          scan_seq_crd_next_state = FREE_CRD;
        end
        else scan_seq_crd_next_state = BLOCK_2_RD;
      end
    BLOCK_2_SIZE_REC: begin
        if (rd_rsp_fifo_valid) begin
          scan_seq_crd_next_state = BLOCK_2_RD;
        end
        else scan_seq_crd_next_state = BLOCK_2_SIZE_REC;
      end
    BLOCK_2_SIZE_REQ: begin
        if (crd_grant_push) begin
          scan_seq_crd_next_state = BLOCK_2_SIZE_REC;
        end
        else scan_seq_crd_next_state = BLOCK_2_SIZE_REQ;
      end
    DENSE_STRM: scan_seq_crd_next_state = DENSE_STRM;
    DONE_CRD: begin
        if ((~spacc_mode) | (spacc_mode & seg_in_done_state)) begin
          scan_seq_crd_next_state = START_CRD;
        end
      end
    FREE_CRD: begin
        if (crd_grant_push & block_mode & (~lookup)) begin
          scan_seq_crd_next_state = FREE_CRD2;
        end
        else if (crd_grant_push & pushed_done_sticky_sticky & spacc_mode) begin
          scan_seq_crd_next_state = PASS_DONE_CRD;
        end
        else if (crd_grant_push & ((~spacc_mode) | (~pushed_done_sticky_sticky))) begin
          scan_seq_crd_next_state = DONE_CRD;
        end
        else scan_seq_crd_next_state = FREE_CRD;
      end
    FREE_CRD2: begin
        if (crd_grant_push) begin
          scan_seq_crd_next_state = DONE_CRD;
        end
        else scan_seq_crd_next_state = FREE_CRD2;
      end
    PASS_DONE_CRD: begin
        if ((~crd_res_fifo_full) & (~pos_fifo_full)) begin
          scan_seq_crd_next_state = DONE_CRD;
        end
      end
    READOUT_SYNC_LOCK: scan_seq_crd_next_state = DONE_CRD;
    SEQ_STRM: begin
        if ((seg_res_fifo_done_out | (spacc_mode & crd_stop_lvl_geq)) & (~crd_res_fifo_full) & (~pos_fifo_full)) begin
          scan_seq_crd_next_state = FREE_CRD;
        end
      end
    START_CRD: begin
        if (block_mode & tile_en) begin
          scan_seq_crd_next_state = BLOCK_1_SIZE_REQ;
        end
        else if (dense & (~lookup) & tile_en) begin
          scan_seq_crd_next_state = DENSE_STRM;
        end
        else if ((~dense) & (~lookup) & tile_en) begin
          scan_seq_crd_next_state = SEQ_STRM;
        end
      end
    default: scan_seq_crd_next_state = scan_seq_crd_current_state;
  endcase
end
always_comb begin
  unique case (scan_seq_crd_current_state)
    BLOCK_1_RD: begin :scan_seq_crd_BLOCK_1_RD_Output
        crd_addr_out_to_fifo = num_req_made_crd;
        crd_op_out_to_fifo = 16'h1;
        crd_ID_out_to_fifo = 16'h0;
        crd_req_push = (num_req_made_crd < ptr_in_d1) & (~crd_res_fifo_full);
        crd_rd_rsp_fifo_pop = num_req_rec_crd < ptr_in_d1;
        pos_out_fifo_push = 1'h0;
        crd_pop_infifo = 1'h0;
        en_reg_data_in = 1'h0;
        pos_out_to_fifo = 17'h0;
        crd_out_to_fifo = 17'h0;
        inc_req_made_crd = (num_req_made_crd < ptr_in_d1) & crd_grant_push & (~crd_res_fifo_full);
        clr_req_made_crd = 1'h0;
        inc_req_rec_crd = (num_req_rec_crd < ptr_in_d1) & rd_rsp_fifo_valid;
        clr_req_rec_crd = 1'h0;
        crd_res_fifo_push_alloc = (num_req_made_crd < ptr_in_d1) & crd_grant_push & (~crd_res_fifo_full);
        crd_res_fifo_push_fill = 1'h0;
        ptr_reg_en = 1'h0;
        seg_res_fifo_pop = 1'h0;
        clr_readout_loop_crd = 1'h0;
        set_readout_loop_crd = 1'h0;
        crd_in_done_state = 1'h0;
        set_pushed_done_crd = 1'h0;
        clr_pushed_done_crd = 1'h0;
      end :scan_seq_crd_BLOCK_1_RD_Output
    BLOCK_1_SIZE_REC: begin :scan_seq_crd_BLOCK_1_SIZE_REC_Output
        crd_addr_out_to_fifo = 16'h0;
        crd_op_out_to_fifo = 16'h0;
        crd_ID_out_to_fifo = 16'h0;
        crd_req_push = 1'h0;
        crd_rd_rsp_fifo_pop = 1'h1;
        pos_out_fifo_push = 1'h0;
        crd_pop_infifo = 1'h0;
        en_reg_data_in = 1'h0;
        pos_out_to_fifo = 17'h0;
        crd_out_to_fifo = 17'h0;
        inc_req_made_crd = 1'h0;
        clr_req_made_crd = 1'h1;
        inc_req_rec_crd = 1'h0;
        clr_req_rec_crd = 1'h0;
        crd_res_fifo_push_alloc = 1'h0;
        crd_res_fifo_push_fill = 1'h0;
        ptr_reg_en = rd_rsp_fifo_valid;
        seg_res_fifo_pop = 1'h0;
        clr_readout_loop_crd = 1'h0;
        set_readout_loop_crd = 1'h0;
        crd_in_done_state = 1'h0;
        set_pushed_done_crd = 1'h0;
        clr_pushed_done_crd = 1'h0;
      end :scan_seq_crd_BLOCK_1_SIZE_REC_Output
    BLOCK_1_SIZE_REQ: begin :scan_seq_crd_BLOCK_1_SIZE_REQ_Output
        crd_addr_out_to_fifo = 16'h0;
        crd_op_out_to_fifo = 16'h2;
        crd_ID_out_to_fifo = 16'h0;
        crd_req_push = ~crd_res_fifo_full;
        crd_rd_rsp_fifo_pop = 1'h0;
        pos_out_fifo_push = 1'h0;
        crd_pop_infifo = 1'h0;
        en_reg_data_in = 1'h0;
        pos_out_to_fifo = 17'h0;
        crd_out_to_fifo = 17'h0;
        inc_req_made_crd = 1'h0;
        clr_req_made_crd = 1'h0;
        inc_req_rec_crd = 1'h0;
        clr_req_rec_crd = 1'h0;
        crd_res_fifo_push_alloc = (~crd_res_fifo_full) & crd_grant_push;
        crd_res_fifo_push_fill = 1'h0;
        ptr_reg_en = 1'h0;
        seg_res_fifo_pop = 1'h0;
        clr_readout_loop_crd = 1'h0;
        set_readout_loop_crd = 1'h0;
        crd_in_done_state = 1'h0;
        set_pushed_done_crd = 1'h0;
        clr_pushed_done_crd = 1'h0;
      end :scan_seq_crd_BLOCK_1_SIZE_REQ_Output
    BLOCK_2_RD: begin :scan_seq_crd_BLOCK_2_RD_Output
        crd_addr_out_to_fifo = num_req_made_crd;
        crd_op_out_to_fifo = 16'h1;
        crd_ID_out_to_fifo = 16'h1;
        crd_req_push = (num_req_made_crd < ptr_in_d1) & (~crd_res_fifo_full);
        crd_rd_rsp_fifo_pop = num_req_rec_crd < ptr_in_d1;
        pos_out_fifo_push = 1'h0;
        crd_pop_infifo = 1'h0;
        en_reg_data_in = 1'h0;
        pos_out_to_fifo = 17'h0;
        crd_out_to_fifo = 17'h0;
        inc_req_made_crd = (num_req_made_crd < ptr_in_d1) & crd_grant_push & (~crd_res_fifo_full);
        clr_req_made_crd = 1'h0;
        inc_req_rec_crd = (num_req_rec_crd < ptr_in_d1) & rd_rsp_fifo_valid;
        clr_req_rec_crd = 1'h0;
        crd_res_fifo_push_alloc = (num_req_made_crd < ptr_in_d1) & crd_grant_push & (~crd_res_fifo_full);
        crd_res_fifo_push_fill = 1'h0;
        ptr_reg_en = 1'h0;
        seg_res_fifo_pop = 1'h0;
        clr_readout_loop_crd = 1'h0;
        set_readout_loop_crd = 1'h0;
        crd_in_done_state = 1'h0;
        set_pushed_done_crd = 1'h0;
        clr_pushed_done_crd = 1'h0;
      end :scan_seq_crd_BLOCK_2_RD_Output
    BLOCK_2_SIZE_REC: begin :scan_seq_crd_BLOCK_2_SIZE_REC_Output
        crd_addr_out_to_fifo = 16'h0;
        crd_op_out_to_fifo = 16'h0;
        crd_ID_out_to_fifo = 16'h0;
        crd_req_push = 1'h0;
        crd_rd_rsp_fifo_pop = 1'h1;
        pos_out_fifo_push = 1'h0;
        crd_pop_infifo = 1'h0;
        en_reg_data_in = 1'h0;
        pos_out_to_fifo = 17'h0;
        crd_out_to_fifo = 17'h0;
        inc_req_made_crd = 1'h0;
        clr_req_made_crd = 1'h1;
        inc_req_rec_crd = 1'h0;
        clr_req_rec_crd = 1'h1;
        crd_res_fifo_push_alloc = 1'h0;
        crd_res_fifo_push_fill = 1'h0;
        ptr_reg_en = rd_rsp_fifo_valid;
        seg_res_fifo_pop = 1'h0;
        clr_readout_loop_crd = 1'h0;
        set_readout_loop_crd = 1'h0;
        crd_in_done_state = 1'h0;
        set_pushed_done_crd = 1'h0;
        clr_pushed_done_crd = 1'h0;
      end :scan_seq_crd_BLOCK_2_SIZE_REC_Output
    BLOCK_2_SIZE_REQ: begin :scan_seq_crd_BLOCK_2_SIZE_REQ_Output
        crd_addr_out_to_fifo = 16'h0;
        crd_op_out_to_fifo = 16'h2;
        crd_ID_out_to_fifo = 16'h1;
        crd_req_push = ~crd_res_fifo_full;
        crd_rd_rsp_fifo_pop = 1'h0;
        pos_out_fifo_push = 1'h0;
        crd_pop_infifo = 1'h0;
        en_reg_data_in = 1'h0;
        pos_out_to_fifo = 17'h0;
        crd_out_to_fifo = 17'h0;
        inc_req_made_crd = 1'h0;
        clr_req_made_crd = 1'h0;
        inc_req_rec_crd = 1'h0;
        clr_req_rec_crd = 1'h0;
        crd_res_fifo_push_alloc = (~crd_res_fifo_full) & crd_grant_push;
        crd_res_fifo_push_fill = 1'h0;
        ptr_reg_en = 1'h0;
        seg_res_fifo_pop = 1'h0;
        clr_readout_loop_crd = 1'h0;
        set_readout_loop_crd = 1'h0;
        crd_in_done_state = 1'h0;
        set_pushed_done_crd = 1'h0;
        clr_pushed_done_crd = 1'h0;
      end :scan_seq_crd_BLOCK_2_SIZE_REQ_Output
    DENSE_STRM: begin :scan_seq_crd_DENSE_STRM_Output
        crd_addr_out_to_fifo = 16'h0;
        crd_op_out_to_fifo = 16'h0;
        crd_ID_out_to_fifo = 16'h0;
        crd_req_push = 1'h0;
        crd_rd_rsp_fifo_pop = 1'h0;
        pos_out_fifo_push = seg_res_fifo_valid & (~pos_fifo_full) & (~crd_res_fifo_full) &
            (seg_res_fifo_data_out_0[16] ? 1'h1: dim_size > num_req_made_crd);
        crd_pop_infifo = 1'h0;
        en_reg_data_in = 1'h0;
        pos_out_to_fifo = seg_res_fifo_data_out_0[16] ? seg_res_fifo_data_out_0:
            17'((seg_res_fifo_data_out_0[15:0] * dim_size) + num_req_made_crd);
        crd_out_to_fifo = seg_res_fifo_data_out_0[16] ? seg_res_fifo_data_out_0: 17'(num_req_made_crd);
        inc_req_made_crd = seg_res_fifo_valid & (dim_size > num_req_made_crd) &
            (~seg_res_fifo_data_out_0[16]) & (~pos_fifo_full) & (~crd_res_fifo_full);
        clr_req_made_crd = seg_res_fifo_valid & seg_res_fifo_data_out_0[16];
        inc_req_rec_crd = 1'h0;
        clr_req_rec_crd = 1'h0;
        crd_res_fifo_push_alloc = seg_res_fifo_valid & (~pos_fifo_full) & (~crd_res_fifo_full) &
            (seg_res_fifo_data_out_0[16] ? 1'h1: dim_size > num_req_made_crd);
        crd_res_fifo_push_fill = seg_res_fifo_valid & (~pos_fifo_full) & (~crd_res_fifo_full) &
            (seg_res_fifo_data_out_0[16] ? 1'h1: dim_size > num_req_made_crd);
        ptr_reg_en = 1'h0;
        seg_res_fifo_pop = seg_res_fifo_valid & (~pos_fifo_full) & (~crd_res_fifo_full) &
            (seg_res_fifo_data_out_0[16] ? 1'h1: ((dim_size - 16'h1) == num_req_made_crd) &
            inc_req_made_crd);
        clr_readout_loop_crd = 1'h0;
        set_readout_loop_crd = 1'h0;
        crd_in_done_state = 1'h0;
        set_pushed_done_crd = 1'h0;
        clr_pushed_done_crd = 1'h0;
      end :scan_seq_crd_DENSE_STRM_Output
    DONE_CRD: begin :scan_seq_crd_DONE_CRD_Output
        crd_addr_out_to_fifo = 16'h0;
        crd_op_out_to_fifo = 16'h0;
        crd_ID_out_to_fifo = 16'h0;
        crd_req_push = 1'h0;
        crd_rd_rsp_fifo_pop = 1'h0;
        pos_out_fifo_push = 1'h0;
        crd_pop_infifo = 1'h0;
        en_reg_data_in = 1'h0;
        pos_out_to_fifo = 17'h0;
        crd_out_to_fifo = 17'h0;
        inc_req_made_crd = 1'h0;
        clr_req_made_crd = 1'h1;
        inc_req_rec_crd = 1'h0;
        clr_req_rec_crd = 1'h1;
        crd_res_fifo_push_alloc = 1'h0;
        crd_res_fifo_push_fill = 1'h0;
        ptr_reg_en = 1'h0;
        seg_res_fifo_pop = 1'h0;
        crd_in_done_state = 1'h1;
        set_readout_loop_crd = 1'h0;
        clr_readout_loop_crd = 1'h0;
        set_pushed_done_crd = 1'h0;
        clr_pushed_done_crd = 1'h0;
      end :scan_seq_crd_DONE_CRD_Output
    FREE_CRD: begin :scan_seq_crd_FREE_CRD_Output
        crd_addr_out_to_fifo = 16'h0;
        crd_op_out_to_fifo = 16'h0;
        crd_ID_out_to_fifo = block_mode ? 16'h0: 16'h1;
        crd_req_push = 1'h1;
        crd_rd_rsp_fifo_pop = 1'h0;
        pos_out_fifo_push = 1'h0;
        crd_pop_infifo = 1'h0;
        en_reg_data_in = 1'h0;
        pos_out_to_fifo = 17'h0;
        crd_out_to_fifo = 17'h0;
        inc_req_made_crd = 1'h0;
        clr_req_made_crd = 1'h1;
        inc_req_rec_crd = 1'h0;
        clr_req_rec_crd = 1'h1;
        crd_res_fifo_push_alloc = 1'h0;
        crd_res_fifo_push_fill = 1'h0;
        ptr_reg_en = 1'h0;
        seg_res_fifo_pop = 1'h0;
        clr_readout_loop_crd = 1'h0;
        set_readout_loop_crd = 1'h0;
        crd_in_done_state = 1'h0;
        set_pushed_done_crd = 1'h0;
        clr_pushed_done_crd = 1'h0;
      end :scan_seq_crd_FREE_CRD_Output
    FREE_CRD2: begin :scan_seq_crd_FREE_CRD2_Output
        crd_addr_out_to_fifo = 16'h0;
        crd_op_out_to_fifo = 16'h0;
        crd_ID_out_to_fifo = 16'h1;
        crd_req_push = 1'h1;
        crd_rd_rsp_fifo_pop = 1'h0;
        pos_out_fifo_push = 1'h0;
        crd_pop_infifo = 1'h0;
        en_reg_data_in = 1'h0;
        pos_out_to_fifo = 17'h0;
        crd_out_to_fifo = 17'h0;
        inc_req_made_crd = 1'h0;
        clr_req_made_crd = 1'h1;
        inc_req_rec_crd = 1'h0;
        clr_req_rec_crd = 1'h1;
        crd_res_fifo_push_alloc = 1'h0;
        crd_res_fifo_push_fill = 1'h0;
        ptr_reg_en = 1'h0;
        seg_res_fifo_pop = 1'h0;
        clr_readout_loop_crd = 1'h0;
        set_readout_loop_crd = 1'h0;
        crd_in_done_state = 1'h0;
        set_pushed_done_crd = 1'h0;
        clr_pushed_done_crd = 1'h0;
      end :scan_seq_crd_FREE_CRD2_Output
    PASS_DONE_CRD: begin :scan_seq_crd_PASS_DONE_CRD_Output
        crd_addr_out_to_fifo = 16'h0;
        crd_op_out_to_fifo = 16'h0;
        crd_ID_out_to_fifo = 16'h0;
        crd_req_push = 1'h0;
        crd_rd_rsp_fifo_pop = 1'h0;
        pos_out_fifo_push = (~pos_fifo_full) & (~crd_res_fifo_full) & seg_res_fifo_done_out &
            seg_res_fifo_valid;
        crd_pop_infifo = 1'h0;
        en_reg_data_in = 1'h0;
        pos_out_to_fifo = {1'h1, 6'h0, 2'h1, 8'h0};
        crd_out_to_fifo = 17'h0;
        inc_req_made_crd = 1'h0;
        clr_req_made_crd = 1'h0;
        inc_req_rec_crd = 1'h0;
        clr_req_rec_crd = 1'h0;
        crd_res_fifo_push_alloc = (~pos_fifo_full) & (~crd_res_fifo_full) & seg_res_fifo_done_out &
            seg_res_fifo_valid;
        crd_res_fifo_push_fill = (~pos_fifo_full) & (~crd_res_fifo_full) & seg_res_fifo_done_out &
            seg_res_fifo_valid;
        ptr_reg_en = 1'h0;
        seg_res_fifo_pop = (~pos_fifo_full) & (~crd_res_fifo_full) & seg_res_fifo_done_out &
            seg_res_fifo_valid;
        clr_pushed_done_crd = 1'h0;
        clr_readout_loop_crd = 1'h0;
        set_readout_loop_crd = 1'h0;
        crd_in_done_state = 1'h0;
        set_pushed_done_crd = 1'h0;
      end :scan_seq_crd_PASS_DONE_CRD_Output
    READOUT_SYNC_LOCK: begin :scan_seq_crd_READOUT_SYNC_LOCK_Output
        crd_addr_out_to_fifo = 16'h0;
        crd_op_out_to_fifo = 16'h0;
        crd_ID_out_to_fifo = 16'h0;
        crd_req_push = 1'h0;
        crd_rd_rsp_fifo_pop = 1'h0;
        pos_out_fifo_push = 1'h0;
        crd_pop_infifo = 1'h0;
        en_reg_data_in = 1'h0;
        pos_out_to_fifo = 17'h0;
        crd_out_to_fifo = 17'h0;
        inc_req_made_crd = 1'h0;
        clr_req_made_crd = 1'h0;
        inc_req_rec_crd = 1'h0;
        clr_req_rec_crd = 1'h0;
        crd_res_fifo_push_alloc = 1'h0;
        crd_res_fifo_push_fill = 1'h0;
        ptr_reg_en = 1'h0;
        seg_res_fifo_pop = 1'h0;
        clr_pushed_done_crd = 1'h1;
        clr_readout_loop_crd = 1'h1;
        set_readout_loop_crd = 1'h0;
        crd_in_done_state = 1'h0;
        set_pushed_done_crd = 1'h0;
      end :scan_seq_crd_READOUT_SYNC_LOCK_Output
    SEQ_STRM: begin :scan_seq_crd_SEQ_STRM_Output
        crd_addr_out_to_fifo = num_req_made_crd + seg_res_fifo_data_out_0[15:0];
        crd_op_out_to_fifo = 16'h1;
        crd_ID_out_to_fifo = 16'h1;
        crd_req_push = seg_res_fifo_valid & (~seg_res_fifo_data_out_0[16]) & (~crd_res_fifo_full) &
            (num_req_made_crd < seq_length_ptr_math) & (~pos_fifo_full);
        crd_rd_rsp_fifo_pop = 1'h1;
        pos_out_fifo_push = seg_res_fifo_data_out_0[16] ? (~pos_fifo_full) & (~crd_res_fifo_full) &
            seg_res_fifo_valid: crd_grant_push & (num_req_made_crd < seq_length_ptr_math) &
            (~pos_fifo_full) & (~crd_res_fifo_full) & seg_res_fifo_valid;
        crd_pop_infifo = 1'h0;
        en_reg_data_in = 1'h0;
        pos_out_to_fifo = seg_res_fifo_data_out_0[16] ? seg_res_fifo_data_out_0: {1'h0, num_req_made_crd +
            seg_res_fifo_data_out_0[15:0]};
        crd_out_to_fifo = 17'h0;
        inc_req_made_crd = crd_grant_push & (num_req_made_crd < seq_length_ptr_math) & (~pos_fifo_full) &
            (~crd_res_fifo_full) & seg_res_fifo_valid;
        clr_req_made_crd = ((crd_grant_push & ((seq_length_ptr_math - 16'h1) == num_req_made_crd)) |
            (seq_length_ptr_math == 16'h0)) & (~pos_fifo_full) & (~crd_res_fifo_full) &
            seg_res_fifo_valid;
        inc_req_rec_crd = 1'h0;
        clr_req_rec_crd = 1'h0;
        crd_res_fifo_push_alloc = seg_res_fifo_data_out_0[16] ? (~pos_fifo_full) & (~crd_res_fifo_full) &
            seg_res_fifo_valid: crd_grant_push & (num_req_made_crd < seq_length_ptr_math) &
            (~pos_fifo_full) & (~crd_res_fifo_full) & seg_res_fifo_valid;
        crd_res_fifo_push_fill = seg_res_fifo_valid & seg_res_fifo_data_out_0[16] & (~pos_fifo_full) &
            (~crd_res_fifo_full);
        ptr_reg_en = 1'h0;
        seg_res_fifo_pop = clr_req_made_crd | (seg_res_fifo_valid & seg_res_fifo_data_out_0[16] &
            (~pos_fifo_full) & (~crd_res_fifo_full));
        clr_readout_loop_crd = 1'h0;
        set_readout_loop_crd = 1'h0;
        crd_in_done_state = 1'h0;
        set_pushed_done_crd = 1'h0;
        clr_pushed_done_crd = 1'h0;
      end :scan_seq_crd_SEQ_STRM_Output
    START_CRD: begin :scan_seq_crd_START_CRD_Output
        crd_addr_out_to_fifo = 16'h0;
        crd_op_out_to_fifo = 16'h0;
        crd_ID_out_to_fifo = 16'h0;
        crd_req_push = 1'h0;
        crd_rd_rsp_fifo_pop = 1'h0;
        pos_out_fifo_push = 1'h0;
        crd_pop_infifo = 1'h0;
        en_reg_data_in = 1'h0;
        pos_out_to_fifo = 17'h0;
        crd_out_to_fifo = 17'h0;
        inc_req_made_crd = 1'h0;
        clr_req_made_crd = 1'h0;
        inc_req_rec_crd = 1'h0;
        clr_req_rec_crd = 1'h0;
        crd_res_fifo_push_alloc = 1'h0;
        crd_res_fifo_push_fill = 1'h0;
        ptr_reg_en = 1'h0;
        seg_res_fifo_pop = 1'h0;
        clr_readout_loop_crd = 1'h0;
        set_readout_loop_crd = 1'h0;
        crd_in_done_state = 1'h0;
        set_pushed_done_crd = 1'h0;
        clr_pushed_done_crd = 1'h0;
      end :scan_seq_crd_START_CRD_Output
    default: begin :scan_seq_crd_default_Output
        crd_addr_out_to_fifo = 16'h0;
        crd_op_out_to_fifo = 16'h0;
        crd_ID_out_to_fifo = 16'h0;
        crd_req_push = 1'h0;
        crd_rd_rsp_fifo_pop = 1'h0;
        pos_out_fifo_push = 1'h0;
        crd_pop_infifo = 1'h0;
        en_reg_data_in = 1'h0;
        pos_out_to_fifo = 17'h0;
        crd_out_to_fifo = 17'h0;
        inc_req_made_crd = 1'h0;
        clr_req_made_crd = 1'h0;
        inc_req_rec_crd = 1'h0;
        clr_req_rec_crd = 1'h0;
        crd_res_fifo_push_alloc = 1'h0;
        crd_res_fifo_push_fill = 1'h0;
        ptr_reg_en = 1'h0;
        seg_res_fifo_pop = 1'h0;
        clr_readout_loop_crd = 1'h0;
        set_readout_loop_crd = 1'h0;
        crd_in_done_state = 1'h0;
        set_pushed_done_crd = 1'h0;
        clr_pushed_done_crd = 1'h0;
      end :scan_seq_crd_default_Output
  endcase
end

always_ff @(posedge clk, negedge rst_n) begin
  if (!rst_n) begin
    scan_seq_seg_current_state <= START_SEG;
  end
  else if (clk_en) begin
    if (flush) begin
      scan_seq_seg_current_state <= START_SEG;
    end
    else scan_seq_seg_current_state <= scan_seq_seg_next_state;
  end
end
always_comb begin
  scan_seq_seg_next_state = scan_seq_seg_current_state;
  unique case (scan_seq_seg_current_state)
    DONE_SEG: begin
        if (lookup ? 1'h1: (~dense) & crd_in_done_state) begin
          scan_seq_seg_next_state = START_SEG;
        end
      end
    FREE_SEG: begin
        if (seg_grant_push) begin
          scan_seq_seg_next_state = DONE_SEG;
        end
      end
    INJECT_0: scan_seq_seg_next_state = INJECT_DONE;
    INJECT_DONE: scan_seq_seg_next_state = READ;
    INJECT_ROUTING: begin
        if (~seg_res_fifo_full) begin
          scan_seq_seg_next_state = READ;
        end
      end
    LOOKUP: begin
        if (((done_in & (~spacc_mode)) | (spacc_mode & seg_stop_lvl_geq & infifo_valid_in & (~pushed_done_sticky_sticky))) & (~crd_res_fifo_full)) begin
          scan_seq_seg_next_state = FREE_SEG;
        end
        else scan_seq_seg_next_state = LOOKUP;
      end
    PASS_DONE_SEG: begin
        if ((readout_loop_sticky_sticky & ((~pushed_done_sticky_sticky) | (~seg_res_fifo_full))) | (~last_stop_done) | (~seg_res_fifo_full)) begin
          scan_seq_seg_next_state = FREE_SEG;
        end
      end
    PASS_STOP_SEG: begin
        if (((infifo_valid_in & (~lookup) & spacc_mode & seg_stop_lvl_geq) | readout_loop_sticky_sticky) & (~seg_res_fifo_full)) begin
          scan_seq_seg_next_state = PASS_DONE_SEG;
        end
        else if (infifo_valid_in & (~lookup) & (~seg_res_fifo_full)) begin
          scan_seq_seg_next_state = READ;
        end
        else scan_seq_seg_next_state = PASS_STOP_SEG;
      end
    READ: begin
        if (maybe_in | (dense & (~done_in) & (~seg_res_fifo_full) & infifo_valid_in) | (((~spacc_mode) | (~readout_loop_sticky_sticky)) & (~dense) & eos_in & ((~spacc_mode) | (~use_data_sticky_sticky)))) begin
          scan_seq_seg_next_state = PASS_STOP_SEG;
        end
        else if (seg_grant_push & (~seg_res_fifo_full)) begin
          scan_seq_seg_next_state = READ_ALT;
        end
        else if (done_in & (~seg_res_fifo_full)) begin
          scan_seq_seg_next_state = FREE_SEG;
        end
        else scan_seq_seg_next_state = READ;
      end
    READ_ALT: begin
        if (seg_grant_push & (~seg_res_fifo_full)) begin
          scan_seq_seg_next_state = PASS_STOP_SEG;
        end
        else scan_seq_seg_next_state = READ_ALT;
      end
    START_SEG: begin
        if (block_mode) begin
          scan_seq_seg_next_state = START_SEG;
        end
        else if ((~root) & (~lookup) & (~block_mode) & (~spacc_mode) & tile_en) begin
          scan_seq_seg_next_state = READ;
        end
        else if ((~root) & (~lookup) & (~block_mode) & (infifo_valid_in | readout_loop_sticky_sticky) & spacc_mode & tile_en) begin
          scan_seq_seg_next_state = INJECT_ROUTING;
        end
        else if (root & (~lookup) & (~block_mode) & tile_en) begin
          scan_seq_seg_next_state = INJECT_0;
        end
        else if ((~root) & lookup & (~block_mode) & tile_en) begin
          scan_seq_seg_next_state = LOOKUP;
        end
      end
    default: scan_seq_seg_next_state = scan_seq_seg_current_state;
  endcase
end
always_comb begin
  unique case (scan_seq_seg_current_state)
    DONE_SEG: begin :scan_seq_seg_DONE_SEG_Output
        seg_addr_out_to_fifo = 16'h0;
        seg_op_out_to_fifo = 16'h0;
        seg_ID_out_to_fifo = 16'h0;
        seg_req_push = 1'h0;
        seg_rd_rsp_fifo_pop = 1'h1;
        seg_pop_infifo = 1'h0;
        inc_req_made_seg = 1'h0;
        clr_req_made_seg = 1'h0;
        inc_req_rec_seg = 1'h0;
        clr_req_rec_seg = 1'h0;
        us_fifo_inject_data = 16'h0;
        us_fifo_inject_eos = 1'h0;
        us_fifo_inject_push = 1'h0;
        seg_res_fifo_push_alloc = 1'h0;
        seg_res_fifo_push_fill = 1'h0;
        seg_res_fifo_fill_data_in = 17'h0;
        set_readout_loop_seg = go_to_readout_sticky_sticky & (~readout_loop_sticky_sticky) & spacc_mode &
            (crd_in_done_state | lookup);
        clr_readout_loop_seg = readout_loop_sticky_sticky & spacc_mode & (crd_in_done_state | lookup);
        seg_in_done_state = 1'h1;
        seg_in_start_state = 1'h0;
        set_pushed_done_seg = 1'h0;
        clr_pushed_done_seg = 1'h0;
      end :scan_seq_seg_DONE_SEG_Output
    FREE_SEG: begin :scan_seq_seg_FREE_SEG_Output
        seg_addr_out_to_fifo = 16'h0;
        seg_op_out_to_fifo = 16'h0;
        seg_ID_out_to_fifo = 16'h0;
        seg_req_push = 1'h1;
        seg_rd_rsp_fifo_pop = 1'h1;
        seg_pop_infifo = 1'h0;
        inc_req_made_seg = 1'h0;
        clr_req_made_seg = 1'h0;
        inc_req_rec_seg = 1'h0;
        clr_req_rec_seg = 1'h0;
        us_fifo_inject_data = 16'h0;
        us_fifo_inject_eos = 1'h0;
        us_fifo_inject_push = 1'h0;
        seg_res_fifo_push_alloc = 1'h0;
        seg_res_fifo_push_fill = 1'h0;
        seg_res_fifo_fill_data_in = 17'h0;
        seg_in_start_state = 1'h0;
        set_readout_loop_seg = 1'h0;
        seg_in_done_state = 1'h0;
        set_pushed_done_seg = 1'h0;
        clr_pushed_done_seg = 1'h0;
        clr_readout_loop_seg = 1'h0;
      end :scan_seq_seg_FREE_SEG_Output
    INJECT_0: begin :scan_seq_seg_INJECT_0_Output
        seg_addr_out_to_fifo = 16'h0;
        seg_op_out_to_fifo = 16'h0;
        seg_ID_out_to_fifo = 16'h0;
        seg_req_push = 1'h0;
        seg_rd_rsp_fifo_pop = 1'h0;
        seg_pop_infifo = 1'h0;
        inc_req_made_seg = 1'h0;
        clr_req_made_seg = 1'h0;
        inc_req_rec_seg = 1'h0;
        clr_req_rec_seg = 1'h0;
        us_fifo_inject_data = 16'h0;
        us_fifo_inject_eos = 1'h0;
        us_fifo_inject_push = 1'h1;
        seg_res_fifo_push_alloc = 1'h0;
        seg_res_fifo_push_fill = 1'h0;
        seg_res_fifo_fill_data_in = 17'h0;
        seg_in_start_state = 1'h0;
        set_readout_loop_seg = 1'h0;
        seg_in_done_state = 1'h0;
        set_pushed_done_seg = 1'h0;
        clr_pushed_done_seg = 1'h0;
        clr_readout_loop_seg = 1'h0;
      end :scan_seq_seg_INJECT_0_Output
    INJECT_DONE: begin :scan_seq_seg_INJECT_DONE_Output
        seg_addr_out_to_fifo = 16'h0;
        seg_op_out_to_fifo = 16'h0;
        seg_ID_out_to_fifo = 16'h0;
        seg_req_push = 1'h0;
        seg_rd_rsp_fifo_pop = 1'h0;
        seg_pop_infifo = 1'h0;
        inc_req_made_seg = 1'h0;
        clr_req_made_seg = 1'h0;
        inc_req_rec_seg = 1'h0;
        clr_req_rec_seg = 1'h0;
        us_fifo_inject_data = 16'h100;
        us_fifo_inject_eos = 1'h1;
        us_fifo_inject_push = 1'h1;
        seg_res_fifo_push_alloc = 1'h0;
        seg_res_fifo_push_fill = 1'h0;
        seg_res_fifo_fill_data_in = 17'h0;
        seg_in_start_state = 1'h0;
        set_readout_loop_seg = 1'h0;
        seg_in_done_state = 1'h0;
        set_pushed_done_seg = 1'h0;
        clr_pushed_done_seg = 1'h0;
        clr_readout_loop_seg = 1'h0;
      end :scan_seq_seg_INJECT_DONE_Output
    INJECT_ROUTING: begin :scan_seq_seg_INJECT_ROUTING_Output
        seg_addr_out_to_fifo = 16'h0;
        seg_op_out_to_fifo = 16'h0;
        seg_ID_out_to_fifo = 16'h0;
        seg_req_push = 1'h0;
        seg_rd_rsp_fifo_pop = 1'h0;
        seg_pop_infifo = 1'h0;
        inc_req_made_seg = 1'h0;
        clr_req_made_seg = 1'h0;
        inc_req_rec_seg = 1'h0;
        clr_req_rec_seg = 1'h0;
        us_fifo_inject_data = 16'h0;
        us_fifo_inject_eos = 1'h0;
        us_fifo_inject_push = 1'h1;
        seg_res_fifo_push_alloc = ~seg_res_fifo_full;
        seg_res_fifo_push_fill = ~seg_res_fifo_full;
        seg_res_fifo_fill_data_in = {1'h1, 6'h0, 2'h3, 7'h0, readout_loop_sticky_sticky};
        seg_in_start_state = 1'h0;
        set_readout_loop_seg = 1'h0;
        seg_in_done_state = 1'h0;
        set_pushed_done_seg = 1'h0;
        clr_pushed_done_seg = 1'h0;
        clr_readout_loop_seg = 1'h0;
      end :scan_seq_seg_INJECT_ROUTING_Output
    LOOKUP: begin :scan_seq_seg_LOOKUP_Output
        seg_addr_out_to_fifo = infifo_pos_in;
        seg_op_out_to_fifo = 16'h1;
        seg_ID_out_to_fifo = 16'h0;
        seg_req_push = infifo_valid_in & (~infifo_eos_in) & (~crd_res_fifo_full);
        seg_rd_rsp_fifo_pop = 1'h1;
        seg_pop_infifo = infifo_valid_in & (~crd_res_fifo_full) & (infifo_eos_in ? 1'h1: seg_grant_push);
        inc_req_made_seg = 1'h0;
        clr_req_made_seg = 1'h1;
        inc_req_rec_seg = 1'h0;
        clr_req_rec_seg = 1'h1;
        us_fifo_inject_data = 16'h0;
        us_fifo_inject_eos = 1'h0;
        us_fifo_inject_push = 1'h0;
        seg_res_fifo_push_alloc = (~crd_res_fifo_full) & (seg_grant_push | (infifo_valid_in & infifo_eos_in));
        seg_res_fifo_push_fill = infifo_valid_in & infifo_eos_in & (~crd_res_fifo_full);
        seg_res_fifo_fill_data_in = (infifo_eos_in & (infifo_pos_in[9:8] == 2'h2)) ? 17'h0: {infifo_eos_in,
            infifo_pos_in};
        set_pushed_done_seg = done_in & (~crd_res_fifo_full) & spacc_mode;
        set_readout_loop_seg = done_in & (~crd_res_fifo_full) & spacc_mode;
        seg_in_start_state = 1'h0;
        seg_in_done_state = 1'h0;
        clr_pushed_done_seg = 1'h0;
        clr_readout_loop_seg = 1'h0;
      end :scan_seq_seg_LOOKUP_Output
    PASS_DONE_SEG: begin :scan_seq_seg_PASS_DONE_SEG_Output
        seg_addr_out_to_fifo = 16'h0;
        seg_op_out_to_fifo = 16'h0;
        seg_ID_out_to_fifo = 16'h0;
        seg_req_push = 1'h0;
        seg_rd_rsp_fifo_pop = 1'h1;
        seg_pop_infifo = (~readout_loop_sticky_sticky) & done_in & (~seg_res_fifo_full);
        inc_req_made_seg = 1'h0;
        clr_req_made_seg = 1'h0;
        inc_req_rec_seg = 1'h0;
        clr_req_rec_seg = 1'h0;
        us_fifo_inject_data = 16'h0;
        us_fifo_inject_eos = 1'h0;
        us_fifo_inject_push = 1'h0;
        seg_res_fifo_push_alloc = ((readout_loop_sticky_sticky & pushed_done_sticky_sticky) |
            ((~readout_loop_sticky_sticky) & last_stop_done)) & (~seg_res_fifo_full);
        seg_res_fifo_push_fill = ((readout_loop_sticky_sticky & pushed_done_sticky_sticky) |
            ((~readout_loop_sticky_sticky) & last_stop_done)) & (~seg_res_fifo_full);
        seg_res_fifo_fill_data_in = {1'h1, 6'h0, 2'h1, 8'h0};
        set_pushed_done_seg = last_stop_done & (~seg_res_fifo_full) & spacc_mode;
        seg_in_start_state = 1'h0;
        set_readout_loop_seg = 1'h0;
        seg_in_done_state = 1'h0;
        clr_pushed_done_seg = 1'h0;
        clr_readout_loop_seg = 1'h0;
      end :scan_seq_seg_PASS_DONE_SEG_Output
    PASS_STOP_SEG: begin :scan_seq_seg_PASS_STOP_SEG_Output
        seg_addr_out_to_fifo = 16'h0;
        seg_op_out_to_fifo = 16'h0;
        seg_ID_out_to_fifo = 16'h0;
        seg_req_push = 1'h0;
        seg_rd_rsp_fifo_pop = 1'h1;
        seg_pop_infifo = (~seg_res_fifo_full) & eos_in & (~readout_loop_sticky_sticky);
        inc_req_made_seg = 1'h0;
        clr_req_made_seg = 1'h1;
        inc_req_rec_seg = 1'h0;
        clr_req_rec_seg = 1'h1;
        us_fifo_inject_data = 16'h0;
        us_fifo_inject_eos = 1'h0;
        us_fifo_inject_push = 1'h0;
        seg_res_fifo_push_alloc = (infifo_valid_in | readout_loop_sticky_sticky) & (~seg_res_fifo_full);
        seg_res_fifo_push_fill = (infifo_valid_in | readout_loop_sticky_sticky) & (~seg_res_fifo_full);
        seg_res_fifo_fill_data_in = readout_loop_sticky_sticky ? last_stop_token - 17'h1: eos_in ? {1'h1,
            infifo_pos_in + 16'h1}: {1'h1, 16'h0};
        seg_in_start_state = 1'h0;
        set_readout_loop_seg = 1'h0;
        seg_in_done_state = 1'h0;
        set_pushed_done_seg = 1'h0;
        clr_pushed_done_seg = 1'h0;
        clr_readout_loop_seg = 1'h0;
      end :scan_seq_seg_PASS_STOP_SEG_Output
    READ: begin :scan_seq_seg_READ_Output
        seg_addr_out_to_fifo = readout_loop_sticky_sticky ? 16'h0: infifo_pos_in;
        seg_op_out_to_fifo = 16'h1;
        seg_ID_out_to_fifo = 16'h0;
        seg_req_push = ((infifo_valid_in & (~infifo_eos_in) & (~dense)) | readout_loop_sticky_sticky) &
            (~seg_res_fifo_full);
        seg_rd_rsp_fifo_pop = 1'h1;
        seg_pop_infifo = (((done_in | (dense & infifo_valid_in)) & (~seg_res_fifo_full)) | maybe_in) &
            (~readout_loop_sticky_sticky);
        inc_req_made_seg = 1'h0;
        clr_req_made_seg = 1'h0;
        inc_req_rec_seg = 1'h0;
        clr_req_rec_seg = 1'h0;
        us_fifo_inject_data = 16'h0;
        us_fifo_inject_eos = 1'h0;
        us_fifo_inject_push = 1'h0;
        seg_res_fifo_push_alloc = (done_in | dense) ? (~seg_res_fifo_full) & infifo_valid_in: (~seg_res_fifo_full)
            & seg_grant_push & (~maybe_in);
        seg_res_fifo_push_fill = (done_in | (dense & infifo_valid_in)) & (~seg_res_fifo_full);
        seg_res_fifo_fill_data_in = {infifo_eos_in, infifo_pos_in};
        seg_in_start_state = 1'h0;
        set_readout_loop_seg = 1'h0;
        seg_in_done_state = 1'h0;
        set_pushed_done_seg = 1'h0;
        clr_pushed_done_seg = 1'h0;
        clr_readout_loop_seg = 1'h0;
      end :scan_seq_seg_READ_Output
    READ_ALT: begin :scan_seq_seg_READ_ALT_Output
        seg_addr_out_to_fifo = readout_loop_sticky_sticky ? 16'h1: infifo_pos_in + 16'h1;
        seg_op_out_to_fifo = 16'h1;
        seg_ID_out_to_fifo = 16'h0;
        seg_req_push = ~seg_res_fifo_full;
        seg_rd_rsp_fifo_pop = 1'h1;
        seg_pop_infifo = seg_grant_push & (~seg_res_fifo_full) & (~readout_loop_sticky_sticky);
        inc_req_made_seg = 1'h0;
        clr_req_made_seg = 1'h0;
        inc_req_rec_seg = 1'h0;
        clr_req_rec_seg = 1'h0;
        us_fifo_inject_data = 16'h0;
        us_fifo_inject_eos = 1'h0;
        us_fifo_inject_push = 1'h0;
        seg_res_fifo_push_alloc = 1'h0;
        seg_res_fifo_push_fill = 1'h0;
        seg_res_fifo_fill_data_in = 17'h0;
        seg_in_start_state = 1'h0;
        set_readout_loop_seg = 1'h0;
        seg_in_done_state = 1'h0;
        set_pushed_done_seg = 1'h0;
        clr_pushed_done_seg = 1'h0;
        clr_readout_loop_seg = 1'h0;
      end :scan_seq_seg_READ_ALT_Output
    START_SEG: begin :scan_seq_seg_START_SEG_Output
        seg_addr_out_to_fifo = 16'h0;
        seg_op_out_to_fifo = 16'h0;
        seg_ID_out_to_fifo = 16'h0;
        seg_req_push = 1'h0;
        seg_rd_rsp_fifo_pop = 1'h0;
        seg_pop_infifo = 1'h0;
        inc_req_made_seg = 1'h0;
        clr_req_made_seg = 1'h0;
        inc_req_rec_seg = 1'h0;
        clr_req_rec_seg = 1'h0;
        us_fifo_inject_data = 16'h0;
        us_fifo_inject_eos = 1'h0;
        us_fifo_inject_push = 1'h0;
        seg_res_fifo_push_alloc = 1'h0;
        seg_res_fifo_push_fill = 1'h0;
        seg_res_fifo_fill_data_in = 17'h0;
        set_readout_loop_seg = 1'h0;
        seg_in_start_state = 1'h1;
        seg_in_done_state = 1'h0;
        set_pushed_done_seg = 1'h0;
        clr_pushed_done_seg = 1'h0;
        clr_readout_loop_seg = 1'h0;
      end :scan_seq_seg_START_SEG_Output
    default: begin :scan_seq_seg_default_Output
        seg_addr_out_to_fifo = 16'h0;
        seg_op_out_to_fifo = 16'h0;
        seg_ID_out_to_fifo = 16'h0;
        seg_req_push = 1'h0;
        seg_rd_rsp_fifo_pop = 1'h0;
        seg_pop_infifo = 1'h0;
        inc_req_made_seg = 1'h0;
        clr_req_made_seg = 1'h0;
        inc_req_rec_seg = 1'h0;
        clr_req_rec_seg = 1'h0;
        us_fifo_inject_data = 16'h0;
        us_fifo_inject_eos = 1'h0;
        us_fifo_inject_push = 1'h0;
        seg_res_fifo_push_alloc = 1'h0;
        seg_res_fifo_push_fill = 1'h0;
        seg_res_fifo_fill_data_in = 17'h0;
        set_readout_loop_seg = 1'h0;
        seg_in_start_state = 1'h1;
        seg_in_done_state = 1'h0;
        set_pushed_done_seg = 1'h0;
        clr_pushed_done_seg = 1'h0;
        clr_readout_loop_seg = 1'h0;
      end :scan_seq_seg_default_Output
  endcase
end
reg_fifo_depth_2_w_17_afd_2 input_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(fifo_us_in_packed),
  .flush(flush),
  .pop(pop_infifo),
  .push(us_fifo_push),
  .rst_n(rst_n),
  .data_out(input_fifo_data_out),
  .empty(input_fifo_empty),
  .full(fifo_us_full)
);

reg_fifo_depth_2_w_17_afd_2 rd_rsp_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(rd_rsp_data_in[0]),
  .flush(flush),
  .pop(1'h1),
  .push(rd_rsp_data_in_valid),
  .rst_n(rst_n),
  .data_out(rd_rsp_fifo_out_data),
  .empty(rd_rsp_fifo_empty),
  .full(rd_rsp_fifo_full)
);

arbiter_2_in_RR_algo rr_arbiter (
  .clk(gclk),
  .clk_en(clk_en),
  .flush(flush),
  .request_in(base_rr),
  .resource_ready(no_outfifo_full),
  .rst_n(rst_n),
  .grant_out(rr_arbiter_grant_out)
);

reg_fifo_depth_2_w_17_afd_2 addr_out_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(addr_out_fifo_data_in),
  .flush(flush),
  .pop(addr_out_ready),
  .push(addr_out_fifo_push),
  .rst_n(rst_n),
  .data_out(addr_out),
  .empty(addr_out_fifo_empty),
  .full(addr_out_fifo_full)
);

reg_fifo_depth_2_w_17_afd_2 op_out_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(op_out_fifo_data_in),
  .flush(flush),
  .pop(op_out_ready),
  .push(op_out_fifo_push),
  .rst_n(rst_n),
  .data_out(op_out),
  .empty(op_out_fifo_empty),
  .full(op_out_fifo_full)
);

reg_fifo_depth_2_w_17_afd_2 ID_out_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(ID_out_fifo_data_in),
  .flush(flush),
  .pop(ID_out_ready),
  .push(ID_out_fifo_push),
  .rst_n(rst_n),
  .data_out(ID_out),
  .empty(ID_out_fifo_empty),
  .full(ID_out_fifo_full)
);

reservation_fifo_depth_8_w_17_num_per_2 seg_res_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in_0(rd_rsp_fifo_out_data),
  .data_in_1(rd_rsp_fifo_out_data),
  .fill_data_in(seg_res_fifo_fill_data_in),
  .flush(flush),
  .pop(seg_res_fifo_pop_0),
  .push_alloc(seg_res_fifo_push_alloc_0),
  .push_fill(seg_res_fifo_push_fill_0),
  .push_reserve(seg_res_fifo_push_reserve_0),
  .rst_n(rst_n),
  .data_out_0(seg_res_fifo_data_out_0),
  .data_out_1(seg_res_fifo_data_out_1),
  .full(seg_res_fifo_full),
  .valid(seg_res_fifo_valid)
);

reservation_fifo_depth_8_w_17_num_per_1 crd_res_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in_0(crd_res_fifo_data_in_0),
  .fill_data_in(crd_res_fifo_fill_data_in),
  .flush(flush),
  .pop(crd_res_fifo_pop),
  .push_alloc(crd_res_fifo_push_alloc_0),
  .push_fill(crd_res_fifo_push_fill_0),
  .push_reserve(crd_res_fifo_push_reserve_0),
  .rst_n(rst_n),
  .data_out_0(crd_res_fifo_data_out),
  .full(crd_res_fifo_full),
  .valid(crd_res_fifo_valid)
);

reg_fifo_depth_0_w_17_afd_2 coordinate_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(coord_fifo_in_packed),
  .flush(flush),
  .pop(coord_out_ready),
  .push(coordinate_fifo_push),
  .rst_n(rst_n),
  .data_out(coord_fifo_out_packed),
  .empty(coordinate_fifo_empty),
  .full(coordinate_fifo_full)
);

reg_fifo_depth_0_w_17_afd_2 pos_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(pos_fifo_in_packed),
  .flush(flush),
  .pop(pos_out_ready),
  .push(pos_out_fifo_push),
  .rst_n(rst_n),
  .data_out(pos_fifo_out_packed),
  .empty(pos_fifo_empty),
  .full(pos_fifo_full)
);

reg_fifo_depth_0_w_17_afd_2 block_rd_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(crd_res_fifo_data_out),
  .flush(flush),
  .pop(block_rd_out_ready),
  .push(block_rd_fifo_push),
  .rst_n(rst_n),
  .data_out(block_rd_out),
  .empty(block_rd_fifo_empty),
  .full(block_rd_fifo_full)
);

endmodule   // scanner_pipe

module sched_gen_3_16 (
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic enable,
  input logic finished,
  input logic flush,
  input logic [1:0] mux_sel,
  input logic rst_n,
  input logic [15:0] sched_addr_gen_starting_addr,
  input logic [15:0] sched_addr_gen_strides_0,
  input logic [15:0] sched_addr_gen_strides_1,
  input logic [15:0] sched_addr_gen_strides_2,
  output logic valid_output
);

logic [15:0] addr_out;
logic [2:0][15:0] sched_addr_gen_strides;
logic valid_gate;
logic valid_gate_inv;
logic valid_out;
assign valid_gate = ~valid_gate_inv;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    valid_gate_inv <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      valid_gate_inv <= 1'h0;
    end
    else if (finished) begin
      valid_gate_inv <= 1'h1;
    end
  end
end
always_comb begin
  valid_out = (cycle_count == addr_out) & valid_gate & enable;
end
always_comb begin
  valid_output = valid_out;
end
assign sched_addr_gen_strides[0] = sched_addr_gen_strides_0;
assign sched_addr_gen_strides[1] = sched_addr_gen_strides_1;
assign sched_addr_gen_strides[2] = sched_addr_gen_strides_2;
addr_gen_3_16 sched_addr_gen (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(mux_sel),
  .restart(finished),
  .rst_n(rst_n),
  .starting_addr(sched_addr_gen_starting_addr),
  .step(valid_out),
  .strides(sched_addr_gen_strides),
  .addr_out(addr_out)
);

endmodule   // sched_gen_3_16

module sched_gen_6_16 (
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic enable,
  input logic finished,
  input logic flush,
  input logic [2:0] mux_sel,
  input logic rst_n,
  input logic [15:0] sched_addr_gen_starting_addr,
  input logic [15:0] sched_addr_gen_strides_0,
  input logic [15:0] sched_addr_gen_strides_1,
  input logic [15:0] sched_addr_gen_strides_2,
  input logic [15:0] sched_addr_gen_strides_3,
  input logic [15:0] sched_addr_gen_strides_4,
  input logic [15:0] sched_addr_gen_strides_5,
  output logic valid_output
);

logic [15:0] addr_out;
logic [5:0][15:0] sched_addr_gen_strides;
logic valid_gate;
logic valid_gate_inv;
logic valid_out;
assign valid_gate = ~valid_gate_inv;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    valid_gate_inv <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      valid_gate_inv <= 1'h0;
    end
    else if (finished) begin
      valid_gate_inv <= 1'h1;
    end
  end
end
always_comb begin
  valid_out = (cycle_count == addr_out) & valid_gate & enable;
end
always_comb begin
  valid_output = valid_out;
end
assign sched_addr_gen_strides[0] = sched_addr_gen_strides_0;
assign sched_addr_gen_strides[1] = sched_addr_gen_strides_1;
assign sched_addr_gen_strides[2] = sched_addr_gen_strides_2;
assign sched_addr_gen_strides[3] = sched_addr_gen_strides_3;
assign sched_addr_gen_strides[4] = sched_addr_gen_strides_4;
assign sched_addr_gen_strides[5] = sched_addr_gen_strides_5;
addr_gen_6_16 sched_addr_gen (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(mux_sel),
  .restart(finished),
  .rst_n(rst_n),
  .starting_addr(sched_addr_gen_starting_addr),
  .step(valid_out),
  .strides(sched_addr_gen_strides),
  .addr_out(addr_out)
);

endmodule   // sched_gen_6_16

module sched_gen_6_16_delay_addr_10_4 (
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic enable,
  input logic finished,
  input logic flush,
  input logic [2:0] mux_sel,
  input logic rst_n,
  input logic [9:0] sched_addr_gen_delay,
  input logic [15:0] sched_addr_gen_starting_addr,
  input logic [15:0] sched_addr_gen_strides_0,
  input logic [15:0] sched_addr_gen_strides_1,
  input logic [15:0] sched_addr_gen_strides_2,
  input logic [15:0] sched_addr_gen_strides_3,
  input logic [15:0] sched_addr_gen_strides_4,
  input logic [15:0] sched_addr_gen_strides_5,
  output logic delay_en_out,
  output logic valid_output,
  output logic valid_output_d
);

logic [3:0][10:0] addr_fifo;
logic addr_fifo_empty_n;
logic [10:0] addr_fifo_in;
logic [10:0] addr_fifo_out;
logic addr_fifo_wr_en;
logic [15:0] addr_out;
logic [15:0] addr_out_d;
logic delay_en;
logic [1:0] next_rd_ptr;
logic [1:0] rd_ptr;
logic [9:0] sched_addr_gen_delay_out;
logic [5:0][15:0] sched_addr_gen_strides;
logic valid_gate;
logic valid_gate_inv;
logic valid_out;
logic valid_out_d;
logic [1:0] wr_ptr;
assign valid_gate = ~valid_gate_inv;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    valid_gate_inv <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      valid_gate_inv <= 1'h0;
    end
    else if (finished) begin
      valid_gate_inv <= 1'h1;
    end
  end
end
assign delay_en_out = delay_en;
assign delay_en = sched_addr_gen_delay_out > 10'h0;
assign next_rd_ptr = rd_ptr + 2'h1;
assign addr_fifo_wr_en = valid_out;
assign addr_fifo_in = addr_out_d[10:0];
assign addr_fifo_out = addr_fifo[rd_ptr];

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    wr_ptr <= 2'h0;
    rd_ptr <= 2'h0;
    addr_fifo <= 44'h0;
    addr_fifo_empty_n <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      wr_ptr <= 2'h0;
      rd_ptr <= 2'h0;
      addr_fifo <= 44'h0;
      addr_fifo_empty_n <= 1'h0;
    end
    else if (delay_en) begin
      if (addr_fifo_wr_en) begin
        wr_ptr <= wr_ptr + 2'h1;
        addr_fifo[wr_ptr] <= addr_fifo_in;
      end
      if (valid_out_d) begin
        rd_ptr <= next_rd_ptr;
      end
      if (addr_fifo_wr_en) begin
        addr_fifo_empty_n <= 1'h1;
      end
      else if (valid_out_d) begin
        addr_fifo_empty_n <= ~(next_rd_ptr == wr_ptr);
      end
      else addr_fifo_empty_n <= addr_fifo_empty_n;
    end
  end
end
always_comb begin
  valid_out_d = (cycle_count[10:0] == addr_fifo_out) & addr_fifo_empty_n & enable;
  valid_output_d = valid_out_d;
end
always_comb begin
  valid_out = (cycle_count == addr_out) & valid_gate & enable;
end
always_comb begin
  valid_output = valid_out;
end
assign sched_addr_gen_strides[0] = sched_addr_gen_strides_0;
assign sched_addr_gen_strides[1] = sched_addr_gen_strides_1;
assign sched_addr_gen_strides[2] = sched_addr_gen_strides_2;
assign sched_addr_gen_strides[3] = sched_addr_gen_strides_3;
assign sched_addr_gen_strides[4] = sched_addr_gen_strides_4;
assign sched_addr_gen_strides[5] = sched_addr_gen_strides_5;
addr_gen_6_16_delay_addr_10 sched_addr_gen (
  .clk(clk),
  .clk_en(clk_en),
  .delay(sched_addr_gen_delay),
  .flush(flush),
  .mux_sel(mux_sel),
  .restart(finished),
  .rst_n(rst_n),
  .starting_addr(sched_addr_gen_starting_addr),
  .step(valid_out),
  .strides(sched_addr_gen_strides),
  .addr_out(addr_out),
  .delay_out(sched_addr_gen_delay_out),
  .delayed_addr_out(addr_out_d)
);

endmodule   // sched_gen_6_16_delay_addr_10_4

module sched_gen_6_16_delay_addr_10_8 (
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic enable,
  input logic finished,
  input logic flush,
  input logic [2:0] mux_sel,
  input logic rst_n,
  input logic [9:0] sched_addr_gen_delay,
  input logic [15:0] sched_addr_gen_starting_addr,
  input logic [15:0] sched_addr_gen_strides_0,
  input logic [15:0] sched_addr_gen_strides_1,
  input logic [15:0] sched_addr_gen_strides_2,
  input logic [15:0] sched_addr_gen_strides_3,
  input logic [15:0] sched_addr_gen_strides_4,
  input logic [15:0] sched_addr_gen_strides_5,
  output logic delay_en_out,
  output logic valid_output,
  output logic valid_output_d
);

logic [7:0][10:0] addr_fifo;
logic addr_fifo_empty_n;
logic [10:0] addr_fifo_in;
logic [10:0] addr_fifo_out;
logic addr_fifo_wr_en;
logic [15:0] addr_out;
logic [15:0] addr_out_d;
logic delay_en;
logic [2:0] next_rd_ptr;
logic [2:0] rd_ptr;
logic [9:0] sched_addr_gen_delay_out;
logic [5:0][15:0] sched_addr_gen_strides;
logic valid_gate;
logic valid_gate_inv;
logic valid_out;
logic valid_out_d;
logic [2:0] wr_ptr;
assign valid_gate = ~valid_gate_inv;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    valid_gate_inv <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      valid_gate_inv <= 1'h0;
    end
    else if (finished) begin
      valid_gate_inv <= 1'h1;
    end
  end
end
assign delay_en_out = delay_en;
assign delay_en = sched_addr_gen_delay_out > 10'h0;
assign next_rd_ptr = rd_ptr + 3'h1;
assign addr_fifo_wr_en = valid_out;
assign addr_fifo_in = addr_out_d[10:0];
assign addr_fifo_out = addr_fifo[rd_ptr];

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    wr_ptr <= 3'h0;
    rd_ptr <= 3'h0;
    addr_fifo <= 88'h0;
    addr_fifo_empty_n <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      wr_ptr <= 3'h0;
      rd_ptr <= 3'h0;
      addr_fifo <= 88'h0;
      addr_fifo_empty_n <= 1'h0;
    end
    else if (delay_en) begin
      if (addr_fifo_wr_en) begin
        wr_ptr <= wr_ptr + 3'h1;
        addr_fifo[wr_ptr] <= addr_fifo_in;
      end
      if (valid_out_d) begin
        rd_ptr <= next_rd_ptr;
      end
      if (addr_fifo_wr_en) begin
        addr_fifo_empty_n <= 1'h1;
      end
      else if (valid_out_d) begin
        addr_fifo_empty_n <= ~(next_rd_ptr == wr_ptr);
      end
      else addr_fifo_empty_n <= addr_fifo_empty_n;
    end
  end
end
always_comb begin
  valid_out_d = (cycle_count[10:0] == addr_fifo_out) & addr_fifo_empty_n & enable;
  valid_output_d = valid_out_d;
end
always_comb begin
  valid_out = (cycle_count == addr_out) & valid_gate & enable;
end
always_comb begin
  valid_output = valid_out;
end
assign sched_addr_gen_strides[0] = sched_addr_gen_strides_0;
assign sched_addr_gen_strides[1] = sched_addr_gen_strides_1;
assign sched_addr_gen_strides[2] = sched_addr_gen_strides_2;
assign sched_addr_gen_strides[3] = sched_addr_gen_strides_3;
assign sched_addr_gen_strides[4] = sched_addr_gen_strides_4;
assign sched_addr_gen_strides[5] = sched_addr_gen_strides_5;
addr_gen_6_16_delay_addr_10 sched_addr_gen (
  .clk(clk),
  .clk_en(clk_en),
  .delay(sched_addr_gen_delay),
  .flush(flush),
  .mux_sel(mux_sel),
  .restart(finished),
  .rst_n(rst_n),
  .starting_addr(sched_addr_gen_starting_addr),
  .step(valid_out),
  .strides(sched_addr_gen_strides),
  .addr_out(addr_out),
  .delay_out(sched_addr_gen_delay_out),
  .delayed_addr_out(addr_out_d)
);

endmodule   // sched_gen_6_16_delay_addr_10_8

module sram_sp__0 (
  input logic clk,
  input logic clk_en,
  input logic [63:0] data_in_p0,
  input logic flush,
  input logic [8:0] read_addr_p0,
  input logic read_enable_p0,
  input logic [8:0] write_addr_p0,
  input logic write_enable_p0,
  output logic [63:0] data_out_p0
);

logic [63:0] data_array [511:0];

always_ff @(posedge clk) begin
  if (clk_en) begin
    if (write_enable_p0 == 1'h1) begin
      data_array[write_addr_p0] <= data_in_p0;
    end
    else if (read_enable_p0) begin
      data_out_p0 <= data_array[read_addr_p0];
    end
  end
end
endmodule   // sram_sp__0

module stencil_valid (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [3:0] loops_stencil_valid_dimensionality,
  input logic [10:0] loops_stencil_valid_ranges_0,
  input logic [10:0] loops_stencil_valid_ranges_1,
  input logic [10:0] loops_stencil_valid_ranges_2,
  input logic [10:0] loops_stencil_valid_ranges_3,
  input logic [10:0] loops_stencil_valid_ranges_4,
  input logic [10:0] loops_stencil_valid_ranges_5,
  input logic rst_n,
  input logic stencil_valid_sched_gen_enable,
  input logic [15:0] stencil_valid_sched_gen_sched_addr_gen_starting_addr,
  input logic [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_0,
  input logic [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_1,
  input logic [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_2,
  input logic [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_3,
  input logic [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_4,
  input logic [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_5,
  output logic stencil_valid
);

logic [15:0] cycle_count;
logic flushed;
logic [2:0] loops_stencil_valid_mux_sel_out;
logic [5:0][10:0] loops_stencil_valid_ranges;
logic loops_stencil_valid_restart;
logic stencil_valid_internal;
assign stencil_valid = stencil_valid_internal & flushed;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    cycle_count <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      cycle_count <= 16'h0;
    end
    else if (flushed) begin
      cycle_count <= cycle_count + 16'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    flushed <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      flushed <= 1'h1;
    end
  end
end
assign loops_stencil_valid_ranges[0] = loops_stencil_valid_ranges_0;
assign loops_stencil_valid_ranges[1] = loops_stencil_valid_ranges_1;
assign loops_stencil_valid_ranges[2] = loops_stencil_valid_ranges_2;
assign loops_stencil_valid_ranges[3] = loops_stencil_valid_ranges_3;
assign loops_stencil_valid_ranges[4] = loops_stencil_valid_ranges_4;
assign loops_stencil_valid_ranges[5] = loops_stencil_valid_ranges_5;
for_loop_6_11 loops_stencil_valid (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_stencil_valid_dimensionality),
  .flush(flush),
  .ranges(loops_stencil_valid_ranges),
  .rst_n(rst_n),
  .step(stencil_valid_internal),
  .mux_sel_out(loops_stencil_valid_mux_sel_out),
  .restart(loops_stencil_valid_restart)
);

sched_gen_6_16 stencil_valid_sched_gen (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(stencil_valid_sched_gen_enable),
  .finished(loops_stencil_valid_restart),
  .flush(flush),
  .mux_sel(loops_stencil_valid_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(stencil_valid_sched_gen_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides_0(stencil_valid_sched_gen_sched_addr_gen_strides_0),
  .sched_addr_gen_strides_1(stencil_valid_sched_gen_sched_addr_gen_strides_1),
  .sched_addr_gen_strides_2(stencil_valid_sched_gen_sched_addr_gen_strides_2),
  .sched_addr_gen_strides_3(stencil_valid_sched_gen_sched_addr_gen_strides_3),
  .sched_addr_gen_strides_4(stencil_valid_sched_gen_sched_addr_gen_strides_4),
  .sched_addr_gen_strides_5(stencil_valid_sched_gen_sched_addr_gen_strides_5),
  .valid_output(stencil_valid_internal)
);

endmodule   // stencil_valid

module stencil_valid_flat (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic rst_n,
  input logic [3:0] stencil_valid_inst_loops_stencil_valid_dimensionality,
  input logic [10:0] stencil_valid_inst_loops_stencil_valid_ranges_0,
  input logic [10:0] stencil_valid_inst_loops_stencil_valid_ranges_1,
  input logic [10:0] stencil_valid_inst_loops_stencil_valid_ranges_2,
  input logic [10:0] stencil_valid_inst_loops_stencil_valid_ranges_3,
  input logic [10:0] stencil_valid_inst_loops_stencil_valid_ranges_4,
  input logic [10:0] stencil_valid_inst_loops_stencil_valid_ranges_5,
  input logic stencil_valid_inst_stencil_valid_sched_gen_enable,
  input logic [15:0] stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr,
  input logic [15:0] stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0,
  input logic [15:0] stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1,
  input logic [15:0] stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2,
  input logic [15:0] stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3,
  input logic [15:0] stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4,
  input logic [15:0] stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5,
  output logic stencil_valid_f_
);

stencil_valid stencil_valid_inst (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .loops_stencil_valid_dimensionality(stencil_valid_inst_loops_stencil_valid_dimensionality),
  .loops_stencil_valid_ranges_0(stencil_valid_inst_loops_stencil_valid_ranges_0),
  .loops_stencil_valid_ranges_1(stencil_valid_inst_loops_stencil_valid_ranges_1),
  .loops_stencil_valid_ranges_2(stencil_valid_inst_loops_stencil_valid_ranges_2),
  .loops_stencil_valid_ranges_3(stencil_valid_inst_loops_stencil_valid_ranges_3),
  .loops_stencil_valid_ranges_4(stencil_valid_inst_loops_stencil_valid_ranges_4),
  .loops_stencil_valid_ranges_5(stencil_valid_inst_loops_stencil_valid_ranges_5),
  .rst_n(rst_n),
  .stencil_valid_sched_gen_enable(stencil_valid_inst_stencil_valid_sched_gen_enable),
  .stencil_valid_sched_gen_sched_addr_gen_starting_addr(stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_starting_addr),
  .stencil_valid_sched_gen_sched_addr_gen_strides_0(stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_0),
  .stencil_valid_sched_gen_sched_addr_gen_strides_1(stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_1),
  .stencil_valid_sched_gen_sched_addr_gen_strides_2(stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_2),
  .stencil_valid_sched_gen_sched_addr_gen_strides_3(stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_3),
  .stencil_valid_sched_gen_sched_addr_gen_strides_4(stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_4),
  .stencil_valid_sched_gen_sched_addr_gen_strides_5(stencil_valid_inst_stencil_valid_sched_gen_sched_addr_gen_strides_5),
  .stencil_valid(stencil_valid_f_)
);

endmodule   // stencil_valid_flat

module storage_config_seq_2_64_16 (
  input logic clk,
  input logic clk_en,
  input logic [7:0] config_addr_in,
  input logic [15:0] config_data_in,
  input logic [1:0] config_en,
  input logic config_rd,
  input logic config_wr,
  input logic flush,
  input logic [0:0][3:0] [15:0] rd_data_stg,
  input logic rst_n,
  output logic [8:0] addr_out,
  output logic [1:0] [15:0] rd_data_out,
  output logic ren_out,
  output logic wen_out,
  output logic [3:0] [15:0] wr_data
);

logic [1:0] cnt;
logic [2:0][15:0] data_wr_reg;
logic [1:0] rd_cnt;
logic rd_valid;
logic [1:0] reduce_en;
logic set_to_addr;
assign reduce_en[0] = |config_en[0];
assign reduce_en[1] = |config_en[1];
always_comb begin
  set_to_addr = 1'h0;
  for (int unsigned i = 0; i < 2; i += 1) begin
      if (reduce_en[1'(i)]) begin
        set_to_addr = 1'(i);
      end
    end
end
assign addr_out = {set_to_addr, config_addr_in};

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    cnt <= 2'h0;
  end
  else if (flush) begin
    cnt <= 2'h0;
  end
  else if (config_wr & (|config_en)) begin
    cnt <= cnt + 2'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    rd_valid <= 1'h0;
  end
  else if (flush) begin
    rd_valid <= 1'h0;
  end
  else rd_valid <= config_rd & (|config_en);
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    rd_cnt <= 2'h0;
  end
  else if (flush) begin
    rd_cnt <= 2'h0;
  end
  else if (rd_valid & (~(config_rd & (|config_en)))) begin
    rd_cnt <= rd_cnt + 2'h1;
  end
end
assign rd_data_out[0] = rd_data_stg[0][rd_cnt];
assign rd_data_out[1] = rd_data_stg[0][rd_cnt];

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    data_wr_reg <= 48'h0;
  end
  else if (flush) begin
    data_wr_reg <= 48'h0;
  end
  else if (config_wr & (cnt < 2'h3)) begin
    data_wr_reg[cnt] <= config_data_in;
  end
end
assign wr_data[0] = data_wr_reg[0];
assign wr_data[1] = data_wr_reg[1];
assign wr_data[2] = data_wr_reg[2];
assign wr_data[3] = config_data_in;
assign wen_out = config_wr & (cnt == 2'h3);
assign ren_out = config_rd;
endmodule   // storage_config_seq_2_64_16

module strg_ram_64_512_delay1 (
  input logic clk,
  input logic clk_en,
  input logic [0:0][3:0] [15:0] data_from_strg,
  input logic [16:0] data_in,
  input logic flush,
  input logic [16:0] rd_addr_in,
  input logic ren,
  input logic rst_n,
  input logic wen,
  input logic [16:0] wr_addr_in,
  output logic [0:0] [8:0] addr_out,
  output logic [16:0] data_out,
  output logic [0:0][3:0] [15:0] data_to_strg,
  output logic ready,
  output logic ren_to_strg,
  output logic valid_out,
  output logic wen_to_strg
);

typedef enum logic[1:0] {
  IDLE = 2'h0,
  MODIFY = 2'h1,
  READ = 2'h2,
  _DEFAULT = 2'h3
} r_w_seq_state;
logic [15:0] addr_to_write;
logic [3:0][15:0] data_combined;
logic [15:0] data_to_write;
r_w_seq_state r_w_seq_current_state;
r_w_seq_state r_w_seq_next_state;
logic [15:0] rd_addr;
logic rd_bank;
logic read_gate;
logic [15:0] wr_addr;
logic write_gate;
assign wr_addr = wr_addr_in[15:0];
assign rd_addr = wr_addr_in[15:0];
assign rd_bank = 1'h0;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    data_to_write <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      data_to_write <= 16'h0;
    end
    else data_to_write <= data_in[15:0];
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    addr_to_write <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      addr_to_write <= 16'h0;
    end
    else addr_to_write <= wr_addr;
  end
end
assign data_to_strg[0] = data_combined;
assign ren_to_strg = (wen | ren) & read_gate;
assign wen_to_strg = write_gate;
always_comb begin
  addr_out[0] = rd_addr[10:2];
  if (wen & (~write_gate)) begin
    addr_out[0] = wr_addr[10:2];
  end
  else if (write_gate) begin
    addr_out[0] = addr_to_write[10:2];
  end
end
always_comb begin
  if (addr_to_write[1:0] == 2'h0) begin
    data_combined[0] = data_to_write;
  end
  else data_combined[0] = data_from_strg[rd_bank][0];
end
always_comb begin
  if (addr_to_write[1:0] == 2'h1) begin
    data_combined[1] = data_to_write;
  end
  else data_combined[1] = data_from_strg[rd_bank][1];
end
always_comb begin
  if (addr_to_write[1:0] == 2'h2) begin
    data_combined[2] = data_to_write;
  end
  else data_combined[2] = data_from_strg[rd_bank][2];
end
always_comb begin
  if (addr_to_write[1:0] == 2'h3) begin
    data_combined[3] = data_to_write;
  end
  else data_combined[3] = data_from_strg[rd_bank][3];
end

always_ff @(posedge clk, negedge rst_n) begin
  if (!rst_n) begin
    r_w_seq_current_state <= IDLE;
  end
  else r_w_seq_current_state <= r_w_seq_next_state;
end
always_comb begin
  r_w_seq_next_state = r_w_seq_current_state;
  unique case (r_w_seq_current_state)
    IDLE: begin
        if ((~wen) & (~ren)) begin
          r_w_seq_next_state = IDLE;
        end
        else if (ren & (~wen)) begin
          r_w_seq_next_state = READ;
        end
        else if (wen) begin
          r_w_seq_next_state = MODIFY;
        end
      end
    MODIFY: begin
        if (1'h1) begin
          r_w_seq_next_state = IDLE;
        end
      end
    READ: begin
        if ((~wen) & (~ren)) begin
          r_w_seq_next_state = IDLE;
        end
        else if (ren & (~wen)) begin
          r_w_seq_next_state = READ;
        end
        else if (wen) begin
          r_w_seq_next_state = MODIFY;
        end
      end
    _DEFAULT: begin
        if (1'h1) begin
          r_w_seq_next_state = _DEFAULT;
        end
      end
    default: begin end
  endcase
end
always_comb begin
  unique case (r_w_seq_current_state)
    IDLE: begin :r_w_seq_IDLE_Output
        ready = 1'h1;
        valid_out = 1'h0;
        data_out[15:0] = 16'h0;
        data_out[16] = 1'h0;
        write_gate = 1'h0;
        read_gate = 1'h1;
      end :r_w_seq_IDLE_Output
    MODIFY: begin :r_w_seq_MODIFY_Output
        ready = 1'h0;
        valid_out = 1'h0;
        data_out[15:0] = 16'h0;
        data_out[16] = 1'h0;
        write_gate = 1'h1;
        read_gate = 1'h0;
      end :r_w_seq_MODIFY_Output
    READ: begin :r_w_seq_READ_Output
        ready = 1'h1;
        valid_out = 1'h1;
        data_out[15:0] = data_from_strg[rd_bank][addr_to_write[1:0]];
        data_out[16] = 1'h0;
        write_gate = 1'h0;
        read_gate = 1'h1;
      end :r_w_seq_READ_Output
    _DEFAULT: begin :r_w_seq__DEFAULT_Output
        ready = 1'h0;
        valid_out = 1'h0;
        data_out[15:0] = 16'h0;
        data_out[16] = 1'h0;
        write_gate = 1'h0;
        read_gate = 1'h0;
      end :r_w_seq__DEFAULT_Output
    default: begin end
  endcase
end
endmodule   // strg_ram_64_512_delay1

module strg_ram_64_512_delay1_flat (
  input logic clk,
  input logic clk_en,
  input logic [0:0] [16:0] data_in_f_,
  input logic flush,
  input logic [0:0] [16:0] rd_addr_in_f_,
  input logic ren_f_,
  input logic rst_n,
  input logic [0:0][3:0] [15:0] strg_ram_64_512_delay1_inst_data_from_strg_lifted,
  input logic wen_f_,
  input logic [0:0] [16:0] wr_addr_in_f_,
  output logic [0:0] [16:0] data_out_f_,
  output logic ready_f_,
  output logic [0:0] [8:0] strg_ram_64_512_delay1_inst_addr_out_lifted,
  output logic [0:0][3:0] [15:0] strg_ram_64_512_delay1_inst_data_to_strg_lifted,
  output logic strg_ram_64_512_delay1_inst_ren_to_strg_lifted,
  output logic strg_ram_64_512_delay1_inst_wen_to_strg_lifted,
  output logic valid_out_f_
);

strg_ram_64_512_delay1 strg_ram_64_512_delay1_inst (
  .clk(clk),
  .clk_en(clk_en),
  .data_from_strg(strg_ram_64_512_delay1_inst_data_from_strg_lifted),
  .data_in(data_in_f_),
  .flush(flush),
  .rd_addr_in(rd_addr_in_f_),
  .ren(ren_f_),
  .rst_n(rst_n),
  .wen(wen_f_),
  .wr_addr_in(wr_addr_in_f_),
  .addr_out(strg_ram_64_512_delay1_inst_addr_out_lifted),
  .data_out(data_out_f_),
  .data_to_strg(strg_ram_64_512_delay1_inst_data_to_strg_lifted),
  .ready(ready_f_),
  .ren_to_strg(strg_ram_64_512_delay1_inst_ren_to_strg_lifted),
  .valid_out(valid_out_f_),
  .wen_to_strg(strg_ram_64_512_delay1_inst_wen_to_strg_lifted)
);

endmodule   // strg_ram_64_512_delay1_flat

module strg_ub_agg_only (
  input logic [1:0] agg_read,
  input logic [2:0] agg_write_addr_gen_0_starting_addr,
  input logic [2:0] agg_write_addr_gen_0_strides_0,
  input logic [2:0] agg_write_addr_gen_0_strides_1,
  input logic [2:0] agg_write_addr_gen_0_strides_2,
  input logic [2:0] agg_write_addr_gen_1_starting_addr,
  input logic [2:0] agg_write_addr_gen_1_strides_0,
  input logic [2:0] agg_write_addr_gen_1_strides_1,
  input logic [2:0] agg_write_addr_gen_1_strides_2,
  input logic agg_write_sched_gen_0_enable,
  input logic [15:0] agg_write_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [15:0] agg_write_sched_gen_0_sched_addr_gen_strides_0,
  input logic [15:0] agg_write_sched_gen_0_sched_addr_gen_strides_1,
  input logic [15:0] agg_write_sched_gen_0_sched_addr_gen_strides_2,
  input logic agg_write_sched_gen_1_enable,
  input logic [15:0] agg_write_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [15:0] agg_write_sched_gen_1_sched_addr_gen_strides_0,
  input logic [15:0] agg_write_sched_gen_1_sched_addr_gen_strides_1,
  input logic [15:0] agg_write_sched_gen_1_sched_addr_gen_strides_2,
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic [1:0] [15:0] data_in,
  input logic flush,
  input logic [2:0] loops_in2buf_0_dimensionality,
  input logic [10:0] loops_in2buf_0_ranges_0,
  input logic [10:0] loops_in2buf_0_ranges_1,
  input logic [10:0] loops_in2buf_0_ranges_2,
  input logic [2:0] loops_in2buf_1_dimensionality,
  input logic [10:0] loops_in2buf_1_ranges_0,
  input logic [10:0] loops_in2buf_1_ranges_1,
  input logic [10:0] loops_in2buf_1_ranges_2,
  input logic rst_n,
  input logic [1:0] [8:0] sram_read_addr_in,
  input logic [1:0] [2:0] tb_read_addr_d_in,
  input logic [1:0] tb_read_d_in,
  input logic [1:0] [1:0] update_mode_in,
  output logic [1:0][3:0] [15:0] agg_data_out,
  output logic [1:0] [1:0] agg_write_addr_l2b_out,
  output logic [1:0] [2:0] agg_write_mux_sel_out,
  output logic [1:0] agg_write_out,
  output logic [1:0] agg_write_restart_out
);

logic [1:0][1:0][3:0][15:0] agg;
logic [1:0] agg_read_addr;
logic [1:0][7:0] agg_read_addr_gen_out;
logic [1:0] agg_read_addr_in;
logic [1:0] agg_write;
logic [1:0][2:0] agg_write_addr;
logic [2:0] agg_write_addr_gen_0_addr_out;
logic [2:0][2:0] agg_write_addr_gen_0_strides;
logic [2:0] agg_write_addr_gen_1_addr_out;
logic [2:0][2:0] agg_write_addr_gen_1_strides;
logic agg_write_sched_gen_0_valid_output;
logic agg_write_sched_gen_1_valid_output;
logic [2:0] fl_mux_sel_0;
logic [2:0] fl_mux_sel_1;
logic [1:0] loops_in2buf_0_mux_sel_out;
logic [2:0][10:0] loops_in2buf_0_ranges;
logic loops_in2buf_0_restart;
logic [1:0] loops_in2buf_1_mux_sel_out;
logic [2:0][10:0] loops_in2buf_1_ranges;
logic loops_in2buf_1_restart;
logic [1:0] mode_0;
logic [1:0] mode_1;
logic [2:0] tb_addr_0;
logic [2:0] tb_addr_1;
logic tb_read_0;
logic tb_read_1;
assign agg_write_out = agg_write;
assign mode_0 = update_mode_in[0];
assign agg_write_addr_l2b_out[0] = agg_write_addr[0][1:0];
assign tb_read_0 = mode_0[0] ? tb_read_d_in[1]: tb_read_d_in[0];
assign tb_addr_0 = mode_0[0] ? tb_read_addr_d_in[1]: tb_read_addr_d_in[0];
assign fl_mux_sel_0[1:0] = loops_in2buf_0_mux_sel_out;
assign fl_mux_sel_0[2] = 1'h0;
assign agg_write_mux_sel_out[0] = fl_mux_sel_0;
assign agg_write_restart_out[0] = loops_in2buf_0_restart;
assign agg_write_addr[0] = mode_0[1] ? tb_addr_0: agg_write_addr_gen_0_addr_out;
assign agg_write[0] = mode_0[1] ? tb_read_0: agg_write_sched_gen_0_valid_output;

always_ff @(posedge clk) begin
  if (clk_en) begin
    if (agg_write[0]) begin
      agg[0][agg_write_addr[0][2]][agg_write_addr[0][1:0]] <= data_in[0];
    end
  end
end
assign agg_read_addr_in[0] = sram_read_addr_in[0][0];
assign agg_read_addr_gen_out[0][0] = agg_read_addr_in[0];
assign agg_read_addr_gen_out[0][7:1] = 7'h0;
assign agg_read_addr[0] = agg_read_addr_gen_out[0][0];
always_comb begin
  agg_data_out[0] = agg[0][agg_read_addr[0]];
end
assign mode_1 = update_mode_in[1];
assign agg_write_addr_l2b_out[1] = agg_write_addr[1][1:0];
assign tb_read_1 = mode_1[0] ? tb_read_d_in[1]: tb_read_d_in[0];
assign tb_addr_1 = mode_1[0] ? tb_read_addr_d_in[1]: tb_read_addr_d_in[0];
assign fl_mux_sel_1[1:0] = loops_in2buf_1_mux_sel_out;
assign fl_mux_sel_1[2] = 1'h0;
assign agg_write_mux_sel_out[1] = fl_mux_sel_1;
assign agg_write_restart_out[1] = loops_in2buf_1_restart;
assign agg_write_addr[1] = mode_1[1] ? tb_addr_1: agg_write_addr_gen_1_addr_out;
assign agg_write[1] = mode_1[1] ? tb_read_1: agg_write_sched_gen_1_valid_output;

always_ff @(posedge clk) begin
  if (clk_en) begin
    if (agg_write[1]) begin
      agg[1][agg_write_addr[1][2]][agg_write_addr[1][1:0]] <= data_in[1];
    end
  end
end
assign agg_read_addr_in[1] = sram_read_addr_in[1][0];
assign agg_read_addr_gen_out[1][0] = agg_read_addr_in[1];
assign agg_read_addr_gen_out[1][7:1] = 7'h0;
assign agg_read_addr[1] = agg_read_addr_gen_out[1][0];
always_comb begin
  agg_data_out[1] = agg[1][agg_read_addr[1]];
end
assign loops_in2buf_0_ranges[0] = loops_in2buf_0_ranges_0;
assign loops_in2buf_0_ranges[1] = loops_in2buf_0_ranges_1;
assign loops_in2buf_0_ranges[2] = loops_in2buf_0_ranges_2;
assign agg_write_addr_gen_0_strides[0] = agg_write_addr_gen_0_strides_0;
assign agg_write_addr_gen_0_strides[1] = agg_write_addr_gen_0_strides_1;
assign agg_write_addr_gen_0_strides[2] = agg_write_addr_gen_0_strides_2;
assign loops_in2buf_1_ranges[0] = loops_in2buf_1_ranges_0;
assign loops_in2buf_1_ranges[1] = loops_in2buf_1_ranges_1;
assign loops_in2buf_1_ranges[2] = loops_in2buf_1_ranges_2;
assign agg_write_addr_gen_1_strides[0] = agg_write_addr_gen_1_strides_0;
assign agg_write_addr_gen_1_strides[1] = agg_write_addr_gen_1_strides_1;
assign agg_write_addr_gen_1_strides[2] = agg_write_addr_gen_1_strides_2;
for_loop_3_11 loops_in2buf_0 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_in2buf_0_dimensionality),
  .flush(flush),
  .ranges(loops_in2buf_0_ranges),
  .rst_n(rst_n),
  .step(agg_write[0]),
  .mux_sel_out(loops_in2buf_0_mux_sel_out),
  .restart(loops_in2buf_0_restart)
);

addr_gen_3_3 agg_write_addr_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(loops_in2buf_0_mux_sel_out),
  .restart(loops_in2buf_0_restart),
  .rst_n(rst_n),
  .starting_addr(agg_write_addr_gen_0_starting_addr),
  .step(agg_write[0]),
  .strides(agg_write_addr_gen_0_strides),
  .addr_out(agg_write_addr_gen_0_addr_out)
);

sched_gen_3_16 agg_write_sched_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(agg_write_sched_gen_0_enable),
  .finished(loops_in2buf_0_restart),
  .flush(flush),
  .mux_sel(loops_in2buf_0_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(agg_write_sched_gen_0_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides_0(agg_write_sched_gen_0_sched_addr_gen_strides_0),
  .sched_addr_gen_strides_1(agg_write_sched_gen_0_sched_addr_gen_strides_1),
  .sched_addr_gen_strides_2(agg_write_sched_gen_0_sched_addr_gen_strides_2),
  .valid_output(agg_write_sched_gen_0_valid_output)
);

for_loop_3_11 loops_in2buf_1 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_in2buf_1_dimensionality),
  .flush(flush),
  .ranges(loops_in2buf_1_ranges),
  .rst_n(rst_n),
  .step(agg_write[1]),
  .mux_sel_out(loops_in2buf_1_mux_sel_out),
  .restart(loops_in2buf_1_restart)
);

addr_gen_3_3 agg_write_addr_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(loops_in2buf_1_mux_sel_out),
  .restart(loops_in2buf_1_restart),
  .rst_n(rst_n),
  .starting_addr(agg_write_addr_gen_1_starting_addr),
  .step(agg_write[1]),
  .strides(agg_write_addr_gen_1_strides),
  .addr_out(agg_write_addr_gen_1_addr_out)
);

sched_gen_3_16 agg_write_sched_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(agg_write_sched_gen_1_enable),
  .finished(loops_in2buf_1_restart),
  .flush(flush),
  .mux_sel(loops_in2buf_1_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(agg_write_sched_gen_1_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides_0(agg_write_sched_gen_1_sched_addr_gen_strides_0),
  .sched_addr_gen_strides_1(agg_write_sched_gen_1_sched_addr_gen_strides_1),
  .sched_addr_gen_strides_2(agg_write_sched_gen_1_sched_addr_gen_strides_2),
  .valid_output(agg_write_sched_gen_1_valid_output)
);

endmodule   // strg_ub_agg_only

module strg_ub_agg_sram_shared (
  input logic [7:0] agg_read_sched_gen_0_agg_read_padding,
  input logic [7:0] agg_read_sched_gen_1_agg_read_padding,
  input logic [8:0] agg_sram_shared_addr_gen_0_starting_addr,
  input logic [8:0] agg_sram_shared_addr_gen_1_starting_addr,
  input logic [1:0] [1:0] agg_write_addr_l2b_in,
  input logic [1:0] agg_write_in,
  input logic [1:0] [2:0] agg_write_mux_sel_in,
  input logic [1:0] agg_write_restart_in,
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [1:0] mode_0,
  input logic [1:0] mode_1,
  input logic rst_n,
  input logic [1:0] [8:0] sram_read_addr_in,
  input logic [1:0] sram_read_d_in,
  input logic [1:0] sram_read_in,
  output logic [1:0] agg_read_out,
  output logic [1:0] [8:0] agg_sram_shared_addr_out,
  output logic [1:0] [1:0] update_mode_out
);

logic [1:0] agg_read;
logic agg_read_sched_gen_0_valid_output;
logic agg_read_sched_gen_1_valid_output;
logic [8:0] agg_sram_shared_addr_gen_0_addr_out;
logic [8:0] agg_sram_shared_addr_gen_1_addr_out;
assign agg_read_out = agg_read;
assign update_mode_out[0] = mode_0;
assign agg_read[0] = agg_read_sched_gen_0_valid_output;
assign agg_sram_shared_addr_out[0] = agg_sram_shared_addr_gen_0_addr_out;
assign update_mode_out[1] = mode_1;
assign agg_read[1] = agg_read_sched_gen_1_valid_output;
assign agg_sram_shared_addr_out[1] = agg_sram_shared_addr_gen_1_addr_out;
agg_sram_shared_sched_gen agg_read_sched_gen_0 (
  .agg_read_padding(agg_read_sched_gen_0_agg_read_padding),
  .agg_write(agg_write_in[0]),
  .agg_write_addr_l2b(agg_write_addr_l2b_in[0]),
  .agg_write_mux_sel(agg_write_mux_sel_in[0]),
  .agg_write_restart(agg_write_restart_in[0]),
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mode(mode_0),
  .rst_n(rst_n),
  .sram_read_d(sram_read_d_in),
  .valid_output(agg_read_sched_gen_0_valid_output)
);

agg_sram_shared_addr_gen agg_sram_shared_addr_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mode(mode_0),
  .rst_n(rst_n),
  .sram_read(sram_read_in),
  .sram_read_addr(sram_read_addr_in),
  .starting_addr(agg_sram_shared_addr_gen_0_starting_addr),
  .step(agg_read[0]),
  .addr_out(agg_sram_shared_addr_gen_0_addr_out)
);

agg_sram_shared_sched_gen agg_read_sched_gen_1 (
  .agg_read_padding(agg_read_sched_gen_1_agg_read_padding),
  .agg_write(agg_write_in[1]),
  .agg_write_addr_l2b(agg_write_addr_l2b_in[1]),
  .agg_write_mux_sel(agg_write_mux_sel_in[1]),
  .agg_write_restart(agg_write_restart_in[1]),
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mode(mode_1),
  .rst_n(rst_n),
  .sram_read_d(sram_read_d_in),
  .valid_output(agg_read_sched_gen_1_valid_output)
);

agg_sram_shared_addr_gen agg_sram_shared_addr_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mode(mode_1),
  .rst_n(rst_n),
  .sram_read(sram_read_in),
  .sram_read_addr(sram_read_addr_in),
  .starting_addr(agg_sram_shared_addr_gen_1_starting_addr),
  .step(agg_read[1]),
  .addr_out(agg_sram_shared_addr_gen_1_addr_out)
);

endmodule   // strg_ub_agg_sram_shared

module strg_ub_sram_only (
  input logic [1:0][3:0] [15:0] agg_data_out,
  input logic [1:0] agg_read,
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic flush,
  input logic [1:0] [2:0] loops_sram2tb_mux_sel,
  input logic [1:0] loops_sram2tb_restart,
  input logic [8:0] output_addr_gen_0_starting_addr,
  input logic [8:0] output_addr_gen_0_strides_0,
  input logic [8:0] output_addr_gen_0_strides_1,
  input logic [8:0] output_addr_gen_0_strides_2,
  input logic [8:0] output_addr_gen_0_strides_3,
  input logic [8:0] output_addr_gen_0_strides_4,
  input logic [8:0] output_addr_gen_0_strides_5,
  input logic [8:0] output_addr_gen_1_starting_addr,
  input logic [8:0] output_addr_gen_1_strides_0,
  input logic [8:0] output_addr_gen_1_strides_1,
  input logic [8:0] output_addr_gen_1_strides_2,
  input logic [8:0] output_addr_gen_1_strides_3,
  input logic [8:0] output_addr_gen_1_strides_4,
  input logic [8:0] output_addr_gen_1_strides_5,
  input logic rst_n,
  input logic [1:0] [8:0] sram_read_addr_in,
  input logic [1:0] t_read,
  output logic [8:0] addr_to_sram,
  output logic cen_to_sram,
  output logic [3:0] [15:0] data_to_sram,
  output logic [1:0] [8:0] sram_read_addr_out,
  output logic wen_to_sram
);

logic [8:0] addr;
logic [3:0][15:0] decode_ret_agg_read_agg_data_out;
logic [15:0] decode_ret_agg_read_s_write_addr;
logic [15:0] decode_ret_t_read_s_read_addr;
logic decode_sel_done_agg_read_agg_data_out;
logic decode_sel_done_agg_read_s_write_addr;
logic decode_sel_done_t_read_s_read_addr;
logic [8:0] output_addr_gen_0_addr_out;
logic [5:0][8:0] output_addr_gen_0_strides;
logic [8:0] output_addr_gen_1_addr_out;
logic [5:0][8:0] output_addr_gen_1_strides;
logic read;
logic [1:0][15:0] s_read_addr;
logic [1:0][15:0] s_write_addr;
logic [3:0][15:0] sram_write_data;
logic write;
assign s_write_addr[0][8:0] = sram_read_addr_in[0];
assign s_write_addr[0][15:9] = 7'h0;
assign s_write_addr[1][8:0] = sram_read_addr_in[1];
assign s_write_addr[1][15:9] = 7'h0;
assign s_read_addr[0][8:0] = output_addr_gen_0_addr_out;
assign s_read_addr[0][15:9] = 7'h0;
assign sram_read_addr_out[0] = output_addr_gen_0_addr_out;
assign s_read_addr[1][8:0] = output_addr_gen_1_addr_out;
assign s_read_addr[1][15:9] = 7'h0;
assign sram_read_addr_out[1] = output_addr_gen_1_addr_out;
assign data_to_sram = sram_write_data;
assign wen_to_sram = write;
always_comb begin
  decode_sel_done_agg_read_s_write_addr = 1'h0;
  decode_ret_agg_read_s_write_addr = 16'h0;
  for (int unsigned i = 0; i < 2; i += 1) begin
      if ((~decode_sel_done_agg_read_s_write_addr) & agg_read[1'(i)]) begin
        decode_ret_agg_read_s_write_addr = s_write_addr[1'(i)];
        decode_sel_done_agg_read_s_write_addr = 1'h1;
      end
    end
end
always_comb begin
  decode_sel_done_t_read_s_read_addr = 1'h0;
  decode_ret_t_read_s_read_addr = 16'h0;
  for (int unsigned i = 0; i < 2; i += 1) begin
      if ((~decode_sel_done_t_read_s_read_addr) & t_read[1'(i)]) begin
        decode_ret_t_read_s_read_addr = s_read_addr[1'(i)];
        decode_sel_done_t_read_s_read_addr = 1'h1;
      end
    end
end
assign cen_to_sram = write | read;
assign addr_to_sram = addr;
always_comb begin
  if (write) begin
    addr = decode_ret_agg_read_s_write_addr[8:0];
  end
  else addr = decode_ret_t_read_s_read_addr[8:0];
end
assign write = |agg_read;
assign read = |t_read;
always_comb begin
  decode_sel_done_agg_read_agg_data_out = 1'h0;
  decode_ret_agg_read_agg_data_out = 64'h0;
  for (int unsigned i = 0; i < 2; i += 1) begin
      if ((~decode_sel_done_agg_read_agg_data_out) & agg_read[1'(i)]) begin
        decode_ret_agg_read_agg_data_out = agg_data_out[1'(i)];
        decode_sel_done_agg_read_agg_data_out = 1'h1;
      end
    end
end
assign sram_write_data = decode_ret_agg_read_agg_data_out;
assign output_addr_gen_0_strides[0] = output_addr_gen_0_strides_0;
assign output_addr_gen_0_strides[1] = output_addr_gen_0_strides_1;
assign output_addr_gen_0_strides[2] = output_addr_gen_0_strides_2;
assign output_addr_gen_0_strides[3] = output_addr_gen_0_strides_3;
assign output_addr_gen_0_strides[4] = output_addr_gen_0_strides_4;
assign output_addr_gen_0_strides[5] = output_addr_gen_0_strides_5;
assign output_addr_gen_1_strides[0] = output_addr_gen_1_strides_0;
assign output_addr_gen_1_strides[1] = output_addr_gen_1_strides_1;
assign output_addr_gen_1_strides[2] = output_addr_gen_1_strides_2;
assign output_addr_gen_1_strides[3] = output_addr_gen_1_strides_3;
assign output_addr_gen_1_strides[4] = output_addr_gen_1_strides_4;
assign output_addr_gen_1_strides[5] = output_addr_gen_1_strides_5;
addr_gen_6_9 output_addr_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(loops_sram2tb_mux_sel[0]),
  .restart(loops_sram2tb_restart[0]),
  .rst_n(rst_n),
  .starting_addr(output_addr_gen_0_starting_addr),
  .step(t_read[0]),
  .strides(output_addr_gen_0_strides),
  .addr_out(output_addr_gen_0_addr_out)
);

addr_gen_6_9 output_addr_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(loops_sram2tb_mux_sel[1]),
  .restart(loops_sram2tb_restart[1]),
  .rst_n(rst_n),
  .starting_addr(output_addr_gen_1_starting_addr),
  .step(t_read[1]),
  .strides(output_addr_gen_1_strides),
  .addr_out(output_addr_gen_1_addr_out)
);

endmodule   // strg_ub_sram_only

module strg_ub_sram_tb_shared (
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic flush,
  input logic [3:0] loops_buf2out_autovec_read_0_dimensionality,
  input logic [10:0] loops_buf2out_autovec_read_0_ranges_0,
  input logic [10:0] loops_buf2out_autovec_read_0_ranges_1,
  input logic [10:0] loops_buf2out_autovec_read_0_ranges_2,
  input logic [10:0] loops_buf2out_autovec_read_0_ranges_3,
  input logic [10:0] loops_buf2out_autovec_read_0_ranges_4,
  input logic [10:0] loops_buf2out_autovec_read_0_ranges_5,
  input logic [3:0] loops_buf2out_autovec_read_1_dimensionality,
  input logic [10:0] loops_buf2out_autovec_read_1_ranges_0,
  input logic [10:0] loops_buf2out_autovec_read_1_ranges_1,
  input logic [10:0] loops_buf2out_autovec_read_1_ranges_2,
  input logic [10:0] loops_buf2out_autovec_read_1_ranges_3,
  input logic [10:0] loops_buf2out_autovec_read_1_ranges_4,
  input logic [10:0] loops_buf2out_autovec_read_1_ranges_5,
  input logic output_sched_gen_0_enable,
  input logic [9:0] output_sched_gen_0_sched_addr_gen_delay,
  input logic [15:0] output_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [15:0] output_sched_gen_0_sched_addr_gen_strides_0,
  input logic [15:0] output_sched_gen_0_sched_addr_gen_strides_1,
  input logic [15:0] output_sched_gen_0_sched_addr_gen_strides_2,
  input logic [15:0] output_sched_gen_0_sched_addr_gen_strides_3,
  input logic [15:0] output_sched_gen_0_sched_addr_gen_strides_4,
  input logic [15:0] output_sched_gen_0_sched_addr_gen_strides_5,
  input logic output_sched_gen_1_enable,
  input logic [9:0] output_sched_gen_1_sched_addr_gen_delay,
  input logic [15:0] output_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [15:0] output_sched_gen_1_sched_addr_gen_strides_0,
  input logic [15:0] output_sched_gen_1_sched_addr_gen_strides_1,
  input logic [15:0] output_sched_gen_1_sched_addr_gen_strides_2,
  input logic [15:0] output_sched_gen_1_sched_addr_gen_strides_3,
  input logic [15:0] output_sched_gen_1_sched_addr_gen_strides_4,
  input logic [15:0] output_sched_gen_1_sched_addr_gen_strides_5,
  input logic rst_n,
  output logic [1:0] [2:0] loops_sram2tb_mux_sel,
  output logic [1:0] loops_sram2tb_restart,
  output logic [1:0] sram_read_d,
  output logic [1:0] t_read_out
);

logic [2:0] loops_buf2out_autovec_read_0_mux_sel_out;
logic [5:0][10:0] loops_buf2out_autovec_read_0_ranges;
logic loops_buf2out_autovec_read_0_restart;
logic [2:0] loops_buf2out_autovec_read_1_mux_sel_out;
logic [5:0][10:0] loops_buf2out_autovec_read_1_ranges;
logic loops_buf2out_autovec_read_1_restart;
logic output_sched_gen_0_valid_output;
logic output_sched_gen_0_valid_output_d;
logic output_sched_gen_1_valid_output;
logic output_sched_gen_1_valid_output_d;
logic [1:0] t_read;
assign t_read_out = t_read;
assign loops_sram2tb_mux_sel[0] = loops_buf2out_autovec_read_0_mux_sel_out;
assign loops_sram2tb_restart[0] = loops_buf2out_autovec_read_0_restart;
assign t_read[0] = output_sched_gen_0_valid_output;
assign sram_read_d[0] = output_sched_gen_0_valid_output_d;
assign loops_sram2tb_mux_sel[1] = loops_buf2out_autovec_read_1_mux_sel_out;
assign loops_sram2tb_restart[1] = loops_buf2out_autovec_read_1_restart;
assign t_read[1] = output_sched_gen_1_valid_output;
assign sram_read_d[1] = output_sched_gen_1_valid_output_d;
assign loops_buf2out_autovec_read_0_ranges[0] = loops_buf2out_autovec_read_0_ranges_0;
assign loops_buf2out_autovec_read_0_ranges[1] = loops_buf2out_autovec_read_0_ranges_1;
assign loops_buf2out_autovec_read_0_ranges[2] = loops_buf2out_autovec_read_0_ranges_2;
assign loops_buf2out_autovec_read_0_ranges[3] = loops_buf2out_autovec_read_0_ranges_3;
assign loops_buf2out_autovec_read_0_ranges[4] = loops_buf2out_autovec_read_0_ranges_4;
assign loops_buf2out_autovec_read_0_ranges[5] = loops_buf2out_autovec_read_0_ranges_5;
assign loops_buf2out_autovec_read_1_ranges[0] = loops_buf2out_autovec_read_1_ranges_0;
assign loops_buf2out_autovec_read_1_ranges[1] = loops_buf2out_autovec_read_1_ranges_1;
assign loops_buf2out_autovec_read_1_ranges[2] = loops_buf2out_autovec_read_1_ranges_2;
assign loops_buf2out_autovec_read_1_ranges[3] = loops_buf2out_autovec_read_1_ranges_3;
assign loops_buf2out_autovec_read_1_ranges[4] = loops_buf2out_autovec_read_1_ranges_4;
assign loops_buf2out_autovec_read_1_ranges[5] = loops_buf2out_autovec_read_1_ranges_5;
for_loop_6_11 loops_buf2out_autovec_read_0 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_buf2out_autovec_read_0_dimensionality),
  .flush(flush),
  .ranges(loops_buf2out_autovec_read_0_ranges),
  .rst_n(rst_n),
  .step(t_read[0]),
  .mux_sel_out(loops_buf2out_autovec_read_0_mux_sel_out),
  .restart(loops_buf2out_autovec_read_0_restart)
);

sched_gen_6_16_delay_addr_10_4 output_sched_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(output_sched_gen_0_enable),
  .finished(loops_buf2out_autovec_read_0_restart),
  .flush(flush),
  .mux_sel(loops_buf2out_autovec_read_0_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_delay(output_sched_gen_0_sched_addr_gen_delay),
  .sched_addr_gen_starting_addr(output_sched_gen_0_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides_0(output_sched_gen_0_sched_addr_gen_strides_0),
  .sched_addr_gen_strides_1(output_sched_gen_0_sched_addr_gen_strides_1),
  .sched_addr_gen_strides_2(output_sched_gen_0_sched_addr_gen_strides_2),
  .sched_addr_gen_strides_3(output_sched_gen_0_sched_addr_gen_strides_3),
  .sched_addr_gen_strides_4(output_sched_gen_0_sched_addr_gen_strides_4),
  .sched_addr_gen_strides_5(output_sched_gen_0_sched_addr_gen_strides_5),
  .valid_output(output_sched_gen_0_valid_output),
  .valid_output_d(output_sched_gen_0_valid_output_d)
);

for_loop_6_11 loops_buf2out_autovec_read_1 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_buf2out_autovec_read_1_dimensionality),
  .flush(flush),
  .ranges(loops_buf2out_autovec_read_1_ranges),
  .rst_n(rst_n),
  .step(t_read[1]),
  .mux_sel_out(loops_buf2out_autovec_read_1_mux_sel_out),
  .restart(loops_buf2out_autovec_read_1_restart)
);

sched_gen_6_16_delay_addr_10_4 output_sched_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(output_sched_gen_1_enable),
  .finished(loops_buf2out_autovec_read_1_restart),
  .flush(flush),
  .mux_sel(loops_buf2out_autovec_read_1_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_delay(output_sched_gen_1_sched_addr_gen_delay),
  .sched_addr_gen_starting_addr(output_sched_gen_1_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides_0(output_sched_gen_1_sched_addr_gen_strides_0),
  .sched_addr_gen_strides_1(output_sched_gen_1_sched_addr_gen_strides_1),
  .sched_addr_gen_strides_2(output_sched_gen_1_sched_addr_gen_strides_2),
  .sched_addr_gen_strides_3(output_sched_gen_1_sched_addr_gen_strides_3),
  .sched_addr_gen_strides_4(output_sched_gen_1_sched_addr_gen_strides_4),
  .sched_addr_gen_strides_5(output_sched_gen_1_sched_addr_gen_strides_5),
  .valid_output(output_sched_gen_1_valid_output),
  .valid_output_d(output_sched_gen_1_valid_output_d)
);

endmodule   // strg_ub_sram_tb_shared

module strg_ub_tb_only (
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic flush,
  input logic [3:0] loops_buf2out_read_0_dimensionality,
  input logic [10:0] loops_buf2out_read_0_ranges_0,
  input logic [10:0] loops_buf2out_read_0_ranges_1,
  input logic [10:0] loops_buf2out_read_0_ranges_2,
  input logic [10:0] loops_buf2out_read_0_ranges_3,
  input logic [10:0] loops_buf2out_read_0_ranges_4,
  input logic [10:0] loops_buf2out_read_0_ranges_5,
  input logic [3:0] loops_buf2out_read_1_dimensionality,
  input logic [10:0] loops_buf2out_read_1_ranges_0,
  input logic [10:0] loops_buf2out_read_1_ranges_1,
  input logic [10:0] loops_buf2out_read_1_ranges_2,
  input logic [10:0] loops_buf2out_read_1_ranges_3,
  input logic [10:0] loops_buf2out_read_1_ranges_4,
  input logic [10:0] loops_buf2out_read_1_ranges_5,
  input logic [1:0] [2:0] loops_sram2tb_mux_sel,
  input logic [1:0] loops_sram2tb_restart,
  input logic rst_n,
  input logic shared_tb_0,
  input logic [3:0] [15:0] sram_read_data,
  input logic [1:0] t_read,
  input logic [3:0] tb_read_addr_gen_0_starting_addr,
  input logic [3:0] tb_read_addr_gen_0_strides_0,
  input logic [3:0] tb_read_addr_gen_0_strides_1,
  input logic [3:0] tb_read_addr_gen_0_strides_2,
  input logic [3:0] tb_read_addr_gen_0_strides_3,
  input logic [3:0] tb_read_addr_gen_0_strides_4,
  input logic [3:0] tb_read_addr_gen_0_strides_5,
  input logic [3:0] tb_read_addr_gen_1_starting_addr,
  input logic [3:0] tb_read_addr_gen_1_strides_0,
  input logic [3:0] tb_read_addr_gen_1_strides_1,
  input logic [3:0] tb_read_addr_gen_1_strides_2,
  input logic [3:0] tb_read_addr_gen_1_strides_3,
  input logic [3:0] tb_read_addr_gen_1_strides_4,
  input logic [3:0] tb_read_addr_gen_1_strides_5,
  input logic tb_read_sched_gen_0_enable,
  input logic [9:0] tb_read_sched_gen_0_sched_addr_gen_delay,
  input logic [15:0] tb_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [15:0] tb_read_sched_gen_0_sched_addr_gen_strides_0,
  input logic [15:0] tb_read_sched_gen_0_sched_addr_gen_strides_1,
  input logic [15:0] tb_read_sched_gen_0_sched_addr_gen_strides_2,
  input logic [15:0] tb_read_sched_gen_0_sched_addr_gen_strides_3,
  input logic [15:0] tb_read_sched_gen_0_sched_addr_gen_strides_4,
  input logic [15:0] tb_read_sched_gen_0_sched_addr_gen_strides_5,
  input logic tb_read_sched_gen_1_enable,
  input logic [9:0] tb_read_sched_gen_1_sched_addr_gen_delay,
  input logic [15:0] tb_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [15:0] tb_read_sched_gen_1_sched_addr_gen_strides_0,
  input logic [15:0] tb_read_sched_gen_1_sched_addr_gen_strides_1,
  input logic [15:0] tb_read_sched_gen_1_sched_addr_gen_strides_2,
  input logic [15:0] tb_read_sched_gen_1_sched_addr_gen_strides_3,
  input logic [15:0] tb_read_sched_gen_1_sched_addr_gen_strides_4,
  input logic [15:0] tb_read_sched_gen_1_sched_addr_gen_strides_5,
  input logic [3:0] tb_write_addr_gen_0_starting_addr,
  input logic [3:0] tb_write_addr_gen_0_strides_0,
  input logic [3:0] tb_write_addr_gen_0_strides_1,
  input logic [3:0] tb_write_addr_gen_0_strides_2,
  input logic [3:0] tb_write_addr_gen_0_strides_3,
  input logic [3:0] tb_write_addr_gen_0_strides_4,
  input logic [3:0] tb_write_addr_gen_0_strides_5,
  input logic [3:0] tb_write_addr_gen_1_starting_addr,
  input logic [3:0] tb_write_addr_gen_1_strides_0,
  input logic [3:0] tb_write_addr_gen_1_strides_1,
  input logic [3:0] tb_write_addr_gen_1_strides_2,
  input logic [3:0] tb_write_addr_gen_1_strides_3,
  input logic [3:0] tb_write_addr_gen_1_strides_4,
  input logic [3:0] tb_write_addr_gen_1_strides_5,
  output logic [1:0] accessor_output,
  output logic [1:0] [15:0] data_out,
  output logic [1:0] [2:0] tb_read_addr_d_out,
  output logic [1:0] tb_read_d_out
);

logic [2:0] addr_fifo_in_0;
logic [2:0] addr_fifo_in_1;
logic delay_en_0;
logic delay_en_1;
logic [2:0] loops_buf2out_read_0_mux_sel_out;
logic [5:0][10:0] loops_buf2out_read_0_ranges;
logic loops_buf2out_read_0_restart;
logic [2:0] loops_buf2out_read_1_mux_sel_out;
logic [5:0][10:0] loops_buf2out_read_1_ranges;
logic loops_buf2out_read_1_restart;
logic [1:0][2:0] mux_sel_d1;
logic [2:0] rd_ptr_0;
logic [2:0] rd_ptr_1;
logic [1:0] restart_d1;
logic [1:0] t_read_d1;
logic [1:0][1:0][3:0][15:0] tb;
logic [7:0][2:0] tb_addr_fifo_0;
logic [7:0][2:0] tb_addr_fifo_1;
logic [1:0] tb_read;
logic [1:0][3:0] tb_read_addr;
logic [3:0] tb_read_addr_gen_0_addr_out;
logic [5:0][3:0] tb_read_addr_gen_0_strides;
logic [3:0] tb_read_addr_gen_1_addr_out;
logic [5:0][3:0] tb_read_addr_gen_1_strides;
logic tb_read_d_0;
logic tb_read_d_1;
logic tb_read_sched_gen_0_valid_output;
logic tb_read_sched_gen_1_valid_output;
logic tb_read_sel_0;
logic [1:0][2:0] tb_write_addr;
logic [3:0] tb_write_addr_gen_0_addr_out;
logic [5:0][3:0] tb_write_addr_gen_0_strides;
logic [3:0] tb_write_addr_gen_1_addr_out;
logic [5:0][3:0] tb_write_addr_gen_1_strides;
logic tb_write_sel_0;
logic [2:0] wr_ptr_0;
logic [2:0] wr_ptr_1;
assign accessor_output = tb_read;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    t_read_d1[0] <= 1'h0;
    mux_sel_d1[0] <= 3'h0;
    restart_d1[0] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      t_read_d1[0] <= 1'h0;
      mux_sel_d1[0] <= 3'h0;
      restart_d1[0] <= 1'h0;
    end
    else begin
      t_read_d1[0] <= t_read[0];
      mux_sel_d1[0] <= loops_sram2tb_mux_sel[0];
      restart_d1[0] <= loops_sram2tb_restart[0];
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    t_read_d1[1] <= 1'h0;
    mux_sel_d1[1] <= 3'h0;
    restart_d1[1] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      t_read_d1[1] <= 1'h0;
      mux_sel_d1[1] <= 3'h0;
      restart_d1[1] <= 1'h0;
    end
    else begin
      t_read_d1[1] <= t_read[1];
      mux_sel_d1[1] <= loops_sram2tb_mux_sel[1];
      restart_d1[1] <= loops_sram2tb_restart[1];
    end
  end
end
assign tb_write_sel_0 = shared_tb_0 ? tb_write_addr[0][1]: 1'h0;
assign tb_read_sel_0 = shared_tb_0 ? tb_read_addr[0][3]: 1'h0;
assign tb_write_addr[0] = tb_write_addr_gen_0_addr_out[2:0];
assign tb_read_addr[0] = tb_read_addr_gen_0_addr_out;
assign tb_read[0] = tb_read_sched_gen_0_valid_output;
assign addr_fifo_in_0 = tb_read_addr_gen_0_addr_out[2:0];

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    wr_ptr_0 <= 3'h0;
    rd_ptr_0 <= 3'h0;
    tb_addr_fifo_0 <= 24'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      wr_ptr_0 <= 3'h0;
      rd_ptr_0 <= 3'h0;
      tb_addr_fifo_0 <= 24'h0;
    end
    else if (delay_en_0) begin
      if (tb_read[0]) begin
        tb_addr_fifo_0[wr_ptr_0] <= addr_fifo_in_0;
        wr_ptr_0 <= wr_ptr_0 + 3'h1;
      end
      if (tb_read_d_0) begin
        rd_ptr_0 <= rd_ptr_0 + 3'h1;
      end
    end
  end
end
assign tb_read_d_out[0] = delay_en_0 ? tb_read_d_0: tb_read[0];
assign tb_read_addr_d_out[0] = delay_en_0 ? tb_addr_fifo_0[rd_ptr_0]: addr_fifo_in_0;
always_comb begin
  data_out[0] = tb[tb_read_sel_0][tb_read_addr[0][2]][tb_read_addr[0][1:0]];
end
assign tb_write_addr[1] = tb_write_addr_gen_1_addr_out[2:0];
assign tb_read_addr[1] = tb_read_addr_gen_1_addr_out;
assign tb_read[1] = tb_read_sched_gen_1_valid_output;
assign addr_fifo_in_1 = tb_read_addr_gen_1_addr_out[2:0];

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    wr_ptr_1 <= 3'h0;
    rd_ptr_1 <= 3'h0;
    tb_addr_fifo_1 <= 24'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      wr_ptr_1 <= 3'h0;
      rd_ptr_1 <= 3'h0;
      tb_addr_fifo_1 <= 24'h0;
    end
    else if (delay_en_1) begin
      if (tb_read[1]) begin
        tb_addr_fifo_1[wr_ptr_1] <= addr_fifo_in_1;
        wr_ptr_1 <= wr_ptr_1 + 3'h1;
      end
      if (tb_read_d_1) begin
        rd_ptr_1 <= rd_ptr_1 + 3'h1;
      end
    end
  end
end
assign tb_read_d_out[1] = delay_en_1 ? tb_read_d_1: tb_read[1];
assign tb_read_addr_d_out[1] = delay_en_1 ? tb_addr_fifo_1[rd_ptr_1]: addr_fifo_in_1;
always_comb begin
  data_out[1] = tb[1][tb_read_addr[1][2]][tb_read_addr[1][1:0]];
end

always_ff @(posedge clk) begin
  if (clk_en) begin
    for (int unsigned i = 0; i < 2; i += 1) begin
        if (t_read_d1[1'(i)]) begin
          if (i == 32'h0) begin
            tb[tb_write_sel_0][tb_write_addr[1'(i)][0]] <= sram_read_data;
          end
          else tb[1'(i)][tb_write_addr[1'(i)][0]] <= sram_read_data;
        end
      end
  end
end
assign tb_write_addr_gen_0_strides[0] = tb_write_addr_gen_0_strides_0;
assign tb_write_addr_gen_0_strides[1] = tb_write_addr_gen_0_strides_1;
assign tb_write_addr_gen_0_strides[2] = tb_write_addr_gen_0_strides_2;
assign tb_write_addr_gen_0_strides[3] = tb_write_addr_gen_0_strides_3;
assign tb_write_addr_gen_0_strides[4] = tb_write_addr_gen_0_strides_4;
assign tb_write_addr_gen_0_strides[5] = tb_write_addr_gen_0_strides_5;
assign loops_buf2out_read_0_ranges[0] = loops_buf2out_read_0_ranges_0;
assign loops_buf2out_read_0_ranges[1] = loops_buf2out_read_0_ranges_1;
assign loops_buf2out_read_0_ranges[2] = loops_buf2out_read_0_ranges_2;
assign loops_buf2out_read_0_ranges[3] = loops_buf2out_read_0_ranges_3;
assign loops_buf2out_read_0_ranges[4] = loops_buf2out_read_0_ranges_4;
assign loops_buf2out_read_0_ranges[5] = loops_buf2out_read_0_ranges_5;
assign tb_read_addr_gen_0_strides[0] = tb_read_addr_gen_0_strides_0;
assign tb_read_addr_gen_0_strides[1] = tb_read_addr_gen_0_strides_1;
assign tb_read_addr_gen_0_strides[2] = tb_read_addr_gen_0_strides_2;
assign tb_read_addr_gen_0_strides[3] = tb_read_addr_gen_0_strides_3;
assign tb_read_addr_gen_0_strides[4] = tb_read_addr_gen_0_strides_4;
assign tb_read_addr_gen_0_strides[5] = tb_read_addr_gen_0_strides_5;
assign tb_write_addr_gen_1_strides[0] = tb_write_addr_gen_1_strides_0;
assign tb_write_addr_gen_1_strides[1] = tb_write_addr_gen_1_strides_1;
assign tb_write_addr_gen_1_strides[2] = tb_write_addr_gen_1_strides_2;
assign tb_write_addr_gen_1_strides[3] = tb_write_addr_gen_1_strides_3;
assign tb_write_addr_gen_1_strides[4] = tb_write_addr_gen_1_strides_4;
assign tb_write_addr_gen_1_strides[5] = tb_write_addr_gen_1_strides_5;
assign loops_buf2out_read_1_ranges[0] = loops_buf2out_read_1_ranges_0;
assign loops_buf2out_read_1_ranges[1] = loops_buf2out_read_1_ranges_1;
assign loops_buf2out_read_1_ranges[2] = loops_buf2out_read_1_ranges_2;
assign loops_buf2out_read_1_ranges[3] = loops_buf2out_read_1_ranges_3;
assign loops_buf2out_read_1_ranges[4] = loops_buf2out_read_1_ranges_4;
assign loops_buf2out_read_1_ranges[5] = loops_buf2out_read_1_ranges_5;
assign tb_read_addr_gen_1_strides[0] = tb_read_addr_gen_1_strides_0;
assign tb_read_addr_gen_1_strides[1] = tb_read_addr_gen_1_strides_1;
assign tb_read_addr_gen_1_strides[2] = tb_read_addr_gen_1_strides_2;
assign tb_read_addr_gen_1_strides[3] = tb_read_addr_gen_1_strides_3;
assign tb_read_addr_gen_1_strides[4] = tb_read_addr_gen_1_strides_4;
assign tb_read_addr_gen_1_strides[5] = tb_read_addr_gen_1_strides_5;
addr_gen_6_4 tb_write_addr_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(mux_sel_d1[0]),
  .restart(restart_d1[0]),
  .rst_n(rst_n),
  .starting_addr(tb_write_addr_gen_0_starting_addr),
  .step(t_read_d1[0]),
  .strides(tb_write_addr_gen_0_strides),
  .addr_out(tb_write_addr_gen_0_addr_out)
);

for_loop_6_11 loops_buf2out_read_0 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_buf2out_read_0_dimensionality),
  .flush(flush),
  .ranges(loops_buf2out_read_0_ranges),
  .rst_n(rst_n),
  .step(tb_read[0]),
  .mux_sel_out(loops_buf2out_read_0_mux_sel_out),
  .restart(loops_buf2out_read_0_restart)
);

addr_gen_6_4 tb_read_addr_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(loops_buf2out_read_0_mux_sel_out),
  .restart(loops_buf2out_read_0_restart),
  .rst_n(rst_n),
  .starting_addr(tb_read_addr_gen_0_starting_addr),
  .step(tb_read[0]),
  .strides(tb_read_addr_gen_0_strides),
  .addr_out(tb_read_addr_gen_0_addr_out)
);

sched_gen_6_16_delay_addr_10_8 tb_read_sched_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(tb_read_sched_gen_0_enable),
  .finished(loops_buf2out_read_0_restart),
  .flush(flush),
  .mux_sel(loops_buf2out_read_0_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_delay(tb_read_sched_gen_0_sched_addr_gen_delay),
  .sched_addr_gen_starting_addr(tb_read_sched_gen_0_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides_0(tb_read_sched_gen_0_sched_addr_gen_strides_0),
  .sched_addr_gen_strides_1(tb_read_sched_gen_0_sched_addr_gen_strides_1),
  .sched_addr_gen_strides_2(tb_read_sched_gen_0_sched_addr_gen_strides_2),
  .sched_addr_gen_strides_3(tb_read_sched_gen_0_sched_addr_gen_strides_3),
  .sched_addr_gen_strides_4(tb_read_sched_gen_0_sched_addr_gen_strides_4),
  .sched_addr_gen_strides_5(tb_read_sched_gen_0_sched_addr_gen_strides_5),
  .delay_en_out(delay_en_0),
  .valid_output(tb_read_sched_gen_0_valid_output),
  .valid_output_d(tb_read_d_0)
);

addr_gen_6_4 tb_write_addr_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(mux_sel_d1[1]),
  .restart(restart_d1[1]),
  .rst_n(rst_n),
  .starting_addr(tb_write_addr_gen_1_starting_addr),
  .step(t_read_d1[1]),
  .strides(tb_write_addr_gen_1_strides),
  .addr_out(tb_write_addr_gen_1_addr_out)
);

for_loop_6_11 loops_buf2out_read_1 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_buf2out_read_1_dimensionality),
  .flush(flush),
  .ranges(loops_buf2out_read_1_ranges),
  .rst_n(rst_n),
  .step(tb_read[1]),
  .mux_sel_out(loops_buf2out_read_1_mux_sel_out),
  .restart(loops_buf2out_read_1_restart)
);

addr_gen_6_4 tb_read_addr_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(loops_buf2out_read_1_mux_sel_out),
  .restart(loops_buf2out_read_1_restart),
  .rst_n(rst_n),
  .starting_addr(tb_read_addr_gen_1_starting_addr),
  .step(tb_read[1]),
  .strides(tb_read_addr_gen_1_strides),
  .addr_out(tb_read_addr_gen_1_addr_out)
);

sched_gen_6_16_delay_addr_10_8 tb_read_sched_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(tb_read_sched_gen_1_enable),
  .finished(loops_buf2out_read_1_restart),
  .flush(flush),
  .mux_sel(loops_buf2out_read_1_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_delay(tb_read_sched_gen_1_sched_addr_gen_delay),
  .sched_addr_gen_starting_addr(tb_read_sched_gen_1_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides_0(tb_read_sched_gen_1_sched_addr_gen_strides_0),
  .sched_addr_gen_strides_1(tb_read_sched_gen_1_sched_addr_gen_strides_1),
  .sched_addr_gen_strides_2(tb_read_sched_gen_1_sched_addr_gen_strides_2),
  .sched_addr_gen_strides_3(tb_read_sched_gen_1_sched_addr_gen_strides_3),
  .sched_addr_gen_strides_4(tb_read_sched_gen_1_sched_addr_gen_strides_4),
  .sched_addr_gen_strides_5(tb_read_sched_gen_1_sched_addr_gen_strides_5),
  .delay_en_out(delay_en_1),
  .valid_output(tb_read_sched_gen_1_valid_output),
  .valid_output_d(tb_read_d_1)
);

endmodule   // strg_ub_tb_only

module strg_ub_vec (
  input logic [2:0] agg_only_agg_write_addr_gen_0_starting_addr,
  input logic [2:0] agg_only_agg_write_addr_gen_0_strides_0,
  input logic [2:0] agg_only_agg_write_addr_gen_0_strides_1,
  input logic [2:0] agg_only_agg_write_addr_gen_0_strides_2,
  input logic [2:0] agg_only_agg_write_addr_gen_1_starting_addr,
  input logic [2:0] agg_only_agg_write_addr_gen_1_strides_0,
  input logic [2:0] agg_only_agg_write_addr_gen_1_strides_1,
  input logic [2:0] agg_only_agg_write_addr_gen_1_strides_2,
  input logic agg_only_agg_write_sched_gen_0_enable,
  input logic [15:0] agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [15:0] agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0,
  input logic [15:0] agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1,
  input logic [15:0] agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2,
  input logic agg_only_agg_write_sched_gen_1_enable,
  input logic [15:0] agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [15:0] agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0,
  input logic [15:0] agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1,
  input logic [15:0] agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2,
  input logic [2:0] agg_only_loops_in2buf_0_dimensionality,
  input logic [10:0] agg_only_loops_in2buf_0_ranges_0,
  input logic [10:0] agg_only_loops_in2buf_0_ranges_1,
  input logic [10:0] agg_only_loops_in2buf_0_ranges_2,
  input logic [2:0] agg_only_loops_in2buf_1_dimensionality,
  input logic [10:0] agg_only_loops_in2buf_1_ranges_0,
  input logic [10:0] agg_only_loops_in2buf_1_ranges_1,
  input logic [10:0] agg_only_loops_in2buf_1_ranges_2,
  input logic [7:0] agg_sram_shared_agg_read_sched_gen_0_agg_read_padding,
  input logic [7:0] agg_sram_shared_agg_read_sched_gen_1_agg_read_padding,
  input logic [8:0] agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr,
  input logic [8:0] agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr,
  input logic [1:0] agg_sram_shared_mode_0,
  input logic [1:0] agg_sram_shared_mode_1,
  input logic chain_chain_en,
  input logic [1:0] [16:0] chain_data_in,
  input logic clk,
  input logic clk_en,
  input logic [3:0] [15:0] data_from_strg,
  input logic [1:0] [16:0] data_in,
  input logic flush,
  input logic rst_n,
  input logic [8:0] sram_only_output_addr_gen_0_starting_addr,
  input logic [8:0] sram_only_output_addr_gen_0_strides_0,
  input logic [8:0] sram_only_output_addr_gen_0_strides_1,
  input logic [8:0] sram_only_output_addr_gen_0_strides_2,
  input logic [8:0] sram_only_output_addr_gen_0_strides_3,
  input logic [8:0] sram_only_output_addr_gen_0_strides_4,
  input logic [8:0] sram_only_output_addr_gen_0_strides_5,
  input logic [8:0] sram_only_output_addr_gen_1_starting_addr,
  input logic [8:0] sram_only_output_addr_gen_1_strides_0,
  input logic [8:0] sram_only_output_addr_gen_1_strides_1,
  input logic [8:0] sram_only_output_addr_gen_1_strides_2,
  input logic [8:0] sram_only_output_addr_gen_1_strides_3,
  input logic [8:0] sram_only_output_addr_gen_1_strides_4,
  input logic [8:0] sram_only_output_addr_gen_1_strides_5,
  input logic [3:0] sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality,
  input logic [10:0] sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0,
  input logic [10:0] sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1,
  input logic [10:0] sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2,
  input logic [10:0] sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3,
  input logic [10:0] sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4,
  input logic [10:0] sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5,
  input logic [3:0] sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality,
  input logic [10:0] sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0,
  input logic [10:0] sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1,
  input logic [10:0] sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2,
  input logic [10:0] sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3,
  input logic [10:0] sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4,
  input logic [10:0] sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5,
  input logic sram_tb_shared_output_sched_gen_0_enable,
  input logic [9:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay,
  input logic [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0,
  input logic [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1,
  input logic [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2,
  input logic [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3,
  input logic [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4,
  input logic [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5,
  input logic sram_tb_shared_output_sched_gen_1_enable,
  input logic [9:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay,
  input logic [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0,
  input logic [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1,
  input logic [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2,
  input logic [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3,
  input logic [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4,
  input logic [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5,
  input logic [3:0] tb_only_loops_buf2out_read_0_dimensionality,
  input logic [10:0] tb_only_loops_buf2out_read_0_ranges_0,
  input logic [10:0] tb_only_loops_buf2out_read_0_ranges_1,
  input logic [10:0] tb_only_loops_buf2out_read_0_ranges_2,
  input logic [10:0] tb_only_loops_buf2out_read_0_ranges_3,
  input logic [10:0] tb_only_loops_buf2out_read_0_ranges_4,
  input logic [10:0] tb_only_loops_buf2out_read_0_ranges_5,
  input logic [3:0] tb_only_loops_buf2out_read_1_dimensionality,
  input logic [10:0] tb_only_loops_buf2out_read_1_ranges_0,
  input logic [10:0] tb_only_loops_buf2out_read_1_ranges_1,
  input logic [10:0] tb_only_loops_buf2out_read_1_ranges_2,
  input logic [10:0] tb_only_loops_buf2out_read_1_ranges_3,
  input logic [10:0] tb_only_loops_buf2out_read_1_ranges_4,
  input logic [10:0] tb_only_loops_buf2out_read_1_ranges_5,
  input logic tb_only_shared_tb_0,
  input logic [3:0] tb_only_tb_read_addr_gen_0_starting_addr,
  input logic [3:0] tb_only_tb_read_addr_gen_0_strides_0,
  input logic [3:0] tb_only_tb_read_addr_gen_0_strides_1,
  input logic [3:0] tb_only_tb_read_addr_gen_0_strides_2,
  input logic [3:0] tb_only_tb_read_addr_gen_0_strides_3,
  input logic [3:0] tb_only_tb_read_addr_gen_0_strides_4,
  input logic [3:0] tb_only_tb_read_addr_gen_0_strides_5,
  input logic [3:0] tb_only_tb_read_addr_gen_1_starting_addr,
  input logic [3:0] tb_only_tb_read_addr_gen_1_strides_0,
  input logic [3:0] tb_only_tb_read_addr_gen_1_strides_1,
  input logic [3:0] tb_only_tb_read_addr_gen_1_strides_2,
  input logic [3:0] tb_only_tb_read_addr_gen_1_strides_3,
  input logic [3:0] tb_only_tb_read_addr_gen_1_strides_4,
  input logic [3:0] tb_only_tb_read_addr_gen_1_strides_5,
  input logic tb_only_tb_read_sched_gen_0_enable,
  input logic [9:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_delay,
  input logic [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0,
  input logic [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1,
  input logic [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2,
  input logic [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3,
  input logic [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4,
  input logic [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5,
  input logic tb_only_tb_read_sched_gen_1_enable,
  input logic [9:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_delay,
  input logic [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0,
  input logic [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1,
  input logic [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2,
  input logic [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3,
  input logic [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4,
  input logic [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5,
  input logic [3:0] tb_only_tb_write_addr_gen_0_starting_addr,
  input logic [3:0] tb_only_tb_write_addr_gen_0_strides_0,
  input logic [3:0] tb_only_tb_write_addr_gen_0_strides_1,
  input logic [3:0] tb_only_tb_write_addr_gen_0_strides_2,
  input logic [3:0] tb_only_tb_write_addr_gen_0_strides_3,
  input logic [3:0] tb_only_tb_write_addr_gen_0_strides_4,
  input logic [3:0] tb_only_tb_write_addr_gen_0_strides_5,
  input logic [3:0] tb_only_tb_write_addr_gen_1_starting_addr,
  input logic [3:0] tb_only_tb_write_addr_gen_1_strides_0,
  input logic [3:0] tb_only_tb_write_addr_gen_1_strides_1,
  input logic [3:0] tb_only_tb_write_addr_gen_1_strides_2,
  input logic [3:0] tb_only_tb_write_addr_gen_1_strides_3,
  input logic [3:0] tb_only_tb_write_addr_gen_1_strides_4,
  input logic [3:0] tb_only_tb_write_addr_gen_1_strides_5,
  output logic [1:0] accessor_output,
  output logic [8:0] addr_out,
  output logic [1:0] [16:0] data_out,
  output logic [3:0] [15:0] data_to_strg,
  output logic ren_to_strg,
  output logic wen_to_strg
);

logic [1:0] accessor_output_int;
logic [1:0][3:0][15:0] agg_only_agg_data_out;
logic [1:0] agg_only_agg_read;
logic [1:0][1:0] agg_only_agg_write_addr_l2b_out;
logic [1:0][2:0] agg_only_agg_write_mux_sel_out;
logic [1:0] agg_only_agg_write_out;
logic [1:0] agg_only_agg_write_restart_out;
logic [1:0][8:0] agg_only_sram_read_addr_in;
logic [1:0][2:0] agg_only_tb_read_addr_d_in;
logic [1:0] agg_only_tb_read_d_in;
logic [1:0][1:0] agg_only_update_mode_in;
logic [1:0] agg_sram_shared_agg_read_out;
logic [1:0][8:0] agg_sram_shared_agg_sram_shared_addr_out;
logic [1:0][8:0] agg_sram_shared_sram_read_addr_in;
logic [1:0] agg_sram_shared_sram_read_d_in;
logic [1:0] agg_sram_shared_sram_read_in;
logic [1:0][15:0] chain_data_in_thin;
logic [15:0] cycle_count;
logic [1:0][15:0] data_in_thin;
logic [1:0][15:0] data_out_int;
logic [1:0][15:0] data_out_int_thin;
logic [1:0][2:0] sram_only_loops_sram2tb_mux_sel;
logic [1:0] sram_only_loops_sram2tb_restart;
logic [1:0] sram_only_t_read;
logic [1:0][2:0] sram_tb_shared_loops_sram2tb_mux_sel;
logic [1:0] sram_tb_shared_loops_sram2tb_restart;
logic [1:0] sram_tb_shared_t_read_out;
assign data_in_thin[0] = data_in[0][15:0];
assign data_in_thin[1] = data_in[1][15:0];
assign data_out[0][15:0] = data_out_int_thin[0];
assign data_out[0][16] = 1'h0;
assign data_out[1][15:0] = data_out_int_thin[1];
assign data_out[1][16] = 1'h0;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    cycle_count <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      cycle_count <= 16'h0;
    end
    else if (1'h1) begin
      cycle_count <= cycle_count + 16'h1;
    end
  end
end
assign agg_only_sram_read_addr_in = agg_sram_shared_agg_sram_shared_addr_out;
assign agg_sram_shared_sram_read_in = sram_tb_shared_t_read_out;
assign agg_only_agg_read = agg_sram_shared_agg_read_out;
assign sram_only_loops_sram2tb_mux_sel = sram_tb_shared_loops_sram2tb_mux_sel;
assign sram_only_loops_sram2tb_restart = sram_tb_shared_loops_sram2tb_restart;
assign sram_only_t_read = sram_tb_shared_t_read_out;
assign ren_to_strg = |sram_tb_shared_t_read_out;
assign chain_data_in_thin[0] = chain_data_in[0][15:0];
assign chain_data_in_thin[1] = chain_data_in[1][15:0];
assign accessor_output = accessor_output_int;
strg_ub_agg_only agg_only (
  .agg_read(agg_only_agg_read),
  .agg_write_addr_gen_0_starting_addr(agg_only_agg_write_addr_gen_0_starting_addr),
  .agg_write_addr_gen_0_strides_0(agg_only_agg_write_addr_gen_0_strides_0),
  .agg_write_addr_gen_0_strides_1(agg_only_agg_write_addr_gen_0_strides_1),
  .agg_write_addr_gen_0_strides_2(agg_only_agg_write_addr_gen_0_strides_2),
  .agg_write_addr_gen_1_starting_addr(agg_only_agg_write_addr_gen_1_starting_addr),
  .agg_write_addr_gen_1_strides_0(agg_only_agg_write_addr_gen_1_strides_0),
  .agg_write_addr_gen_1_strides_1(agg_only_agg_write_addr_gen_1_strides_1),
  .agg_write_addr_gen_1_strides_2(agg_only_agg_write_addr_gen_1_strides_2),
  .agg_write_sched_gen_0_enable(agg_only_agg_write_sched_gen_0_enable),
  .agg_write_sched_gen_0_sched_addr_gen_starting_addr(agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr),
  .agg_write_sched_gen_0_sched_addr_gen_strides_0(agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0),
  .agg_write_sched_gen_0_sched_addr_gen_strides_1(agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1),
  .agg_write_sched_gen_0_sched_addr_gen_strides_2(agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2),
  .agg_write_sched_gen_1_enable(agg_only_agg_write_sched_gen_1_enable),
  .agg_write_sched_gen_1_sched_addr_gen_starting_addr(agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr),
  .agg_write_sched_gen_1_sched_addr_gen_strides_0(agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0),
  .agg_write_sched_gen_1_sched_addr_gen_strides_1(agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1),
  .agg_write_sched_gen_1_sched_addr_gen_strides_2(agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2),
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .data_in(data_in_thin),
  .flush(flush),
  .loops_in2buf_0_dimensionality(agg_only_loops_in2buf_0_dimensionality),
  .loops_in2buf_0_ranges_0(agg_only_loops_in2buf_0_ranges_0),
  .loops_in2buf_0_ranges_1(agg_only_loops_in2buf_0_ranges_1),
  .loops_in2buf_0_ranges_2(agg_only_loops_in2buf_0_ranges_2),
  .loops_in2buf_1_dimensionality(agg_only_loops_in2buf_1_dimensionality),
  .loops_in2buf_1_ranges_0(agg_only_loops_in2buf_1_ranges_0),
  .loops_in2buf_1_ranges_1(agg_only_loops_in2buf_1_ranges_1),
  .loops_in2buf_1_ranges_2(agg_only_loops_in2buf_1_ranges_2),
  .rst_n(rst_n),
  .sram_read_addr_in(agg_only_sram_read_addr_in),
  .tb_read_addr_d_in(agg_only_tb_read_addr_d_in),
  .tb_read_d_in(agg_only_tb_read_d_in),
  .update_mode_in(agg_only_update_mode_in),
  .agg_data_out(agg_only_agg_data_out),
  .agg_write_addr_l2b_out(agg_only_agg_write_addr_l2b_out),
  .agg_write_mux_sel_out(agg_only_agg_write_mux_sel_out),
  .agg_write_out(agg_only_agg_write_out),
  .agg_write_restart_out(agg_only_agg_write_restart_out)
);

strg_ub_agg_sram_shared agg_sram_shared (
  .agg_read_sched_gen_0_agg_read_padding(agg_sram_shared_agg_read_sched_gen_0_agg_read_padding),
  .agg_read_sched_gen_1_agg_read_padding(agg_sram_shared_agg_read_sched_gen_1_agg_read_padding),
  .agg_sram_shared_addr_gen_0_starting_addr(agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr),
  .agg_sram_shared_addr_gen_1_starting_addr(agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr),
  .agg_write_addr_l2b_in(agg_only_agg_write_addr_l2b_out),
  .agg_write_in(agg_only_agg_write_out),
  .agg_write_mux_sel_in(agg_only_agg_write_mux_sel_out),
  .agg_write_restart_in(agg_only_agg_write_restart_out),
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mode_0(agg_sram_shared_mode_0),
  .mode_1(agg_sram_shared_mode_1),
  .rst_n(rst_n),
  .sram_read_addr_in(agg_sram_shared_sram_read_addr_in),
  .sram_read_d_in(agg_sram_shared_sram_read_d_in),
  .sram_read_in(agg_sram_shared_sram_read_in),
  .agg_read_out(agg_sram_shared_agg_read_out),
  .agg_sram_shared_addr_out(agg_sram_shared_agg_sram_shared_addr_out),
  .update_mode_out(agg_only_update_mode_in)
);

strg_ub_sram_only sram_only (
  .agg_data_out(agg_only_agg_data_out),
  .agg_read(agg_sram_shared_agg_read_out),
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .flush(flush),
  .loops_sram2tb_mux_sel(sram_only_loops_sram2tb_mux_sel),
  .loops_sram2tb_restart(sram_only_loops_sram2tb_restart),
  .output_addr_gen_0_starting_addr(sram_only_output_addr_gen_0_starting_addr),
  .output_addr_gen_0_strides_0(sram_only_output_addr_gen_0_strides_0),
  .output_addr_gen_0_strides_1(sram_only_output_addr_gen_0_strides_1),
  .output_addr_gen_0_strides_2(sram_only_output_addr_gen_0_strides_2),
  .output_addr_gen_0_strides_3(sram_only_output_addr_gen_0_strides_3),
  .output_addr_gen_0_strides_4(sram_only_output_addr_gen_0_strides_4),
  .output_addr_gen_0_strides_5(sram_only_output_addr_gen_0_strides_5),
  .output_addr_gen_1_starting_addr(sram_only_output_addr_gen_1_starting_addr),
  .output_addr_gen_1_strides_0(sram_only_output_addr_gen_1_strides_0),
  .output_addr_gen_1_strides_1(sram_only_output_addr_gen_1_strides_1),
  .output_addr_gen_1_strides_2(sram_only_output_addr_gen_1_strides_2),
  .output_addr_gen_1_strides_3(sram_only_output_addr_gen_1_strides_3),
  .output_addr_gen_1_strides_4(sram_only_output_addr_gen_1_strides_4),
  .output_addr_gen_1_strides_5(sram_only_output_addr_gen_1_strides_5),
  .rst_n(rst_n),
  .sram_read_addr_in(agg_sram_shared_agg_sram_shared_addr_out),
  .t_read(sram_only_t_read),
  .addr_to_sram(addr_out),
  .data_to_sram(data_to_strg),
  .sram_read_addr_out(agg_sram_shared_sram_read_addr_in),
  .wen_to_sram(wen_to_strg)
);

strg_ub_sram_tb_shared sram_tb_shared (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .flush(flush),
  .loops_buf2out_autovec_read_0_dimensionality(sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality),
  .loops_buf2out_autovec_read_0_ranges_0(sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0),
  .loops_buf2out_autovec_read_0_ranges_1(sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1),
  .loops_buf2out_autovec_read_0_ranges_2(sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2),
  .loops_buf2out_autovec_read_0_ranges_3(sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3),
  .loops_buf2out_autovec_read_0_ranges_4(sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4),
  .loops_buf2out_autovec_read_0_ranges_5(sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5),
  .loops_buf2out_autovec_read_1_dimensionality(sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality),
  .loops_buf2out_autovec_read_1_ranges_0(sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0),
  .loops_buf2out_autovec_read_1_ranges_1(sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1),
  .loops_buf2out_autovec_read_1_ranges_2(sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2),
  .loops_buf2out_autovec_read_1_ranges_3(sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3),
  .loops_buf2out_autovec_read_1_ranges_4(sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4),
  .loops_buf2out_autovec_read_1_ranges_5(sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5),
  .output_sched_gen_0_enable(sram_tb_shared_output_sched_gen_0_enable),
  .output_sched_gen_0_sched_addr_gen_delay(sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay),
  .output_sched_gen_0_sched_addr_gen_starting_addr(sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr),
  .output_sched_gen_0_sched_addr_gen_strides_0(sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0),
  .output_sched_gen_0_sched_addr_gen_strides_1(sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1),
  .output_sched_gen_0_sched_addr_gen_strides_2(sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2),
  .output_sched_gen_0_sched_addr_gen_strides_3(sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3),
  .output_sched_gen_0_sched_addr_gen_strides_4(sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4),
  .output_sched_gen_0_sched_addr_gen_strides_5(sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5),
  .output_sched_gen_1_enable(sram_tb_shared_output_sched_gen_1_enable),
  .output_sched_gen_1_sched_addr_gen_delay(sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay),
  .output_sched_gen_1_sched_addr_gen_starting_addr(sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr),
  .output_sched_gen_1_sched_addr_gen_strides_0(sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0),
  .output_sched_gen_1_sched_addr_gen_strides_1(sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1),
  .output_sched_gen_1_sched_addr_gen_strides_2(sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2),
  .output_sched_gen_1_sched_addr_gen_strides_3(sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3),
  .output_sched_gen_1_sched_addr_gen_strides_4(sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4),
  .output_sched_gen_1_sched_addr_gen_strides_5(sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5),
  .rst_n(rst_n),
  .loops_sram2tb_mux_sel(sram_tb_shared_loops_sram2tb_mux_sel),
  .loops_sram2tb_restart(sram_tb_shared_loops_sram2tb_restart),
  .sram_read_d(agg_sram_shared_sram_read_d_in),
  .t_read_out(sram_tb_shared_t_read_out)
);

strg_ub_tb_only tb_only (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .flush(flush),
  .loops_buf2out_read_0_dimensionality(tb_only_loops_buf2out_read_0_dimensionality),
  .loops_buf2out_read_0_ranges_0(tb_only_loops_buf2out_read_0_ranges_0),
  .loops_buf2out_read_0_ranges_1(tb_only_loops_buf2out_read_0_ranges_1),
  .loops_buf2out_read_0_ranges_2(tb_only_loops_buf2out_read_0_ranges_2),
  .loops_buf2out_read_0_ranges_3(tb_only_loops_buf2out_read_0_ranges_3),
  .loops_buf2out_read_0_ranges_4(tb_only_loops_buf2out_read_0_ranges_4),
  .loops_buf2out_read_0_ranges_5(tb_only_loops_buf2out_read_0_ranges_5),
  .loops_buf2out_read_1_dimensionality(tb_only_loops_buf2out_read_1_dimensionality),
  .loops_buf2out_read_1_ranges_0(tb_only_loops_buf2out_read_1_ranges_0),
  .loops_buf2out_read_1_ranges_1(tb_only_loops_buf2out_read_1_ranges_1),
  .loops_buf2out_read_1_ranges_2(tb_only_loops_buf2out_read_1_ranges_2),
  .loops_buf2out_read_1_ranges_3(tb_only_loops_buf2out_read_1_ranges_3),
  .loops_buf2out_read_1_ranges_4(tb_only_loops_buf2out_read_1_ranges_4),
  .loops_buf2out_read_1_ranges_5(tb_only_loops_buf2out_read_1_ranges_5),
  .loops_sram2tb_mux_sel(sram_tb_shared_loops_sram2tb_mux_sel),
  .loops_sram2tb_restart(sram_tb_shared_loops_sram2tb_restart),
  .rst_n(rst_n),
  .shared_tb_0(tb_only_shared_tb_0),
  .sram_read_data(data_from_strg),
  .t_read(sram_tb_shared_t_read_out),
  .tb_read_addr_gen_0_starting_addr(tb_only_tb_read_addr_gen_0_starting_addr),
  .tb_read_addr_gen_0_strides_0(tb_only_tb_read_addr_gen_0_strides_0),
  .tb_read_addr_gen_0_strides_1(tb_only_tb_read_addr_gen_0_strides_1),
  .tb_read_addr_gen_0_strides_2(tb_only_tb_read_addr_gen_0_strides_2),
  .tb_read_addr_gen_0_strides_3(tb_only_tb_read_addr_gen_0_strides_3),
  .tb_read_addr_gen_0_strides_4(tb_only_tb_read_addr_gen_0_strides_4),
  .tb_read_addr_gen_0_strides_5(tb_only_tb_read_addr_gen_0_strides_5),
  .tb_read_addr_gen_1_starting_addr(tb_only_tb_read_addr_gen_1_starting_addr),
  .tb_read_addr_gen_1_strides_0(tb_only_tb_read_addr_gen_1_strides_0),
  .tb_read_addr_gen_1_strides_1(tb_only_tb_read_addr_gen_1_strides_1),
  .tb_read_addr_gen_1_strides_2(tb_only_tb_read_addr_gen_1_strides_2),
  .tb_read_addr_gen_1_strides_3(tb_only_tb_read_addr_gen_1_strides_3),
  .tb_read_addr_gen_1_strides_4(tb_only_tb_read_addr_gen_1_strides_4),
  .tb_read_addr_gen_1_strides_5(tb_only_tb_read_addr_gen_1_strides_5),
  .tb_read_sched_gen_0_enable(tb_only_tb_read_sched_gen_0_enable),
  .tb_read_sched_gen_0_sched_addr_gen_delay(tb_only_tb_read_sched_gen_0_sched_addr_gen_delay),
  .tb_read_sched_gen_0_sched_addr_gen_starting_addr(tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr),
  .tb_read_sched_gen_0_sched_addr_gen_strides_0(tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0),
  .tb_read_sched_gen_0_sched_addr_gen_strides_1(tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1),
  .tb_read_sched_gen_0_sched_addr_gen_strides_2(tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2),
  .tb_read_sched_gen_0_sched_addr_gen_strides_3(tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3),
  .tb_read_sched_gen_0_sched_addr_gen_strides_4(tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4),
  .tb_read_sched_gen_0_sched_addr_gen_strides_5(tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5),
  .tb_read_sched_gen_1_enable(tb_only_tb_read_sched_gen_1_enable),
  .tb_read_sched_gen_1_sched_addr_gen_delay(tb_only_tb_read_sched_gen_1_sched_addr_gen_delay),
  .tb_read_sched_gen_1_sched_addr_gen_starting_addr(tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr),
  .tb_read_sched_gen_1_sched_addr_gen_strides_0(tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0),
  .tb_read_sched_gen_1_sched_addr_gen_strides_1(tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1),
  .tb_read_sched_gen_1_sched_addr_gen_strides_2(tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2),
  .tb_read_sched_gen_1_sched_addr_gen_strides_3(tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3),
  .tb_read_sched_gen_1_sched_addr_gen_strides_4(tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4),
  .tb_read_sched_gen_1_sched_addr_gen_strides_5(tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5),
  .tb_write_addr_gen_0_starting_addr(tb_only_tb_write_addr_gen_0_starting_addr),
  .tb_write_addr_gen_0_strides_0(tb_only_tb_write_addr_gen_0_strides_0),
  .tb_write_addr_gen_0_strides_1(tb_only_tb_write_addr_gen_0_strides_1),
  .tb_write_addr_gen_0_strides_2(tb_only_tb_write_addr_gen_0_strides_2),
  .tb_write_addr_gen_0_strides_3(tb_only_tb_write_addr_gen_0_strides_3),
  .tb_write_addr_gen_0_strides_4(tb_only_tb_write_addr_gen_0_strides_4),
  .tb_write_addr_gen_0_strides_5(tb_only_tb_write_addr_gen_0_strides_5),
  .tb_write_addr_gen_1_starting_addr(tb_only_tb_write_addr_gen_1_starting_addr),
  .tb_write_addr_gen_1_strides_0(tb_only_tb_write_addr_gen_1_strides_0),
  .tb_write_addr_gen_1_strides_1(tb_only_tb_write_addr_gen_1_strides_1),
  .tb_write_addr_gen_1_strides_2(tb_only_tb_write_addr_gen_1_strides_2),
  .tb_write_addr_gen_1_strides_3(tb_only_tb_write_addr_gen_1_strides_3),
  .tb_write_addr_gen_1_strides_4(tb_only_tb_write_addr_gen_1_strides_4),
  .tb_write_addr_gen_1_strides_5(tb_only_tb_write_addr_gen_1_strides_5),
  .accessor_output(accessor_output_int),
  .data_out(data_out_int),
  .tb_read_addr_d_out(agg_only_tb_read_addr_d_in),
  .tb_read_d_out(agg_only_tb_read_d_in)
);

Chain_2_16 chain (
  .accessor_output(accessor_output_int),
  .chain_data_in(chain_data_in_thin),
  .chain_en(chain_chain_en),
  .clk_en(clk_en),
  .curr_tile_data_out(data_out_int),
  .flush(flush),
  .data_out_tile(data_out_int_thin)
);

endmodule   // strg_ub_vec

module strg_ub_vec_flat (
  input logic [0:0] [16:0] chain_data_in_f_0,
  input logic [0:0] [16:0] chain_data_in_f_1,
  input logic clk,
  input logic clk_en,
  input logic [0:0] [16:0] data_in_f_0,
  input logic [0:0] [16:0] data_in_f_1,
  input logic flush,
  input logic rst_n,
  input logic [2:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr,
  input logic [2:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0,
  input logic [2:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1,
  input logic [2:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2,
  input logic [2:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr,
  input logic [2:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0,
  input logic [2:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1,
  input logic [2:0] strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2,
  input logic strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable,
  input logic [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0,
  input logic [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1,
  input logic [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2,
  input logic strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable,
  input logic [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0,
  input logic [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1,
  input logic [15:0] strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2,
  input logic [2:0] strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality,
  input logic [10:0] strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0,
  input logic [10:0] strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1,
  input logic [10:0] strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2,
  input logic [2:0] strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality,
  input logic [10:0] strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0,
  input logic [10:0] strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1,
  input logic [10:0] strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2,
  input logic [7:0] strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_agg_read_padding,
  input logic [7:0] strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_agg_read_padding,
  input logic [8:0] strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr,
  input logic [8:0] strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr,
  input logic [1:0] strg_ub_vec_inst_agg_sram_shared_mode_0,
  input logic [1:0] strg_ub_vec_inst_agg_sram_shared_mode_1,
  input logic strg_ub_vec_inst_chain_chain_en,
  input logic [3:0] [15:0] strg_ub_vec_inst_data_from_strg_lifted,
  input logic [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr,
  input logic [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0,
  input logic [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1,
  input logic [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2,
  input logic [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3,
  input logic [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4,
  input logic [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5,
  input logic [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr,
  input logic [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0,
  input logic [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1,
  input logic [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2,
  input logic [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3,
  input logic [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4,
  input logic [8:0] strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5,
  input logic [3:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality,
  input logic [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0,
  input logic [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1,
  input logic [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2,
  input logic [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3,
  input logic [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4,
  input logic [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5,
  input logic [3:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality,
  input logic [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0,
  input logic [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1,
  input logic [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2,
  input logic [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3,
  input logic [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4,
  input logic [10:0] strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5,
  input logic strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable,
  input logic [9:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay,
  input logic [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0,
  input logic [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1,
  input logic [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2,
  input logic [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3,
  input logic [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4,
  input logic [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5,
  input logic strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable,
  input logic [9:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay,
  input logic [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0,
  input logic [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1,
  input logic [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2,
  input logic [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3,
  input logic [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4,
  input logic [15:0] strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5,
  input logic [3:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality,
  input logic [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0,
  input logic [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1,
  input logic [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2,
  input logic [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3,
  input logic [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4,
  input logic [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5,
  input logic [3:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality,
  input logic [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0,
  input logic [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1,
  input logic [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2,
  input logic [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3,
  input logic [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4,
  input logic [10:0] strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5,
  input logic strg_ub_vec_inst_tb_only_shared_tb_0,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5,
  input logic strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable,
  input logic [9:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_delay,
  input logic [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0,
  input logic [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1,
  input logic [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2,
  input logic [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3,
  input logic [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4,
  input logic [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5,
  input logic strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable,
  input logic [9:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_delay,
  input logic [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0,
  input logic [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1,
  input logic [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2,
  input logic [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3,
  input logic [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4,
  input logic [15:0] strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4,
  input logic [3:0] strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5,
  output logic accessor_output_f_b_0,
  output logic accessor_output_f_b_1,
  output logic [0:0] [16:0] data_out_f_0,
  output logic [0:0] [16:0] data_out_f_1,
  output logic [8:0] strg_ub_vec_inst_addr_out_lifted,
  output logic [3:0] [15:0] strg_ub_vec_inst_data_to_strg_lifted,
  output logic strg_ub_vec_inst_ren_to_strg_lifted,
  output logic strg_ub_vec_inst_wen_to_strg_lifted
);

logic [1:0] strg_ub_vec_inst_accessor_output;
logic [1:0][16:0] strg_ub_vec_inst_chain_data_in;
logic [1:0][16:0] strg_ub_vec_inst_data_in;
logic [1:0][16:0] strg_ub_vec_inst_data_out;
assign strg_ub_vec_inst_data_in[0] = data_in_f_0;
assign strg_ub_vec_inst_data_in[1] = data_in_f_1;
assign strg_ub_vec_inst_chain_data_in[0] = chain_data_in_f_0;
assign strg_ub_vec_inst_chain_data_in[1] = chain_data_in_f_1;
assign accessor_output_f_b_0 = strg_ub_vec_inst_accessor_output[0];
assign accessor_output_f_b_1 = strg_ub_vec_inst_accessor_output[1];
assign data_out_f_0 = strg_ub_vec_inst_data_out[0];
assign data_out_f_1 = strg_ub_vec_inst_data_out[1];
strg_ub_vec strg_ub_vec_inst (
  .agg_only_agg_write_addr_gen_0_starting_addr(strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_starting_addr),
  .agg_only_agg_write_addr_gen_0_strides_0(strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_0),
  .agg_only_agg_write_addr_gen_0_strides_1(strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_1),
  .agg_only_agg_write_addr_gen_0_strides_2(strg_ub_vec_inst_agg_only_agg_write_addr_gen_0_strides_2),
  .agg_only_agg_write_addr_gen_1_starting_addr(strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_starting_addr),
  .agg_only_agg_write_addr_gen_1_strides_0(strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_0),
  .agg_only_agg_write_addr_gen_1_strides_1(strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_1),
  .agg_only_agg_write_addr_gen_1_strides_2(strg_ub_vec_inst_agg_only_agg_write_addr_gen_1_strides_2),
  .agg_only_agg_write_sched_gen_0_enable(strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_enable),
  .agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr),
  .agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0(strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0),
  .agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1(strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1),
  .agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2(strg_ub_vec_inst_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2),
  .agg_only_agg_write_sched_gen_1_enable(strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_enable),
  .agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr),
  .agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0(strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0),
  .agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1(strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1),
  .agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2(strg_ub_vec_inst_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2),
  .agg_only_loops_in2buf_0_dimensionality(strg_ub_vec_inst_agg_only_loops_in2buf_0_dimensionality),
  .agg_only_loops_in2buf_0_ranges_0(strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_0),
  .agg_only_loops_in2buf_0_ranges_1(strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_1),
  .agg_only_loops_in2buf_0_ranges_2(strg_ub_vec_inst_agg_only_loops_in2buf_0_ranges_2),
  .agg_only_loops_in2buf_1_dimensionality(strg_ub_vec_inst_agg_only_loops_in2buf_1_dimensionality),
  .agg_only_loops_in2buf_1_ranges_0(strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_0),
  .agg_only_loops_in2buf_1_ranges_1(strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_1),
  .agg_only_loops_in2buf_1_ranges_2(strg_ub_vec_inst_agg_only_loops_in2buf_1_ranges_2),
  .agg_sram_shared_agg_read_sched_gen_0_agg_read_padding(strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_0_agg_read_padding),
  .agg_sram_shared_agg_read_sched_gen_1_agg_read_padding(strg_ub_vec_inst_agg_sram_shared_agg_read_sched_gen_1_agg_read_padding),
  .agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr(strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_0_starting_addr),
  .agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr(strg_ub_vec_inst_agg_sram_shared_agg_sram_shared_addr_gen_1_starting_addr),
  .agg_sram_shared_mode_0(strg_ub_vec_inst_agg_sram_shared_mode_0),
  .agg_sram_shared_mode_1(strg_ub_vec_inst_agg_sram_shared_mode_1),
  .chain_chain_en(strg_ub_vec_inst_chain_chain_en),
  .chain_data_in(strg_ub_vec_inst_chain_data_in),
  .clk(clk),
  .clk_en(clk_en),
  .data_from_strg(strg_ub_vec_inst_data_from_strg_lifted),
  .data_in(strg_ub_vec_inst_data_in),
  .flush(flush),
  .rst_n(rst_n),
  .sram_only_output_addr_gen_0_starting_addr(strg_ub_vec_inst_sram_only_output_addr_gen_0_starting_addr),
  .sram_only_output_addr_gen_0_strides_0(strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_0),
  .sram_only_output_addr_gen_0_strides_1(strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_1),
  .sram_only_output_addr_gen_0_strides_2(strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_2),
  .sram_only_output_addr_gen_0_strides_3(strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_3),
  .sram_only_output_addr_gen_0_strides_4(strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_4),
  .sram_only_output_addr_gen_0_strides_5(strg_ub_vec_inst_sram_only_output_addr_gen_0_strides_5),
  .sram_only_output_addr_gen_1_starting_addr(strg_ub_vec_inst_sram_only_output_addr_gen_1_starting_addr),
  .sram_only_output_addr_gen_1_strides_0(strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_0),
  .sram_only_output_addr_gen_1_strides_1(strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_1),
  .sram_only_output_addr_gen_1_strides_2(strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_2),
  .sram_only_output_addr_gen_1_strides_3(strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_3),
  .sram_only_output_addr_gen_1_strides_4(strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_4),
  .sram_only_output_addr_gen_1_strides_5(strg_ub_vec_inst_sram_only_output_addr_gen_1_strides_5),
  .sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality),
  .sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0),
  .sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1),
  .sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2),
  .sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3),
  .sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4),
  .sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5),
  .sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality),
  .sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0),
  .sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1),
  .sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2),
  .sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3),
  .sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4),
  .sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5(strg_ub_vec_inst_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5),
  .sram_tb_shared_output_sched_gen_0_enable(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_enable),
  .sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_delay),
  .sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr),
  .sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0),
  .sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1),
  .sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2),
  .sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3),
  .sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4),
  .sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5),
  .sram_tb_shared_output_sched_gen_1_enable(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_enable),
  .sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_delay),
  .sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr),
  .sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0),
  .sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1),
  .sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2),
  .sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3),
  .sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4),
  .sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5(strg_ub_vec_inst_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5),
  .tb_only_loops_buf2out_read_0_dimensionality(strg_ub_vec_inst_tb_only_loops_buf2out_read_0_dimensionality),
  .tb_only_loops_buf2out_read_0_ranges_0(strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_0),
  .tb_only_loops_buf2out_read_0_ranges_1(strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_1),
  .tb_only_loops_buf2out_read_0_ranges_2(strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_2),
  .tb_only_loops_buf2out_read_0_ranges_3(strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_3),
  .tb_only_loops_buf2out_read_0_ranges_4(strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_4),
  .tb_only_loops_buf2out_read_0_ranges_5(strg_ub_vec_inst_tb_only_loops_buf2out_read_0_ranges_5),
  .tb_only_loops_buf2out_read_1_dimensionality(strg_ub_vec_inst_tb_only_loops_buf2out_read_1_dimensionality),
  .tb_only_loops_buf2out_read_1_ranges_0(strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_0),
  .tb_only_loops_buf2out_read_1_ranges_1(strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_1),
  .tb_only_loops_buf2out_read_1_ranges_2(strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_2),
  .tb_only_loops_buf2out_read_1_ranges_3(strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_3),
  .tb_only_loops_buf2out_read_1_ranges_4(strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_4),
  .tb_only_loops_buf2out_read_1_ranges_5(strg_ub_vec_inst_tb_only_loops_buf2out_read_1_ranges_5),
  .tb_only_shared_tb_0(strg_ub_vec_inst_tb_only_shared_tb_0),
  .tb_only_tb_read_addr_gen_0_starting_addr(strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_starting_addr),
  .tb_only_tb_read_addr_gen_0_strides_0(strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_0),
  .tb_only_tb_read_addr_gen_0_strides_1(strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_1),
  .tb_only_tb_read_addr_gen_0_strides_2(strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_2),
  .tb_only_tb_read_addr_gen_0_strides_3(strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_3),
  .tb_only_tb_read_addr_gen_0_strides_4(strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_4),
  .tb_only_tb_read_addr_gen_0_strides_5(strg_ub_vec_inst_tb_only_tb_read_addr_gen_0_strides_5),
  .tb_only_tb_read_addr_gen_1_starting_addr(strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_starting_addr),
  .tb_only_tb_read_addr_gen_1_strides_0(strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_0),
  .tb_only_tb_read_addr_gen_1_strides_1(strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_1),
  .tb_only_tb_read_addr_gen_1_strides_2(strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_2),
  .tb_only_tb_read_addr_gen_1_strides_3(strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_3),
  .tb_only_tb_read_addr_gen_1_strides_4(strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_4),
  .tb_only_tb_read_addr_gen_1_strides_5(strg_ub_vec_inst_tb_only_tb_read_addr_gen_1_strides_5),
  .tb_only_tb_read_sched_gen_0_enable(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_enable),
  .tb_only_tb_read_sched_gen_0_sched_addr_gen_delay(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_delay),
  .tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr),
  .tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0),
  .tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1),
  .tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2),
  .tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3),
  .tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4),
  .tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5(strg_ub_vec_inst_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5),
  .tb_only_tb_read_sched_gen_1_enable(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_enable),
  .tb_only_tb_read_sched_gen_1_sched_addr_gen_delay(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_delay),
  .tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr),
  .tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0),
  .tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1),
  .tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2),
  .tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3),
  .tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4),
  .tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5(strg_ub_vec_inst_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5),
  .tb_only_tb_write_addr_gen_0_starting_addr(strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_starting_addr),
  .tb_only_tb_write_addr_gen_0_strides_0(strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_0),
  .tb_only_tb_write_addr_gen_0_strides_1(strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_1),
  .tb_only_tb_write_addr_gen_0_strides_2(strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_2),
  .tb_only_tb_write_addr_gen_0_strides_3(strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_3),
  .tb_only_tb_write_addr_gen_0_strides_4(strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_4),
  .tb_only_tb_write_addr_gen_0_strides_5(strg_ub_vec_inst_tb_only_tb_write_addr_gen_0_strides_5),
  .tb_only_tb_write_addr_gen_1_starting_addr(strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_starting_addr),
  .tb_only_tb_write_addr_gen_1_strides_0(strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_0),
  .tb_only_tb_write_addr_gen_1_strides_1(strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_1),
  .tb_only_tb_write_addr_gen_1_strides_2(strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_2),
  .tb_only_tb_write_addr_gen_1_strides_3(strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_3),
  .tb_only_tb_write_addr_gen_1_strides_4(strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_4),
  .tb_only_tb_write_addr_gen_1_strides_5(strg_ub_vec_inst_tb_only_tb_write_addr_gen_1_strides_5),
  .accessor_output(strg_ub_vec_inst_accessor_output),
  .addr_out(strg_ub_vec_inst_addr_out_lifted),
  .data_out(strg_ub_vec_inst_data_out),
  .data_to_strg(strg_ub_vec_inst_data_to_strg_lifted),
  .ren_to_strg(strg_ub_vec_inst_ren_to_strg_lifted),
  .wen_to_strg(strg_ub_vec_inst_wen_to_strg_lifted)
);

endmodule   // strg_ub_vec_flat

module write_scanner (
  input logic ID_out_ready,
  input logic [16:0] addr_in,
  input logic addr_in_valid,
  input logic addr_out_ready,
  input logic block_mode,
  input logic [16:0] block_wr_in,
  input logic block_wr_in_valid,
  input logic clk,
  input logic clk_en,
  input logic compressed,
  input logic [16:0] data_in,
  input logic data_in_valid,
  input logic data_out_ready,
  input logic flush,
  input logic init_blank,
  input logic lowest_level,
  input logic rst_n,
  input logic spacc_mode,
  input logic [15:0] stop_lvl,
  input logic tile_en,
  output logic [16:0] ID_out,
  output logic ID_out_valid,
  output logic addr_in_ready,
  output logic [16:0] addr_out,
  output logic addr_out_valid,
  output logic block_wr_in_ready,
  output logic data_in_ready,
  output logic [16:0] data_out,
  output logic data_out_valid
);

typedef enum logic[4:0] {
  ALLOCATE1 = 5'h0,
  ALLOCATE2 = 5'h1,
  BLOCK_1_SZ = 5'h2,
  BLOCK_1_WR = 5'h3,
  BLOCK_2_SZ = 5'h4,
  BLOCK_2_WR = 5'h5,
  ComLL = 5'h6,
  DONE = 5'h7,
  FINALIZE1 = 5'h8,
  FINALIZE2 = 5'h9,
  LL = 5'hA,
  START = 5'hB,
  UL = 5'hC,
  UL_EMIT_COORD = 5'hD,
  UL_EMIT_SEG = 5'hE,
  UL_WZ = 5'hF,
  UnLL = 5'h10
} scan_seq_state;
logic [0:0][16:0] ID_out_fifo_data_in;
logic ID_out_fifo_empty;
logic ID_out_fifo_full;
logic ID_out_fifo_push;
logic [15:0] ID_to_fifo;
logic addr_done_in;
logic [15:0] addr_infifo_data_in;
logic addr_infifo_eos_in;
logic [16:0] addr_infifo_in_packed;
logic [16:0] addr_infifo_out_packed;
logic addr_infifo_valid_in;
logic addr_input_fifo_empty;
logic addr_input_fifo_full;
logic [0:0][16:0] addr_out_fifo_data_in;
logic addr_out_fifo_empty;
logic addr_out_fifo_full;
logic addr_out_fifo_push;
logic [15:0] addr_to_fifo;
logic blank_done_stick_sticky;
logic blank_done_stick_was_high;
logic [15:0] block_size;
logic block_wr_fifo_valid;
logic [0:0][15:0] block_wr_input_fifo_data_out;
logic block_wr_input_fifo_empty;
logic block_wr_input_fifo_full;
logic [15:0] block_write_count;
logic clr_blank_done;
logic clr_block_write;
logic clr_coord_addr;
logic clr_curr_coord;
logic clr_seg_addr;
logic clr_seg_ctr;
logic clr_wen_made;
logic [15:0] coord_addr;
logic data_done_in;
logic [15:0] data_infifo_data_in;
logic [15:0] data_infifo_data_in_d1;
logic data_infifo_eos_in;
logic [16:0] data_infifo_in_packed;
logic [16:0] data_infifo_out_packed;
logic data_infifo_valid_in;
logic data_input_fifo_empty;
logic data_input_fifo_full;
logic [0:0][16:0] data_out_fifo_data_in;
logic data_out_fifo_empty;
logic data_out_fifo_full;
logic data_out_fifo_push;
logic [15:0] data_to_fifo;
logic gclk;
logic inc_block_write;
logic inc_coord_addr;
logic inc_seg_addr;
logic inc_seg_ctr;
logic [1:0] infifo_pop;
logic matching_stop;
logic new_coord;
logic op_to_fifo;
logic pop_block_wr;
logic push_to_outs;
scan_seq_state scan_seq_current_state;
scan_seq_state scan_seq_next_state;
logic [15:0] segment_addr;
logic [15:0] segment_counter;
logic set_blank_done;
logic set_block_size;
logic set_curr_coord;
logic stop_in;
logic stop_lvl_geq;
logic stop_lvl_geq_p1;
logic stop_lvl_new_blank_sticky_sticky;
logic stop_lvl_new_blank_sticky_was_high;
logic valid_coord_sticky_sticky;
logic valid_coord_sticky_was_high;
logic wen_made_sticky;
logic wen_made_was_high;
assign gclk = clk & tile_en;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    blank_done_stick_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      blank_done_stick_was_high <= 1'h0;
    end
    else if (clr_blank_done) begin
      blank_done_stick_was_high <= 1'h0;
    end
    else if (set_blank_done) begin
      blank_done_stick_was_high <= 1'h1;
    end
  end
end
assign blank_done_stick_sticky = blank_done_stick_was_high;
assign data_infifo_in_packed[16] = data_in[16];
assign data_infifo_in_packed[15:0] = data_in[15:0];
assign data_infifo_eos_in = data_infifo_out_packed[16];
assign data_infifo_data_in = data_infifo_out_packed[15:0];
assign data_in_ready = ~data_input_fifo_full;
assign data_infifo_valid_in = ~data_input_fifo_empty;
assign addr_infifo_in_packed[16] = addr_in[16];
assign addr_infifo_in_packed[15:0] = addr_in[15:0];
assign addr_infifo_eos_in = addr_infifo_out_packed[16];
assign addr_infifo_data_in = addr_infifo_out_packed[15:0];
assign addr_in_ready = ~addr_input_fifo_full;
assign addr_infifo_valid_in = ~addr_input_fifo_empty;
assign block_wr_in_ready = ~block_wr_input_fifo_full;
assign block_wr_fifo_valid = ~block_wr_input_fifo_empty;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    block_size <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      block_size <= 16'h0;
    end
    else if (1'h0) begin
      block_size <= 16'h0;
    end
    else if (set_block_size) begin
      block_size <= block_wr_input_fifo_data_out;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    block_write_count <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      block_write_count <= 16'h0;
    end
    else if (clr_block_write) begin
      block_write_count <= 16'h0;
    end
    else if (inc_block_write) begin
      block_write_count <= block_write_count + 16'h1;
    end
  end
end
assign data_out_fifo_data_in = {op_to_fifo, data_to_fifo};
assign data_out_valid = ~data_out_fifo_empty;
assign addr_out_fifo_data_in = {1'h0, addr_to_fifo};
assign addr_out_valid = ~addr_out_fifo_empty;
assign ID_out_fifo_data_in = {1'h0, ID_to_fifo};
assign ID_out_valid = ~ID_out_fifo_empty;
assign {data_out_fifo_push, addr_out_fifo_push, ID_out_fifo_push} = {push_to_outs, push_to_outs, push_to_outs};
assign stop_lvl_geq = data_infifo_eos_in & data_infifo_valid_in & (data_infifo_data_in[9:8] == 2'h0) &
    (data_infifo_data_in[7:0] >= stop_lvl[7:0]);
assign stop_lvl_geq_p1 = data_infifo_eos_in & data_infifo_valid_in & (data_infifo_data_in[9:8] == 2'h0) &
    (data_infifo_data_in[7:0] >= (stop_lvl[7:0] + 8'h1));

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    stop_lvl_new_blank_sticky_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      stop_lvl_new_blank_sticky_was_high <= 1'h0;
    end
    else if (clr_blank_done) begin
      stop_lvl_new_blank_sticky_was_high <= 1'h0;
    end
    else if (stop_lvl_geq_p1) begin
      stop_lvl_new_blank_sticky_was_high <= 1'h1;
    end
  end
end
assign stop_lvl_new_blank_sticky_sticky = stop_lvl_new_blank_sticky_was_high;
assign data_done_in = data_infifo_valid_in & data_infifo_eos_in & (data_infifo_data_in[9:8] == 2'h1);
assign addr_done_in = addr_infifo_valid_in & addr_infifo_eos_in & (addr_infifo_data_in[9:8] == 2'h1);

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    segment_addr <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      segment_addr <= 16'h0;
    end
    else if (clr_seg_addr) begin
      segment_addr <= 16'h0;
    end
    else if (inc_seg_addr) begin
      segment_addr <= segment_addr + 16'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    coord_addr <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      coord_addr <= 16'h0;
    end
    else if (clr_coord_addr) begin
      coord_addr <= 16'h0;
    end
    else if (inc_coord_addr) begin
      coord_addr <= coord_addr + 16'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    segment_counter <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      segment_counter <= 16'h0;
    end
    else if (clr_seg_ctr) begin
      segment_counter <= 16'h0;
    end
    else if (inc_seg_ctr) begin
      segment_counter <= segment_counter + 16'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    data_infifo_data_in_d1 <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      data_infifo_data_in_d1 <= 16'h0;
    end
    else if (1'h0) begin
      data_infifo_data_in_d1 <= 16'h0;
    end
    else if (set_curr_coord) begin
      data_infifo_data_in_d1 <= data_infifo_data_in;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    valid_coord_sticky_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      valid_coord_sticky_was_high <= 1'h0;
    end
    else if (clr_curr_coord) begin
      valid_coord_sticky_was_high <= 1'h0;
    end
    else if (set_curr_coord) begin
      valid_coord_sticky_was_high <= 1'h1;
    end
  end
end
assign valid_coord_sticky_sticky = valid_coord_sticky_was_high;
assign new_coord = data_infifo_valid_in & (~data_infifo_eos_in) & ((~valid_coord_sticky_sticky) |
    (data_infifo_data_in != data_infifo_data_in_d1));
assign stop_in = data_infifo_valid_in & data_infifo_eos_in;
assign matching_stop = data_infifo_valid_in & data_infifo_eos_in;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    wen_made_was_high <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      wen_made_was_high <= 1'h0;
    end
    else if (clr_wen_made) begin
      wen_made_was_high <= 1'h0;
    end
    else if (push_to_outs) begin
      wen_made_was_high <= 1'h1;
    end
  end
end
assign wen_made_sticky = wen_made_was_high;

always_ff @(posedge clk, negedge rst_n) begin
  if (!rst_n) begin
    scan_seq_current_state <= START;
  end
  else if (clk_en) begin
    if (flush) begin
      scan_seq_current_state <= START;
    end
    else scan_seq_current_state <= scan_seq_next_state;
  end
end
always_comb begin
  scan_seq_next_state = scan_seq_current_state;
  unique case (scan_seq_current_state)
    ALLOCATE1: begin
        if (~(&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}))) begin
          scan_seq_next_state = ALLOCATE1;
        end
        else if ((~lowest_level) & (&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}))) begin
          scan_seq_next_state = ALLOCATE2;
        end
        else if (lowest_level & block_mode & (&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}))) begin
          scan_seq_next_state = BLOCK_1_SZ;
        end
        else if (lowest_level & (~block_mode) & (&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}))) begin
          scan_seq_next_state = LL;
        end
      end
    ALLOCATE2: begin
        if (~(&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}))) begin
          scan_seq_next_state = ALLOCATE2;
        end
        else if (block_mode & (&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}))) begin
          scan_seq_next_state = BLOCK_1_SZ;
        end
        else if ((~block_mode) & (&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}))) begin
          scan_seq_next_state = UL_WZ;
        end
      end
    BLOCK_1_SZ: begin
        if (block_wr_fifo_valid) begin
          scan_seq_next_state = BLOCK_1_WR;
        end
        else scan_seq_next_state = BLOCK_1_SZ;
      end
    BLOCK_1_WR: begin
        if ((block_write_count == block_size) & (~lowest_level)) begin
          scan_seq_next_state = BLOCK_2_SZ;
        end
        else if ((block_write_count == block_size) & lowest_level) begin
          scan_seq_next_state = FINALIZE2;
        end
        else scan_seq_next_state = BLOCK_1_WR;
      end
    BLOCK_2_SZ: begin
        if (block_wr_fifo_valid) begin
          scan_seq_next_state = BLOCK_2_WR;
        end
        else scan_seq_next_state = BLOCK_2_SZ;
      end
    BLOCK_2_WR: begin
        if (block_write_count == block_size) begin
          scan_seq_next_state = FINALIZE1;
        end
        else scan_seq_next_state = BLOCK_2_WR;
      end
    ComLL: begin
        if (data_done_in | (spacc_mode & stop_lvl_geq)) begin
          scan_seq_next_state = FINALIZE2;
        end
        else scan_seq_next_state = ComLL;
      end
    DONE: scan_seq_next_state = START;
    FINALIZE1: begin
        if (&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full})) begin
          scan_seq_next_state = FINALIZE2;
        end
        else scan_seq_next_state = FINALIZE1;
      end
    FINALIZE2: begin
        if (&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full})) begin
          scan_seq_next_state = DONE;
        end
        else scan_seq_next_state = FINALIZE2;
      end
    LL: begin
        if (init_blank & (~blank_done_stick_sticky)) begin
          scan_seq_next_state = FINALIZE2;
        end
        else if (compressed & ((~init_blank) | blank_done_stick_sticky)) begin
          scan_seq_next_state = ComLL;
        end
        else if ((~compressed) & ((~init_blank) | blank_done_stick_sticky)) begin
          scan_seq_next_state = UnLL;
        end
      end
    START: begin
        if (tile_en) begin
          scan_seq_next_state = ALLOCATE1;
        end
        else scan_seq_next_state = START;
      end
    UL: begin
        if (new_coord) begin
          scan_seq_next_state = UL_EMIT_COORD;
        end
        else if (matching_stop | (init_blank & (~blank_done_stick_sticky))) begin
          scan_seq_next_state = UL_EMIT_SEG;
        end
        else scan_seq_next_state = UL;
      end
    UL_EMIT_COORD: begin
        if (new_coord | stop_in) begin
          scan_seq_next_state = UL;
        end
        else scan_seq_next_state = UL_EMIT_COORD;
      end
    UL_EMIT_SEG: begin
        if (init_blank ? data_infifo_valid_in & (~data_infifo_eos_in) & blank_done_stick_sticky: data_infifo_valid_in & (~data_infifo_eos_in)) begin
          scan_seq_next_state = UL;
        end
        else if (spacc_mode ? data_done_in | (init_blank & (~blank_done_stick_sticky)) | stop_lvl_geq: data_done_in) begin
          scan_seq_next_state = FINALIZE1;
        end
        else scan_seq_next_state = UL_EMIT_SEG;
      end
    UL_WZ: begin
        if (&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full})) begin
          scan_seq_next_state = UL;
        end
        else if (~(&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}))) begin
          scan_seq_next_state = UL_WZ;
        end
      end
    UnLL: begin
        if ((data_done_in & addr_done_in) | (spacc_mode & stop_lvl_geq)) begin
          scan_seq_next_state = FINALIZE2;
        end
        else scan_seq_next_state = UnLL;
      end
    default: scan_seq_next_state = scan_seq_current_state;
  endcase
end
always_comb begin
  unique case (scan_seq_current_state)
    ALLOCATE1: begin :scan_seq_ALLOCATE1_Output
        data_to_fifo = 16'h0;
        op_to_fifo = 1'h0;
        addr_to_fifo = 16'h0;
        ID_to_fifo = 16'h0;
        push_to_outs = 1'h1;
        inc_seg_addr = 1'h0;
        clr_seg_addr = 1'h0;
        inc_coord_addr = 1'h0;
        clr_coord_addr = 1'h0;
        inc_seg_ctr = 1'h0;
        clr_seg_ctr = 1'h0;
        set_curr_coord = 1'h0;
        clr_curr_coord = 1'h0;
        infifo_pop[0] = 1'h0;
        infifo_pop[1] = 1'h0;
        clr_wen_made = 1'h0;
        set_block_size = 1'h0;
        inc_block_write = 1'h0;
        clr_block_write = 1'h0;
        clr_blank_done = 1'h0;
        set_blank_done = 1'h0;
        pop_block_wr = 1'h0;
      end :scan_seq_ALLOCATE1_Output
    ALLOCATE2: begin :scan_seq_ALLOCATE2_Output
        data_to_fifo = 16'h0;
        op_to_fifo = 1'h0;
        addr_to_fifo = 16'h0;
        ID_to_fifo = 16'h1;
        push_to_outs = 1'h1;
        inc_seg_addr = 1'h0;
        clr_seg_addr = 1'h0;
        inc_coord_addr = 1'h0;
        clr_coord_addr = 1'h0;
        inc_seg_ctr = 1'h0;
        clr_seg_ctr = 1'h0;
        set_curr_coord = 1'h0;
        clr_curr_coord = 1'h0;
        infifo_pop[0] = 1'h0;
        infifo_pop[1] = 1'h0;
        clr_wen_made = 1'h0;
        set_block_size = 1'h0;
        inc_block_write = 1'h0;
        clr_block_write = 1'h0;
        clr_blank_done = 1'h0;
        set_blank_done = 1'h0;
        pop_block_wr = 1'h0;
      end :scan_seq_ALLOCATE2_Output
    BLOCK_1_SZ: begin :scan_seq_BLOCK_1_SZ_Output
        data_to_fifo = 16'h0;
        op_to_fifo = 1'h0;
        addr_to_fifo = 16'h0;
        ID_to_fifo = 16'h1;
        push_to_outs = 1'h0;
        inc_seg_addr = 1'h0;
        clr_seg_addr = 1'h0;
        inc_coord_addr = 1'h0;
        clr_coord_addr = 1'h0;
        inc_seg_ctr = 1'h0;
        clr_seg_ctr = 1'h0;
        set_curr_coord = 1'h0;
        clr_curr_coord = 1'h0;
        infifo_pop[0] = 1'h0;
        infifo_pop[1] = 1'h0;
        clr_wen_made = 1'h0;
        set_block_size = block_wr_fifo_valid;
        inc_block_write = 1'h0;
        clr_block_write = 1'h1;
        pop_block_wr = block_wr_fifo_valid;
        clr_blank_done = 1'h0;
        set_blank_done = 1'h0;
      end :scan_seq_BLOCK_1_SZ_Output
    BLOCK_1_WR: begin :scan_seq_BLOCK_1_WR_Output
        data_to_fifo = block_wr_input_fifo_data_out;
        op_to_fifo = 1'h1;
        addr_to_fifo = block_write_count;
        ID_to_fifo = 16'h0;
        push_to_outs = block_wr_fifo_valid & (block_write_count < block_size);
        inc_seg_addr = 1'h0;
        clr_seg_addr = 1'h0;
        inc_coord_addr = 1'h0;
        clr_coord_addr = 1'h0;
        inc_seg_ctr = 1'h0;
        clr_seg_ctr = 1'h0;
        set_curr_coord = 1'h0;
        clr_curr_coord = 1'h0;
        infifo_pop[0] = 1'h0;
        infifo_pop[1] = 1'h0;
        clr_wen_made = 1'h0;
        set_block_size = 1'h0;
        inc_block_write = block_wr_fifo_valid & (block_write_count < block_size) &
            (&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}));
        clr_block_write = 1'h0;
        pop_block_wr = block_wr_fifo_valid & (block_write_count < block_size) &
            (&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}));
        clr_blank_done = 1'h0;
        set_blank_done = 1'h0;
      end :scan_seq_BLOCK_1_WR_Output
    BLOCK_2_SZ: begin :scan_seq_BLOCK_2_SZ_Output
        data_to_fifo = 16'h0;
        op_to_fifo = 1'h0;
        addr_to_fifo = 16'h0;
        ID_to_fifo = 16'h0;
        push_to_outs = 1'h0;
        inc_seg_addr = 1'h0;
        clr_seg_addr = 1'h0;
        inc_coord_addr = 1'h0;
        clr_coord_addr = 1'h0;
        inc_seg_ctr = 1'h0;
        clr_seg_ctr = 1'h0;
        set_curr_coord = 1'h0;
        clr_curr_coord = 1'h0;
        infifo_pop[0] = 1'h0;
        infifo_pop[1] = 1'h0;
        clr_wen_made = 1'h0;
        set_block_size = block_wr_fifo_valid;
        inc_block_write = 1'h0;
        clr_block_write = 1'h1;
        pop_block_wr = block_wr_fifo_valid;
        clr_blank_done = 1'h0;
        set_blank_done = 1'h0;
      end :scan_seq_BLOCK_2_SZ_Output
    BLOCK_2_WR: begin :scan_seq_BLOCK_2_WR_Output
        data_to_fifo = block_wr_input_fifo_data_out;
        op_to_fifo = 1'h1;
        addr_to_fifo = block_write_count;
        ID_to_fifo = 16'h1;
        push_to_outs = block_wr_fifo_valid & (block_write_count < block_size);
        inc_seg_addr = 1'h0;
        clr_seg_addr = 1'h0;
        inc_coord_addr = 1'h0;
        clr_coord_addr = 1'h0;
        inc_seg_ctr = 1'h0;
        clr_seg_ctr = 1'h0;
        set_curr_coord = 1'h0;
        clr_curr_coord = 1'h0;
        infifo_pop[0] = 1'h0;
        infifo_pop[1] = 1'h0;
        clr_wen_made = 1'h0;
        set_block_size = 1'h0;
        inc_block_write = block_wr_fifo_valid & (block_write_count < block_size) &
            (&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}));
        clr_block_write = 1'h0;
        pop_block_wr = block_wr_fifo_valid & (block_write_count < block_size) &
            (&(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full}));
        clr_blank_done = 1'h0;
        set_blank_done = 1'h0;
      end :scan_seq_BLOCK_2_WR_Output
    ComLL: begin :scan_seq_ComLL_Output
        data_to_fifo = data_infifo_data_in;
        op_to_fifo = 1'h1;
        addr_to_fifo = segment_addr;
        ID_to_fifo = 16'h0;
        push_to_outs = data_infifo_valid_in & (~data_infifo_eos_in);
        inc_seg_addr = data_infifo_valid_in & (~data_infifo_eos_in) & (&(~{data_out_fifo_full,
            addr_out_fifo_full, ID_out_fifo_full}));
        clr_seg_addr = 1'h0;
        inc_coord_addr = 1'h0;
        clr_coord_addr = 1'h0;
        inc_seg_ctr = 1'h0;
        clr_seg_ctr = 1'h0;
        set_curr_coord = 1'h0;
        clr_curr_coord = 1'h0;
        infifo_pop[0] = data_infifo_valid_in & (data_infifo_eos_in | (&(~{data_out_fifo_full,
            addr_out_fifo_full, ID_out_fifo_full})));
        infifo_pop[1] = 1'h0;
        clr_wen_made = 1'h0;
        set_block_size = 1'h0;
        inc_block_write = 1'h0;
        clr_block_write = 1'h0;
        clr_blank_done = 1'h0;
        set_blank_done = 1'h0;
        pop_block_wr = 1'h0;
      end :scan_seq_ComLL_Output
    DONE: begin :scan_seq_DONE_Output
        data_to_fifo = 16'h0;
        op_to_fifo = 1'h0;
        addr_to_fifo = 16'h0;
        ID_to_fifo = 16'h0;
        push_to_outs = 1'h0;
        inc_seg_addr = 1'h0;
        clr_seg_addr = 1'h0;
        inc_coord_addr = 1'h0;
        clr_coord_addr = 1'h0;
        inc_seg_ctr = 1'h0;
        clr_seg_ctr = 1'h0;
        set_curr_coord = 1'h0;
        clr_curr_coord = 1'h0;
        infifo_pop[0] = data_done_in;
        infifo_pop[1] = 1'h0;
        clr_wen_made = 1'h0;
        set_block_size = 1'h0;
        inc_block_write = 1'h0;
        clr_block_write = 1'h0;
        set_blank_done = init_blank & (~blank_done_stick_sticky) & spacc_mode;
        clr_blank_done = init_blank & blank_done_stick_sticky & stop_lvl_new_blank_sticky_sticky &
            spacc_mode;
        pop_block_wr = 1'h0;
      end :scan_seq_DONE_Output
    FINALIZE1: begin :scan_seq_FINALIZE1_Output
        data_to_fifo = 16'h0;
        op_to_fifo = 1'h0;
        addr_to_fifo = 16'h0;
        ID_to_fifo = 16'h1;
        push_to_outs = 1'h1;
        inc_seg_addr = 1'h0;
        clr_seg_addr = 1'h0;
        inc_coord_addr = 1'h0;
        clr_coord_addr = 1'h0;
        inc_seg_ctr = 1'h0;
        clr_seg_ctr = 1'h0;
        set_curr_coord = 1'h0;
        clr_curr_coord = 1'h0;
        infifo_pop[0] = 1'h0;
        infifo_pop[1] = 1'h0;
        clr_wen_made = 1'h0;
        set_block_size = 1'h0;
        inc_block_write = 1'h0;
        clr_block_write = 1'h0;
        clr_blank_done = 1'h0;
        set_blank_done = 1'h0;
        pop_block_wr = 1'h0;
      end :scan_seq_FINALIZE1_Output
    FINALIZE2: begin :scan_seq_FINALIZE2_Output
        data_to_fifo = 16'h0;
        op_to_fifo = 1'h0;
        addr_to_fifo = 16'h0;
        ID_to_fifo = 16'h0;
        push_to_outs = 1'h1;
        inc_seg_addr = 1'h0;
        clr_seg_addr = 1'h0;
        inc_coord_addr = 1'h0;
        clr_coord_addr = 1'h0;
        inc_seg_ctr = 1'h0;
        clr_seg_ctr = 1'h0;
        set_curr_coord = 1'h0;
        clr_curr_coord = 1'h0;
        infifo_pop[0] = 1'h0;
        infifo_pop[1] = 1'h0;
        clr_wen_made = 1'h0;
        set_block_size = 1'h0;
        inc_block_write = 1'h0;
        clr_block_write = 1'h0;
        clr_blank_done = 1'h0;
        set_blank_done = 1'h0;
        pop_block_wr = 1'h0;
      end :scan_seq_FINALIZE2_Output
    LL: begin :scan_seq_LL_Output
        data_to_fifo = 16'h0;
        op_to_fifo = 1'h0;
        addr_to_fifo = 16'h0;
        ID_to_fifo = 16'h0;
        push_to_outs = 1'h0;
        inc_seg_addr = 1'h0;
        clr_seg_addr = 1'h0;
        inc_coord_addr = 1'h0;
        clr_coord_addr = 1'h0;
        inc_seg_ctr = 1'h0;
        clr_seg_ctr = 1'h0;
        set_curr_coord = 1'h0;
        clr_curr_coord = 1'h0;
        infifo_pop[0] = 1'h0;
        infifo_pop[1] = 1'h0;
        clr_wen_made = 1'h0;
        set_block_size = 1'h0;
        inc_block_write = 1'h0;
        clr_block_write = 1'h0;
        clr_blank_done = 1'h0;
        set_blank_done = 1'h0;
        pop_block_wr = 1'h0;
      end :scan_seq_LL_Output
    START: begin :scan_seq_START_Output
        data_to_fifo = 16'h0;
        op_to_fifo = 1'h0;
        addr_to_fifo = 16'h0;
        ID_to_fifo = 16'h0;
        push_to_outs = 1'h0;
        inc_seg_addr = 1'h0;
        clr_seg_addr = 1'h1;
        inc_coord_addr = 1'h0;
        clr_coord_addr = 1'h1;
        inc_seg_ctr = 1'h0;
        clr_seg_ctr = 1'h1;
        set_curr_coord = 1'h0;
        clr_curr_coord = 1'h1;
        infifo_pop[0] = 1'h0;
        infifo_pop[1] = 1'h0;
        clr_wen_made = 1'h1;
        set_block_size = 1'h0;
        inc_block_write = 1'h0;
        clr_block_write = 1'h1;
        clr_blank_done = 1'h0;
        set_blank_done = 1'h0;
        pop_block_wr = 1'h0;
      end :scan_seq_START_Output
    UL: begin :scan_seq_UL_Output
        data_to_fifo = 16'h0;
        op_to_fifo = 1'h0;
        addr_to_fifo = 16'h0;
        ID_to_fifo = 16'h0;
        push_to_outs = 1'h0;
        inc_seg_addr = 1'h0;
        clr_seg_addr = 1'h0;
        inc_coord_addr = 1'h0;
        clr_coord_addr = 1'h0;
        inc_seg_ctr = 1'h0;
        clr_seg_ctr = 1'h0;
        set_curr_coord = new_coord;
        clr_curr_coord = 1'h0;
        infifo_pop[0] = 1'h0;
        infifo_pop[1] = 1'h0;
        clr_wen_made = 1'h1;
        set_block_size = 1'h0;
        inc_block_write = 1'h0;
        clr_block_write = 1'h0;
        clr_blank_done = 1'h0;
        set_blank_done = 1'h0;
        pop_block_wr = 1'h0;
      end :scan_seq_UL_Output
    UL_EMIT_COORD: begin :scan_seq_UL_EMIT_COORD_Output
        data_to_fifo = data_infifo_data_in_d1;
        op_to_fifo = 1'h1;
        addr_to_fifo = coord_addr;
        ID_to_fifo = 16'h1;
        push_to_outs = (~wen_made_sticky) & (&(~{data_out_fifo_full, addr_out_fifo_full,
            ID_out_fifo_full}));
        inc_seg_addr = 1'h0;
        clr_seg_addr = 1'h0;
        inc_coord_addr = (~wen_made_sticky) & (&(~{data_out_fifo_full, addr_out_fifo_full,
            ID_out_fifo_full}));
        clr_coord_addr = 1'h0;
        inc_seg_ctr = (~wen_made_sticky) & (&(~{data_out_fifo_full, addr_out_fifo_full,
            ID_out_fifo_full}));
        clr_seg_ctr = 1'h0;
        set_curr_coord = 1'h0;
        clr_curr_coord = 1'h0;
        infifo_pop[0] = (~new_coord) & (~stop_in);
        infifo_pop[1] = 1'h0;
        clr_wen_made = 1'h0;
        set_block_size = 1'h0;
        inc_block_write = 1'h0;
        clr_block_write = 1'h0;
        clr_blank_done = 1'h0;
        set_blank_done = 1'h0;
        pop_block_wr = 1'h0;
      end :scan_seq_UL_EMIT_COORD_Output
    UL_EMIT_SEG: begin :scan_seq_UL_EMIT_SEG_Output
        data_to_fifo = segment_counter;
        op_to_fifo = 1'h1;
        addr_to_fifo = segment_addr;
        ID_to_fifo = 16'h0;
        push_to_outs = (~wen_made_sticky) & (&(~{data_out_fifo_full, addr_out_fifo_full,
            ID_out_fifo_full}));
        inc_seg_addr = (~wen_made_sticky) & (&(~{data_out_fifo_full, addr_out_fifo_full,
            ID_out_fifo_full}));
        clr_seg_addr = 1'h0;
        inc_coord_addr = 1'h0;
        clr_coord_addr = 1'h0;
        inc_seg_ctr = 1'h0;
        clr_seg_ctr = 1'h0;
        set_curr_coord = 1'h0;
        clr_curr_coord = 1'h1;
        infifo_pop[0] = data_infifo_valid_in & data_infifo_eos_in & (~(init_blank &
            (~blank_done_stick_sticky))) & (~data_done_in);
        infifo_pop[1] = 1'h0;
        clr_wen_made = 1'h0;
        set_block_size = 1'h0;
        inc_block_write = 1'h0;
        clr_block_write = 1'h0;
        clr_blank_done = 1'h0;
        set_blank_done = 1'h0;
        pop_block_wr = 1'h0;
      end :scan_seq_UL_EMIT_SEG_Output
    UL_WZ: begin :scan_seq_UL_WZ_Output
        data_to_fifo = 16'h0;
        op_to_fifo = 1'h1;
        addr_to_fifo = segment_addr;
        ID_to_fifo = 16'h0;
        push_to_outs = 1'h1;
        inc_seg_addr = &(~{data_out_fifo_full, addr_out_fifo_full, ID_out_fifo_full});
        clr_seg_addr = 1'h0;
        inc_coord_addr = 1'h0;
        clr_coord_addr = 1'h0;
        inc_seg_ctr = 1'h0;
        clr_seg_ctr = 1'h0;
        set_curr_coord = 1'h0;
        clr_curr_coord = 1'h0;
        infifo_pop[0] = 1'h0;
        infifo_pop[1] = 1'h0;
        clr_wen_made = 1'h0;
        set_block_size = 1'h0;
        inc_block_write = 1'h0;
        clr_block_write = 1'h0;
        clr_blank_done = 1'h0;
        set_blank_done = 1'h0;
        pop_block_wr = 1'h0;
      end :scan_seq_UL_WZ_Output
    UnLL: begin :scan_seq_UnLL_Output
        data_to_fifo = data_infifo_data_in;
        op_to_fifo = 1'h1;
        addr_to_fifo = addr_infifo_data_in;
        ID_to_fifo = 16'h0;
        push_to_outs = data_infifo_valid_in & addr_infifo_valid_in & (~(data_infifo_eos_in |
            addr_infifo_eos_in));
        inc_seg_addr = 1'h0;
        clr_seg_addr = 1'h0;
        inc_coord_addr = 1'h0;
        clr_coord_addr = 1'h0;
        inc_seg_ctr = 1'h0;
        clr_seg_ctr = 1'h0;
        set_curr_coord = 1'h0;
        clr_curr_coord = 1'h0;
        infifo_pop[0] = data_infifo_valid_in & addr_infifo_valid_in & ((data_infifo_eos_in &
            addr_infifo_eos_in) | (&(~{data_out_fifo_full, addr_out_fifo_full,
            ID_out_fifo_full})));
        infifo_pop[1] = data_infifo_valid_in & addr_infifo_valid_in & ((data_infifo_eos_in &
            addr_infifo_eos_in) | (&(~{data_out_fifo_full, addr_out_fifo_full,
            ID_out_fifo_full})));
        clr_wen_made = 1'h0;
        set_block_size = 1'h0;
        inc_block_write = 1'h0;
        clr_block_write = 1'h0;
        clr_blank_done = 1'h0;
        set_blank_done = 1'h0;
        pop_block_wr = 1'h0;
      end :scan_seq_UnLL_Output
    default: begin :scan_seq_default_Output
        data_to_fifo = 16'h0;
        op_to_fifo = 1'h0;
        addr_to_fifo = 16'h0;
        ID_to_fifo = 16'h0;
        push_to_outs = 1'h0;
        inc_seg_addr = 1'h0;
        clr_seg_addr = 1'h1;
        inc_coord_addr = 1'h0;
        clr_coord_addr = 1'h1;
        inc_seg_ctr = 1'h0;
        clr_seg_ctr = 1'h1;
        set_curr_coord = 1'h0;
        clr_curr_coord = 1'h1;
        infifo_pop[0] = 1'h0;
        infifo_pop[1] = 1'h0;
        clr_wen_made = 1'h1;
        set_block_size = 1'h0;
        inc_block_write = 1'h0;
        clr_block_write = 1'h1;
        clr_blank_done = 1'h0;
        set_blank_done = 1'h0;
        pop_block_wr = 1'h0;
      end :scan_seq_default_Output
  endcase
end
reg_fifo_depth_0_w_17_afd_2 data_input_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(data_infifo_in_packed),
  .flush(flush),
  .pop(infifo_pop[0]),
  .push(data_in_valid),
  .rst_n(rst_n),
  .data_out(data_infifo_out_packed),
  .empty(data_input_fifo_empty),
  .full(data_input_fifo_full)
);

reg_fifo_depth_0_w_17_afd_2 addr_input_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(addr_infifo_in_packed),
  .flush(flush),
  .pop(infifo_pop[1]),
  .push(addr_in_valid),
  .rst_n(rst_n),
  .data_out(addr_infifo_out_packed),
  .empty(addr_input_fifo_empty),
  .full(addr_input_fifo_full)
);

reg_fifo_depth_0_w_16_afd_2 block_wr_input_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(block_wr_in[15:0]),
  .flush(flush),
  .pop(pop_block_wr),
  .push(block_wr_in_valid),
  .rst_n(rst_n),
  .data_out(block_wr_input_fifo_data_out),
  .empty(block_wr_input_fifo_empty),
  .full(block_wr_input_fifo_full)
);

reg_fifo_depth_2_w_17_afd_2 data_out_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(data_out_fifo_data_in),
  .flush(flush),
  .pop(data_out_ready),
  .push(data_out_fifo_push),
  .rst_n(rst_n),
  .data_out(data_out),
  .empty(data_out_fifo_empty),
  .full(data_out_fifo_full)
);

reg_fifo_depth_2_w_17_afd_2 addr_out_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(addr_out_fifo_data_in),
  .flush(flush),
  .pop(addr_out_ready),
  .push(addr_out_fifo_push),
  .rst_n(rst_n),
  .data_out(addr_out),
  .empty(addr_out_fifo_empty),
  .full(addr_out_fifo_full)
);

reg_fifo_depth_2_w_17_afd_2 ID_out_fifo (
  .clk(gclk),
  .clk_en(clk_en),
  .data_in(ID_out_fifo_data_in),
  .flush(flush),
  .pop(ID_out_ready),
  .push(ID_out_fifo_push),
  .rst_n(rst_n),
  .data_out(ID_out),
  .empty(ID_out_fifo_empty),
  .full(ID_out_fifo_full)
);

endmodule   // write_scanner


module FanoutHash_F95D10B01D02012 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[0]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[0]) | I3;
assign sel4 = (~E4) | (~S4[0]) | I4;
assign sel5 = (~E5) | (~S5[0]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_F95D10B01D02012


module FanoutHash_F8E7A0823DC8CDD (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[11]) | I3;
assign sel4 = (~E4) | (~S4[11]) | I4;
assign sel5 = (~E5) | (~S5[11]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_F8E7A0823DC8CDD


module FanoutHash_F689C91787363AB (
  input logic E0,
  input logic E1,
  input logic E10,
  input logic E11,
  input logic E12,
  input logic E13,
  input logic E14,
  input logic E15,
  input logic E16,
  input logic E17,
  input logic E18,
  input logic E19,
  input logic E2,
  input logic E20,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic E9,
  input logic I0,
  input logic I1,
  input logic I10,
  input logic I11,
  input logic I12,
  input logic I13,
  input logic I14,
  input logic I15,
  input logic I16,
  input logic I17,
  input logic I18,
  input logic I19,
  input logic I2,
  input logic I20,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic I9,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S10,
  input logic [7:0] S11,
  input logic [7:0] S12,
  input logic [7:0] S13,
  input logic [7:0] S14,
  input logic [7:0] S15,
  input logic [7:0] S16,
  input logic [7:0] S17,
  input logic [7:0] S18,
  input logic [7:0] S19,
  input logic [7:0] S2,
  input logic [31:0] S20,
  input logic [7:0] S3,
  input logic [7:0] S4,
  input logic [7:0] S5,
  input logic [7:0] S6,
  input logic [7:0] S7,
  input logic [7:0] S8,
  input logic [7:0] S9,
  output logic O
);

logic sel0;
logic sel1;
logic sel10;
logic sel11;
logic sel12;
logic sel13;
logic sel14;
logic sel15;
logic sel16;
logic sel17;
logic sel18;
logic sel19;
logic sel2;
logic sel20;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
logic sel9;
assign sel0 = (~E0) | (~S0[4]) | I0;
assign sel1 = (~E1) | (~S1[4]) | I1;
assign sel2 = (~E2) | (~S2[4]) | I2;
assign sel3 = (~E3) | (~S3[4]) | I3;
assign sel4 = (~E4) | (~S4[4]) | I4;
assign sel5 = (~E5) | (~S5[4]) | I5;
assign sel6 = (~E6) | (~S6[4]) | I6;
assign sel7 = (~E7) | (~S7[4]) | I7;
assign sel8 = (~E8) | (~S8[4]) | I8;
assign sel9 = (~E9) | (~S9[4]) | I9;
assign sel10 = (~E10) | (~S10[4]) | I10;
assign sel11 = (~E11) | (~S11[4]) | I11;
assign sel12 = (~E12) | (~S12[4]) | I12;
assign sel13 = (~E13) | (~S13[4]) | I13;
assign sel14 = (~E14) | (~S14[4]) | I14;
assign sel15 = (~E15) | (~S15[4]) | I15;
assign sel16 = (~E16) | (~S16[4]) | I16;
assign sel17 = (~E17) | (~S17[4]) | I17;
assign sel18 = (~E18) | (~S18[4]) | I18;
assign sel19 = (~E19) | (~S19[4]) | I19;
assign sel20 = (~E20) | (~S20[20]) | I20;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8 & sel9 & sel10 &
    sel11 & sel12 & sel13 & sel14 & sel15 & sel16 & sel17 & sel18 & sel19 & sel20;
endmodule   // FanoutHash_F689C91787363AB


module FanoutHash_E70AF988E4250F5 (
  input logic E0,
  input logic E1,
  input logic E10,
  input logic E11,
  input logic E12,
  input logic E13,
  input logic E14,
  input logic E15,
  input logic E16,
  input logic E17,
  input logic E18,
  input logic E19,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic E9,
  input logic I0,
  input logic I1,
  input logic I10,
  input logic I11,
  input logic I12,
  input logic I13,
  input logic I14,
  input logic I15,
  input logic I16,
  input logic I17,
  input logic I18,
  input logic I19,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic I9,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S10,
  input logic [7:0] S11,
  input logic [7:0] S12,
  input logic [7:0] S13,
  input logic [7:0] S14,
  input logic [7:0] S15,
  input logic [7:0] S16,
  input logic [7:0] S17,
  input logic [7:0] S18,
  input logic [7:0] S19,
  input logic [7:0] S2,
  input logic [7:0] S3,
  input logic [7:0] S4,
  input logic [7:0] S5,
  input logic [7:0] S6,
  input logic [7:0] S7,
  input logic [7:0] S8,
  input logic [7:0] S9,
  output logic O
);

logic sel0;
logic sel1;
logic sel10;
logic sel11;
logic sel12;
logic sel13;
logic sel14;
logic sel15;
logic sel16;
logic sel17;
logic sel18;
logic sel19;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
logic sel9;
assign sel0 = (~E0) | (~S0[3]) | I0;
assign sel1 = (~E1) | (~S1[3]) | I1;
assign sel2 = (~E2) | (~S2[3]) | I2;
assign sel3 = (~E3) | (~S3[3]) | I3;
assign sel4 = (~E4) | (~S4[3]) | I4;
assign sel5 = (~E5) | (~S5[3]) | I5;
assign sel6 = (~E6) | (~S6[3]) | I6;
assign sel7 = (~E7) | (~S7[3]) | I7;
assign sel8 = (~E8) | (~S8[3]) | I8;
assign sel9 = (~E9) | (~S9[3]) | I9;
assign sel10 = (~E10) | (~S10[3]) | I10;
assign sel11 = (~E11) | (~S11[3]) | I11;
assign sel12 = (~E12) | (~S12[3]) | I12;
assign sel13 = (~E13) | (~S13[3]) | I13;
assign sel14 = (~E14) | (~S14[3]) | I14;
assign sel15 = (~E15) | (~S15[3]) | I15;
assign sel16 = (~E16) | (~S16[3]) | I16;
assign sel17 = (~E17) | (~S17[3]) | I17;
assign sel18 = (~E18) | (~S18[3]) | I18;
assign sel19 = (~E19) | (~S19[3]) | I19;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8 & sel9 & sel10 &
    sel11 & sel12 & sel13 & sel14 & sel15 & sel16 & sel17 & sel18 & sel19;
endmodule   // FanoutHash_E70AF988E4250F5


module FanoutHash_D70CFBE8EA3CE7F (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[0]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[14]) | I3;
assign sel4 = (~E4) | (~S4[14]) | I4;
assign sel5 = (~E5) | (~S5[14]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_D70CFBE8EA3CE7F


module FanoutHash_CE1AA874B742213 (
  input logic E0,
  input logic E1,
  input logic E10,
  input logic E11,
  input logic E12,
  input logic E13,
  input logic E14,
  input logic E15,
  input logic E16,
  input logic E17,
  input logic E18,
  input logic E19,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic E9,
  input logic I0,
  input logic I1,
  input logic I10,
  input logic I11,
  input logic I12,
  input logic I13,
  input logic I14,
  input logic I15,
  input logic I16,
  input logic I17,
  input logic I18,
  input logic I19,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic I9,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S10,
  input logic [7:0] S11,
  input logic [7:0] S12,
  input logic [7:0] S13,
  input logic [7:0] S14,
  input logic [7:0] S15,
  input logic [7:0] S16,
  input logic [7:0] S17,
  input logic [7:0] S18,
  input logic [7:0] S19,
  input logic [7:0] S2,
  input logic [7:0] S3,
  input logic [7:0] S4,
  input logic [7:0] S5,
  input logic [7:0] S6,
  input logic [7:0] S7,
  input logic [7:0] S8,
  input logic [7:0] S9,
  output logic O
);

logic sel0;
logic sel1;
logic sel10;
logic sel11;
logic sel12;
logic sel13;
logic sel14;
logic sel15;
logic sel16;
logic sel17;
logic sel18;
logic sel19;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
logic sel9;
assign sel0 = (~E0) | (~S0[5]) | I0;
assign sel1 = (~E1) | (~S1[5]) | I1;
assign sel2 = (~E2) | (~S2[5]) | I2;
assign sel3 = (~E3) | (~S3[5]) | I3;
assign sel4 = (~E4) | (~S4[5]) | I4;
assign sel5 = (~E5) | (~S5[5]) | I5;
assign sel6 = (~E6) | (~S6[5]) | I6;
assign sel7 = (~E7) | (~S7[5]) | I7;
assign sel8 = (~E8) | (~S8[5]) | I8;
assign sel9 = (~E9) | (~S9[5]) | I9;
assign sel10 = (~E10) | (~S10[5]) | I10;
assign sel11 = (~E11) | (~S11[5]) | I11;
assign sel12 = (~E12) | (~S12[5]) | I12;
assign sel13 = (~E13) | (~S13[5]) | I13;
assign sel14 = (~E14) | (~S14[5]) | I14;
assign sel15 = (~E15) | (~S15[5]) | I15;
assign sel16 = (~E16) | (~S16[5]) | I16;
assign sel17 = (~E17) | (~S17[5]) | I17;
assign sel18 = (~E18) | (~S18[5]) | I18;
assign sel19 = (~E19) | (~S19[5]) | I19;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8 & sel9 & sel10 &
    sel11 & sel12 & sel13 & sel14 & sel15 & sel16 & sel17 & sel18 & sel19;
endmodule   // FanoutHash_CE1AA874B742213


module FanoutHash_AE7392256DF8B0F (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[17]) | I3;
assign sel4 = (~E4) | (~S4[17]) | I4;
assign sel5 = (~E5) | (~S5[17]) | I5;
assign sel6 = (~E6) | (~S6[17]) | I6;
assign sel7 = (~E7) | (~S7[17]) | I7;
assign sel8 = (~E8) | (~S8[17]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_AE7392256DF8B0F


module FanoutHash_99D793215CEDDD5 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[1]) | I3;
assign sel4 = (~E4) | (~S4[1]) | I4;
assign sel5 = (~E5) | (~S5[1]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_99D793215CEDDD5


module FanoutHash_87642A353688B49 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[0]) | I1;
assign sel2 = (~E2) | (~S2[0]) | I2;
assign sel3 = (~E3) | (~S3[3]) | I3;
assign sel4 = (~E4) | (~S4[3]) | I4;
assign sel5 = (~E5) | (~S5[3]) | I5;
assign sel6 = (~E6) | (~S6[3]) | I6;
assign sel7 = (~E7) | (~S7[3]) | I7;
assign sel8 = (~E8) | (~S8[3]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_87642A353688B49


module FanoutHash_82899D6851EDC11 (
  input logic E0,
  input logic E1,
  input logic E10,
  input logic E11,
  input logic E12,
  input logic E13,
  input logic E14,
  input logic E15,
  input logic E16,
  input logic E17,
  input logic E18,
  input logic E19,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic E9,
  input logic I0,
  input logic I1,
  input logic I10,
  input logic I11,
  input logic I12,
  input logic I13,
  input logic I14,
  input logic I15,
  input logic I16,
  input logic I17,
  input logic I18,
  input logic I19,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic I9,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S10,
  input logic [7:0] S11,
  input logic [7:0] S12,
  input logic [7:0] S13,
  input logic [7:0] S14,
  input logic [7:0] S15,
  input logic [7:0] S16,
  input logic [7:0] S17,
  input logic [7:0] S18,
  input logic [7:0] S19,
  input logic [7:0] S2,
  input logic [7:0] S3,
  input logic [7:0] S4,
  input logic [7:0] S5,
  input logic [7:0] S6,
  input logic [7:0] S7,
  input logic [7:0] S8,
  input logic [7:0] S9,
  output logic O
);

logic sel0;
logic sel1;
logic sel10;
logic sel11;
logic sel12;
logic sel13;
logic sel14;
logic sel15;
logic sel16;
logic sel17;
logic sel18;
logic sel19;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
logic sel9;
assign sel0 = (~E0) | (~S0[4]) | I0;
assign sel1 = (~E1) | (~S1[4]) | I1;
assign sel2 = (~E2) | (~S2[4]) | I2;
assign sel3 = (~E3) | (~S3[4]) | I3;
assign sel4 = (~E4) | (~S4[4]) | I4;
assign sel5 = (~E5) | (~S5[4]) | I5;
assign sel6 = (~E6) | (~S6[4]) | I6;
assign sel7 = (~E7) | (~S7[4]) | I7;
assign sel8 = (~E8) | (~S8[4]) | I8;
assign sel9 = (~E9) | (~S9[4]) | I9;
assign sel10 = (~E10) | (~S10[4]) | I10;
assign sel11 = (~E11) | (~S11[4]) | I11;
assign sel12 = (~E12) | (~S12[4]) | I12;
assign sel13 = (~E13) | (~S13[4]) | I13;
assign sel14 = (~E14) | (~S14[4]) | I14;
assign sel15 = (~E15) | (~S15[4]) | I15;
assign sel16 = (~E16) | (~S16[4]) | I16;
assign sel17 = (~E17) | (~S17[4]) | I17;
assign sel18 = (~E18) | (~S18[4]) | I18;
assign sel19 = (~E19) | (~S19[4]) | I19;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8 & sel9 & sel10 &
    sel11 & sel12 & sel13 & sel14 & sel15 & sel16 & sel17 & sel18 & sel19;
endmodule   // FanoutHash_82899D6851EDC11


module FanoutHash_7FDF2D3240D4A947 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[2]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[15]) | I3;
assign sel4 = (~E4) | (~S4[15]) | I4;
assign sel5 = (~E5) | (~S5[15]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_7FDF2D3240D4A947


module FanoutHash_7F4660D1463D9234 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[0]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[10]) | I3;
assign sel4 = (~E4) | (~S4[10]) | I4;
assign sel5 = (~E5) | (~S5[10]) | I5;
assign sel6 = (~E6) | (~S6[10]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_7F4660D1463D9234


module FanoutHash_7ED1C80229B84786 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[7]) | I3;
assign sel4 = (~E4) | (~S4[7]) | I4;
assign sel5 = (~E5) | (~S5[7]) | I5;
assign sel6 = (~E6) | (~S6[7]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_7ED1C80229B84786


module FanoutHash_7E22D83B42537D1D (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[0]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[12]) | I3;
assign sel4 = (~E4) | (~S4[12]) | I4;
assign sel5 = (~E5) | (~S5[12]) | I5;
assign sel6 = (~E6) | (~S6[12]) | I6;
assign sel7 = (~E7) | (~S7[12]) | I7;
assign sel8 = (~E8) | (~S8[12]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_7E22D83B42537D1D


module FanoutHash_752C11B748DD905C (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[11]) | I3;
assign sel4 = (~E4) | (~S4[11]) | I4;
assign sel5 = (~E5) | (~S5[11]) | I5;
assign sel6 = (~E6) | (~S6[11]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_752C11B748DD905C


module FanoutHash_74A3E41836ECED62 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[0]) | I2;
assign sel3 = (~E3) | (~S3[8]) | I3;
assign sel4 = (~E4) | (~S4[8]) | I4;
assign sel5 = (~E5) | (~S5[8]) | I5;
assign sel6 = (~E6) | (~S6[8]) | I6;
assign sel7 = (~E7) | (~S7[8]) | I7;
assign sel8 = (~E8) | (~S8[8]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_74A3E41836ECED62


module FanoutHash_6EB42FA08A9B7B5B (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[0]) | I2;
assign sel3 = (~E3) | (~S3[8]) | I3;
assign sel4 = (~E4) | (~S4[8]) | I4;
assign sel5 = (~E5) | (~S5[8]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_6EB42FA08A9B7B5B


module FanoutHash_6E1094CE0D0F6DFA (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[2]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[19]) | I3;
assign sel4 = (~E4) | (~S4[19]) | I4;
assign sel5 = (~E5) | (~S5[19]) | I5;
assign sel6 = (~E6) | (~S6[19]) | I6;
assign sel7 = (~E7) | (~S7[19]) | I7;
assign sel8 = (~E8) | (~S8[19]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_6E1094CE0D0F6DFA


module FanoutHash_69376833A2418E2 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[0]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[12]) | I3;
assign sel4 = (~E4) | (~S4[12]) | I4;
assign sel5 = (~E5) | (~S5[12]) | I5;
assign sel6 = (~E6) | (~S6[12]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_69376833A2418E2


module FanoutHash_66A75CC8494A4D6B (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[13]) | I3;
assign sel4 = (~E4) | (~S4[13]) | I4;
assign sel5 = (~E5) | (~S5[13]) | I5;
assign sel6 = (~E6) | (~S6[13]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_66A75CC8494A4D6B


module FanoutHash_660E59B0DDACF452 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[2]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[19]) | I3;
assign sel4 = (~E4) | (~S4[19]) | I4;
assign sel5 = (~E5) | (~S5[19]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_660E59B0DDACF452


module FanoutHash_65A468071775C7BB (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[0]) | I1;
assign sel2 = (~E2) | (~S2[0]) | I2;
assign sel3 = (~E3) | (~S3[3]) | I3;
assign sel4 = (~E4) | (~S4[3]) | I4;
assign sel5 = (~E5) | (~S5[3]) | I5;
assign sel6 = (~E6) | (~S6[3]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_65A468071775C7BB


module FanoutHash_653384C8EF52B5E3 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[7]) | I3;
assign sel4 = (~E4) | (~S4[7]) | I4;
assign sel5 = (~E5) | (~S5[7]) | I5;
assign sel6 = (~E6) | (~S6[7]) | I6;
assign sel7 = (~E7) | (~S7[7]) | I7;
assign sel8 = (~E8) | (~S8[7]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_653384C8EF52B5E3


module FanoutHash_5DE101F5B6936D07 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[0]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[12]) | I3;
assign sel4 = (~E4) | (~S4[12]) | I4;
assign sel5 = (~E5) | (~S5[12]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_5DE101F5B6936D07


module FanoutHash_5D7AEC1255CDC1CC (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[18]) | I3;
assign sel4 = (~E4) | (~S4[18]) | I4;
assign sel5 = (~E5) | (~S5[18]) | I5;
assign sel6 = (~E6) | (~S6[18]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_5D7AEC1255CDC1CC


module FanoutHash_5CD8077D054B887B (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[0]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[10]) | I3;
assign sel4 = (~E4) | (~S4[10]) | I4;
assign sel5 = (~E5) | (~S5[10]) | I5;
assign sel6 = (~E6) | (~S6[10]) | I6;
assign sel7 = (~E7) | (~S7[10]) | I7;
assign sel8 = (~E8) | (~S8[10]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_5CD8077D054B887B


module FanoutHash_59B7E37DAE2221E3 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[13]) | I3;
assign sel4 = (~E4) | (~S4[13]) | I4;
assign sel5 = (~E5) | (~S5[13]) | I5;
assign sel6 = (~E6) | (~S6[13]) | I6;
assign sel7 = (~E7) | (~S7[13]) | I7;
assign sel8 = (~E8) | (~S8[13]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_59B7E37DAE2221E3


module FanoutHash_55B00FA90A0098BB (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[2]) | I0;
assign sel1 = (~E1) | (~S1[0]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[2]) | I3;
assign sel4 = (~E4) | (~S4[2]) | I4;
assign sel5 = (~E5) | (~S5[2]) | I5;
assign sel6 = (~E6) | (~S6[2]) | I6;
assign sel7 = (~E7) | (~S7[2]) | I7;
assign sel8 = (~E8) | (~S8[2]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_55B00FA90A0098BB


module FanoutHash_55169EB19E10AA09 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[18]) | I3;
assign sel4 = (~E4) | (~S4[18]) | I4;
assign sel5 = (~E5) | (~S5[18]) | I5;
assign sel6 = (~E6) | (~S6[18]) | I6;
assign sel7 = (~E7) | (~S7[18]) | I7;
assign sel8 = (~E8) | (~S8[18]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_55169EB19E10AA09


module FanoutHash_4FF010386DB0B737 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[5]) | I3;
assign sel4 = (~E4) | (~S4[5]) | I4;
assign sel5 = (~E5) | (~S5[5]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_4FF010386DB0B737


module FanoutHash_4FADDC8F90390680 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[0]) | I2;
assign sel3 = (~E3) | (~S3[4]) | I3;
assign sel4 = (~E4) | (~S4[4]) | I4;
assign sel5 = (~E5) | (~S5[4]) | I5;
assign sel6 = (~E6) | (~S6[4]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_4FADDC8F90390680


module FanoutHash_4F83851A40824F89 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[0]) | I2;
assign sel3 = (~E3) | (~S3[6]) | I3;
assign sel4 = (~E4) | (~S4[6]) | I4;
assign sel5 = (~E5) | (~S5[6]) | I5;
assign sel6 = (~E6) | (~S6[6]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_4F83851A40824F89


module FanoutHash_4A74B16B611BA7E4 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[11]) | I3;
assign sel4 = (~E4) | (~S4[11]) | I4;
assign sel5 = (~E5) | (~S5[11]) | I5;
assign sel6 = (~E6) | (~S6[11]) | I6;
assign sel7 = (~E7) | (~S7[11]) | I7;
assign sel8 = (~E8) | (~S8[11]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_4A74B16B611BA7E4


module FanoutHash_47712AAC902ADA2 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[0]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[0]) | I3;
assign sel4 = (~E4) | (~S4[0]) | I4;
assign sel5 = (~E5) | (~S5[0]) | I5;
assign sel6 = (~E6) | (~S6[0]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_47712AAC902ADA2


module FanoutHash_4678C6877F96240E (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[2]) | I0;
assign sel1 = (~E1) | (~S1[0]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[2]) | I3;
assign sel4 = (~E4) | (~S4[2]) | I4;
assign sel5 = (~E5) | (~S5[2]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_4678C6877F96240E


module FanoutHash_466EB88CFD0CAD7B (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[5]) | I3;
assign sel4 = (~E4) | (~S4[5]) | I4;
assign sel5 = (~E5) | (~S5[5]) | I5;
assign sel6 = (~E6) | (~S6[5]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_466EB88CFD0CAD7B


module FanoutHash_43D5C80ABD816837 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[0]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[14]) | I3;
assign sel4 = (~E4) | (~S4[14]) | I4;
assign sel5 = (~E5) | (~S5[14]) | I5;
assign sel6 = (~E6) | (~S6[14]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_43D5C80ABD816837


module FanoutHash_41D739158D58E184 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[2]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[15]) | I3;
assign sel4 = (~E4) | (~S4[15]) | I4;
assign sel5 = (~E5) | (~S5[15]) | I5;
assign sel6 = (~E6) | (~S6[15]) | I6;
assign sel7 = (~E7) | (~S7[15]) | I7;
assign sel8 = (~E8) | (~S8[15]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_41D739158D58E184


module FanoutHash_3E05574A9CE9CA8A (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[1]) | I3;
assign sel4 = (~E4) | (~S4[1]) | I4;
assign sel5 = (~E5) | (~S5[1]) | I5;
assign sel6 = (~E6) | (~S6[1]) | I6;
assign sel7 = (~E7) | (~S7[1]) | I7;
assign sel8 = (~E8) | (~S8[1]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_3E05574A9CE9CA8A


module FanoutHash_3B67229CB02928BA (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[0]) | I2;
assign sel3 = (~E3) | (~S3[8]) | I3;
assign sel4 = (~E4) | (~S4[8]) | I4;
assign sel5 = (~E5) | (~S5[8]) | I5;
assign sel6 = (~E6) | (~S6[8]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_3B67229CB02928BA


module FanoutHash_3A6A5822E84DCC71 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[0]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[0]) | I3;
assign sel4 = (~E4) | (~S4[0]) | I4;
assign sel5 = (~E5) | (~S5[0]) | I5;
assign sel6 = (~E6) | (~S6[0]) | I6;
assign sel7 = (~E7) | (~S7[0]) | I7;
assign sel8 = (~E8) | (~S8[0]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_3A6A5822E84DCC71


module FanoutHash_3A0064632A577CF5 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[0]) | I1;
assign sel2 = (~E2) | (~S2[0]) | I2;
assign sel3 = (~E3) | (~S3[3]) | I3;
assign sel4 = (~E4) | (~S4[3]) | I4;
assign sel5 = (~E5) | (~S5[3]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_3A0064632A577CF5


module FanoutHash_37E9FE88073C5BAC (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[0]) | I2;
assign sel3 = (~E3) | (~S3[4]) | I3;
assign sel4 = (~E4) | (~S4[4]) | I4;
assign sel5 = (~E5) | (~S5[4]) | I5;
assign sel6 = (~E6) | (~S6[4]) | I6;
assign sel7 = (~E7) | (~S7[4]) | I7;
assign sel8 = (~E8) | (~S8[4]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_37E9FE88073C5BAC


module FanoutHash_37B926A0CDF82FCC (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[16]) | I3;
assign sel4 = (~E4) | (~S4[16]) | I4;
assign sel5 = (~E5) | (~S5[16]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_37B926A0CDF82FCC


module FanoutHash_330DF95D65589621 (
  input logic E0,
  input logic E1,
  input logic E10,
  input logic E11,
  input logic E12,
  input logic E13,
  input logic E14,
  input logic E15,
  input logic E16,
  input logic E17,
  input logic E18,
  input logic E19,
  input logic E2,
  input logic E20,
  input logic E21,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic E9,
  input logic I0,
  input logic I1,
  input logic I10,
  input logic I11,
  input logic I12,
  input logic I13,
  input logic I14,
  input logic I15,
  input logic I16,
  input logic I17,
  input logic I18,
  input logic I19,
  input logic I2,
  input logic I20,
  input logic I21,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic I9,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S10,
  input logic [7:0] S11,
  input logic [7:0] S12,
  input logic [7:0] S13,
  input logic [7:0] S14,
  input logic [7:0] S15,
  input logic [7:0] S16,
  input logic [7:0] S17,
  input logic [7:0] S18,
  input logic [7:0] S19,
  input logic [7:0] S2,
  input logic [31:0] S20,
  input logic [31:0] S21,
  input logic [7:0] S3,
  input logic [7:0] S4,
  input logic [7:0] S5,
  input logic [7:0] S6,
  input logic [7:0] S7,
  input logic [7:0] S8,
  input logic [7:0] S9,
  output logic O
);

logic sel0;
logic sel1;
logic sel10;
logic sel11;
logic sel12;
logic sel13;
logic sel14;
logic sel15;
logic sel16;
logic sel17;
logic sel18;
logic sel19;
logic sel2;
logic sel20;
logic sel21;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
logic sel9;
assign sel0 = (~E0) | (~S0[3]) | I0;
assign sel1 = (~E1) | (~S1[3]) | I1;
assign sel2 = (~E2) | (~S2[3]) | I2;
assign sel3 = (~E3) | (~S3[3]) | I3;
assign sel4 = (~E4) | (~S4[3]) | I4;
assign sel5 = (~E5) | (~S5[3]) | I5;
assign sel6 = (~E6) | (~S6[3]) | I6;
assign sel7 = (~E7) | (~S7[3]) | I7;
assign sel8 = (~E8) | (~S8[3]) | I8;
assign sel9 = (~E9) | (~S9[3]) | I9;
assign sel10 = (~E10) | (~S10[3]) | I10;
assign sel11 = (~E11) | (~S11[3]) | I11;
assign sel12 = (~E12) | (~S12[3]) | I12;
assign sel13 = (~E13) | (~S13[3]) | I13;
assign sel14 = (~E14) | (~S14[3]) | I14;
assign sel15 = (~E15) | (~S15[3]) | I15;
assign sel16 = (~E16) | (~S16[3]) | I16;
assign sel17 = (~E17) | (~S17[3]) | I17;
assign sel18 = (~E18) | (~S18[3]) | I18;
assign sel19 = (~E19) | (~S19[3]) | I19;
assign sel20 = (~E20) | (~S20[20]) | I20;
assign sel21 = (~E21) | (~S21[20]) | I21;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8 & sel9 & sel10 &
    sel11 & sel12 & sel13 & sel14 & sel15 & sel16 & sel17 & sel18 & sel19 & sel20 &
    sel21;
endmodule   // FanoutHash_330DF95D65589621


module FanoutHash_31AE65CCDD94603 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[2]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[15]) | I3;
assign sel4 = (~E4) | (~S4[15]) | I4;
assign sel5 = (~E5) | (~S5[15]) | I5;
assign sel6 = (~E6) | (~S6[15]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_31AE65CCDD94603


module FanoutHash_31555E0CDC460B97 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[0]) | I2;
assign sel3 = (~E3) | (~S3[4]) | I3;
assign sel4 = (~E4) | (~S4[4]) | I4;
assign sel5 = (~E5) | (~S5[4]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_31555E0CDC460B97


module FanoutHash_308BAC760F688049 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[2]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[9]) | I3;
assign sel4 = (~E4) | (~S4[9]) | I4;
assign sel5 = (~E5) | (~S5[9]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_308BAC760F688049


module FanoutHash_302974B49BE3F0C4 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[2]) | I0;
assign sel1 = (~E1) | (~S1[0]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[2]) | I3;
assign sel4 = (~E4) | (~S4[2]) | I4;
assign sel5 = (~E5) | (~S5[2]) | I5;
assign sel6 = (~E6) | (~S6[2]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_302974B49BE3F0C4


module FanoutHash_2F92967E9F56D548 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[5]) | I3;
assign sel4 = (~E4) | (~S4[5]) | I4;
assign sel5 = (~E5) | (~S5[5]) | I5;
assign sel6 = (~E6) | (~S6[5]) | I6;
assign sel7 = (~E7) | (~S7[5]) | I7;
assign sel8 = (~E8) | (~S8[5]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_2F92967E9F56D548


module FanoutHash_2CE3041FDDDDEC1A (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[2]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[9]) | I3;
assign sel4 = (~E4) | (~S4[9]) | I4;
assign sel5 = (~E5) | (~S5[9]) | I5;
assign sel6 = (~E6) | (~S6[9]) | I6;
assign sel7 = (~E7) | (~S7[9]) | I7;
assign sel8 = (~E8) | (~S8[9]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_2CE3041FDDDDEC1A


module FanoutHash_28125A548B305607 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[2]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[9]) | I3;
assign sel4 = (~E4) | (~S4[9]) | I4;
assign sel5 = (~E5) | (~S5[9]) | I5;
assign sel6 = (~E6) | (~S6[9]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_28125A548B305607


module FanoutHash_2785CE916183C5C (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[1]) | I3;
assign sel4 = (~E4) | (~S4[1]) | I4;
assign sel5 = (~E5) | (~S5[1]) | I5;
assign sel6 = (~E6) | (~S6[1]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_2785CE916183C5C


module FanoutHash_278348DB702230E6 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[0]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[10]) | I3;
assign sel4 = (~E4) | (~S4[10]) | I4;
assign sel5 = (~E5) | (~S5[10]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_278348DB702230E6


module FanoutHash_276F8381CE025648 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[0]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[14]) | I3;
assign sel4 = (~E4) | (~S4[14]) | I4;
assign sel5 = (~E5) | (~S5[14]) | I5;
assign sel6 = (~E6) | (~S6[14]) | I6;
assign sel7 = (~E7) | (~S7[14]) | I7;
assign sel8 = (~E8) | (~S8[14]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_276F8381CE025648


module FanoutHash_26B6474864379B6A (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[17]) | I3;
assign sel4 = (~E4) | (~S4[17]) | I4;
assign sel5 = (~E5) | (~S5[17]) | I5;
assign sel6 = (~E6) | (~S6[17]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_26B6474864379B6A


module FanoutHash_245560850976C879 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[0]) | I2;
assign sel3 = (~E3) | (~S3[6]) | I3;
assign sel4 = (~E4) | (~S4[6]) | I4;
assign sel5 = (~E5) | (~S5[6]) | I5;
assign sel6 = (~E6) | (~S6[6]) | I6;
assign sel7 = (~E7) | (~S7[6]) | I7;
assign sel8 = (~E8) | (~S8[6]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_245560850976C879


module FanoutHash_244497FCED8BEB80 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[16]) | I3;
assign sel4 = (~E4) | (~S4[16]) | I4;
assign sel5 = (~E5) | (~S5[16]) | I5;
assign sel6 = (~E6) | (~S6[16]) | I6;
assign sel7 = (~E7) | (~S7[16]) | I7;
assign sel8 = (~E8) | (~S8[16]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_244497FCED8BEB80


module FanoutHash_1EBD0270673B29D7 (
  input logic E0,
  input logic E1,
  input logic E10,
  input logic E11,
  input logic E12,
  input logic E13,
  input logic E14,
  input logic E15,
  input logic E16,
  input logic E17,
  input logic E18,
  input logic E19,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic E9,
  input logic I0,
  input logic I1,
  input logic I10,
  input logic I11,
  input logic I12,
  input logic I13,
  input logic I14,
  input logic I15,
  input logic I16,
  input logic I17,
  input logic I18,
  input logic I19,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic I9,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S10,
  input logic [7:0] S11,
  input logic [7:0] S12,
  input logic [7:0] S13,
  input logic [7:0] S14,
  input logic [7:0] S15,
  input logic [7:0] S16,
  input logic [7:0] S17,
  input logic [7:0] S18,
  input logic [7:0] S19,
  input logic [7:0] S2,
  input logic [7:0] S3,
  input logic [7:0] S4,
  input logic [7:0] S5,
  input logic [7:0] S6,
  input logic [7:0] S7,
  input logic [7:0] S8,
  input logic [7:0] S9,
  output logic O
);

logic sel0;
logic sel1;
logic sel10;
logic sel11;
logic sel12;
logic sel13;
logic sel14;
logic sel15;
logic sel16;
logic sel17;
logic sel18;
logic sel19;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
logic sel9;
assign sel0 = (~E0) | (~S0[6]) | I0;
assign sel1 = (~E1) | (~S1[6]) | I1;
assign sel2 = (~E2) | (~S2[6]) | I2;
assign sel3 = (~E3) | (~S3[6]) | I3;
assign sel4 = (~E4) | (~S4[6]) | I4;
assign sel5 = (~E5) | (~S5[6]) | I5;
assign sel6 = (~E6) | (~S6[6]) | I6;
assign sel7 = (~E7) | (~S7[6]) | I7;
assign sel8 = (~E8) | (~S8[6]) | I8;
assign sel9 = (~E9) | (~S9[6]) | I9;
assign sel10 = (~E10) | (~S10[6]) | I10;
assign sel11 = (~E11) | (~S11[6]) | I11;
assign sel12 = (~E12) | (~S12[6]) | I12;
assign sel13 = (~E13) | (~S13[6]) | I13;
assign sel14 = (~E14) | (~S14[6]) | I14;
assign sel15 = (~E15) | (~S15[6]) | I15;
assign sel16 = (~E16) | (~S16[6]) | I16;
assign sel17 = (~E17) | (~S17[6]) | I17;
assign sel18 = (~E18) | (~S18[6]) | I18;
assign sel19 = (~E19) | (~S19[6]) | I19;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8 & sel9 & sel10 &
    sel11 & sel12 & sel13 & sel14 & sel15 & sel16 & sel17 & sel18 & sel19;
endmodule   // FanoutHash_1EBD0270673B29D7


module FanoutHash_1B10C32F008C11AC (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[17]) | I3;
assign sel4 = (~E4) | (~S4[17]) | I4;
assign sel5 = (~E5) | (~S5[17]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_1B10C32F008C11AC


module FanoutHash_1A568579D8E9714B (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[7]) | I3;
assign sel4 = (~E4) | (~S4[7]) | I4;
assign sel5 = (~E5) | (~S5[7]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_1A568579D8E9714B


module FanoutHash_184DFC10DAF19BE9 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[16]) | I3;
assign sel4 = (~E4) | (~S4[16]) | I4;
assign sel5 = (~E5) | (~S5[16]) | I5;
assign sel6 = (~E6) | (~S6[16]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_184DFC10DAF19BE9


module FanoutHash_1816466D6957000 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[2]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[19]) | I3;
assign sel4 = (~E4) | (~S4[19]) | I4;
assign sel5 = (~E5) | (~S5[19]) | I5;
assign sel6 = (~E6) | (~S6[19]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_1816466D6957000


module FanoutHash_14EBE1E8E49CA541 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic [31:0] S0,
  input logic [31:0] S1,
  input logic [31:0] S2,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
assign sel0 = (~E0) | (~S0[20]) | I0;
assign sel1 = (~E1) | (~S1[20]) | I1;
assign sel2 = (~E2) | (~S2[20]) | I2;
assign O = sel0 & sel1 & sel2;
endmodule   // FanoutHash_14EBE1E8E49CA541


module FanoutHash_13B77C2790BDE4E2 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[1]) | I2;
assign sel3 = (~E3) | (~S3[13]) | I3;
assign sel4 = (~E4) | (~S4[13]) | I4;
assign sel5 = (~E5) | (~S5[13]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_13B77C2790BDE4E2


module FanoutHash_11B554A18790BBBC (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[18]) | I3;
assign sel4 = (~E4) | (~S4[18]) | I4;
assign sel5 = (~E5) | (~S5[18]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_11B554A18790BBBC


module FanoutHash_1130FCC7DFE98006 (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[2]) | I1;
assign sel2 = (~E2) | (~S2[0]) | I2;
assign sel3 = (~E3) | (~S3[6]) | I3;
assign sel4 = (~E4) | (~S4[6]) | I4;
assign sel5 = (~E5) | (~S5[6]) | I5;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5;
endmodule   // FanoutHash_1130FCC7DFE98006


module ExclusiveNodeFanout_H2 (
  input logic [1:0] I,
  input logic [1:0] S,
  output logic O
);

assign O = (I[0] & S[0]) | (I[1] & S[1]);
endmodule   // ExclusiveNodeFanout_H2


module Decode98 (
    input [7:0] I,
    output O
);
wire [7:0] const_9_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h09),
    .width(8)
) const_9_8 (
    .out(const_9_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_9_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode88 (
    input [7:0] I,
    output O
);
wire [7:0] const_8_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h08),
    .width(8)
) const_8_8 (
    .out(const_8_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_8_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode78 (
    input [7:0] I,
    output O
);
wire [7:0] const_7_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h07),
    .width(8)
) const_7_8 (
    .out(const_7_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_7_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode68 (
    input [7:0] I,
    output O
);
wire [7:0] const_6_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h06),
    .width(8)
) const_6_8 (
    .out(const_6_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_6_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode58 (
    input [7:0] I,
    output O
);
wire [7:0] const_5_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h05),
    .width(8)
) const_5_8 (
    .out(const_5_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_5_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode48 (
    input [7:0] I,
    output O
);
wire [7:0] const_4_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h04),
    .width(8)
) const_4_8 (
    .out(const_4_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_4_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode38 (
    input [7:0] I,
    output O
);
wire [7:0] const_3_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h03),
    .width(8)
) const_3_8 (
    .out(const_3_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_3_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode28 (
    input [7:0] I,
    output O
);
wire [7:0] const_2_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h02),
    .width(8)
) const_2_8 (
    .out(const_2_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_2_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode18 (
    input [7:0] I,
    output O
);
wire [7:0] const_1_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h01),
    .width(8)
) const_1_8 (
    .out(const_1_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_1_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode158 (
    input [7:0] I,
    output O
);
wire [7:0] const_15_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0f),
    .width(8)
) const_15_8 (
    .out(const_15_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_15_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode148 (
    input [7:0] I,
    output O
);
wire [7:0] const_14_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0e),
    .width(8)
) const_14_8 (
    .out(const_14_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_14_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode138 (
    input [7:0] I,
    output O
);
wire [7:0] const_13_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0d),
    .width(8)
) const_13_8 (
    .out(const_13_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_13_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode128 (
    input [7:0] I,
    output O
);
wire [7:0] const_12_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0c),
    .width(8)
) const_12_8 (
    .out(const_12_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_12_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode118 (
    input [7:0] I,
    output O
);
wire [7:0] const_11_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0b),
    .width(8)
) const_11_8 (
    .out(const_11_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_11_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode108 (
    input [7:0] I,
    output O
);
wire [7:0] const_10_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0a),
    .width(8)
) const_10_8 (
    .out(const_10_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_10_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode08 (
    input [7:0] I,
    output O
);
wire [7:0] const_0_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_0_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module ConfigRegister_6_8_32_0 (
    input clk,
    input reset,
    output [5:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [5:0] Register_inst0_O;
wire [7:0] const_0_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq2 Register_inst0 (
    .I(config_data[5:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_0_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_9 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_9_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h09),
    .width(8)
) const_9_8 (
    .out(const_9_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_9_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_8 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_8_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h08),
    .width(8)
) const_8_8 (
    .out(const_8_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_8_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_7 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_7_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h07),
    .width(8)
) const_7_8 (
    .out(const_7_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_7_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_6 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_6_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h06),
    .width(8)
) const_6_8 (
    .out(const_6_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_6_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_5 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_5_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h05),
    .width(8)
) const_5_8 (
    .out(const_5_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_5_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_45 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_45_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h2d),
    .width(8)
) const_45_8 (
    .out(const_45_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_45_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_44 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_44_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h2c),
    .width(8)
) const_44_8 (
    .out(const_44_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_44_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_43 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_43_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h2b),
    .width(8)
) const_43_8 (
    .out(const_43_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_43_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_42 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_42_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h2a),
    .width(8)
) const_42_8 (
    .out(const_42_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_42_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_41 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_41_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h29),
    .width(8)
) const_41_8 (
    .out(const_41_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_41_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_4 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_4_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h04),
    .width(8)
) const_4_8 (
    .out(const_4_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_4_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_39 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_39_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h27),
    .width(8)
) const_39_8 (
    .out(const_39_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_39_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_38 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_38_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h26),
    .width(8)
) const_38_8 (
    .out(const_38_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_38_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_37 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_37_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h25),
    .width(8)
) const_37_8 (
    .out(const_37_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_37_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_36 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_36_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h24),
    .width(8)
) const_36_8 (
    .out(const_36_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_36_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_35 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_35_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h23),
    .width(8)
) const_35_8 (
    .out(const_35_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_35_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_34 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_34_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h22),
    .width(8)
) const_34_8 (
    .out(const_34_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_34_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_33 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_33_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h21),
    .width(8)
) const_33_8 (
    .out(const_33_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_33_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_32 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_32_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h20),
    .width(8)
) const_32_8 (
    .out(const_32_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_32_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_31 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_31_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h1f),
    .width(8)
) const_31_8 (
    .out(const_31_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_31_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_30 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_30_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h1e),
    .width(8)
) const_30_8 (
    .out(const_30_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_30_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_3 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_3_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h03),
    .width(8)
) const_3_8 (
    .out(const_3_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_3_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_29 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_29_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h1d),
    .width(8)
) const_29_8 (
    .out(const_29_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_29_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_28 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_28_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h1c),
    .width(8)
) const_28_8 (
    .out(const_28_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_28_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_27 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_27_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h1b),
    .width(8)
) const_27_8 (
    .out(const_27_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_27_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_26 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_26_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h1a),
    .width(8)
) const_26_8 (
    .out(const_26_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_26_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_25 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_25_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h19),
    .width(8)
) const_25_8 (
    .out(const_25_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_25_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_24 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_24_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h18),
    .width(8)
) const_24_8 (
    .out(const_24_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_24_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_23 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_23_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h17),
    .width(8)
) const_23_8 (
    .out(const_23_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_23_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_22 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_22_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h16),
    .width(8)
) const_22_8 (
    .out(const_22_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_22_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_21 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_21_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h15),
    .width(8)
) const_21_8 (
    .out(const_21_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_21_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_20 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_20_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h14),
    .width(8)
) const_20_8 (
    .out(const_20_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_20_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_2 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_2_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h02),
    .width(8)
) const_2_8 (
    .out(const_2_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_2_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_19 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_19_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h13),
    .width(8)
) const_19_8 (
    .out(const_19_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_19_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_18 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_18_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h12),
    .width(8)
) const_18_8 (
    .out(const_18_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_18_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_17 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_17_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h11),
    .width(8)
) const_17_8 (
    .out(const_17_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_17_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_16 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_16_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h10),
    .width(8)
) const_16_8 (
    .out(const_16_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_16_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_15 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_15_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0f),
    .width(8)
) const_15_8 (
    .out(const_15_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_15_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_14 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_14_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0e),
    .width(8)
) const_14_8 (
    .out(const_14_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_14_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_13 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_13_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0d),
    .width(8)
) const_13_8 (
    .out(const_13_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_13_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_12 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_12_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0c),
    .width(8)
) const_12_8 (
    .out(const_12_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_12_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_11 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_11_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0b),
    .width(8)
) const_11_8 (
    .out(const_11_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_11_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_10 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_10_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0a),
    .width(8)
) const_10_8 (
    .out(const_10_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_10_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_1 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_1_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h01),
    .width(8)
) const_1_8 (
    .out(const_1_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_1_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_32_8_32_0 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_inst0_O;
wire [7:0] const_0_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register Register_inst0 (
    .I(config_data),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_0_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_31_8_32_3 (
    input clk,
    input reset,
    output [30:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [30:0] Register_inst0_O;
wire [7:0] const_3_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq5 Register_inst0 (
    .I(config_data[30:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h03),
    .width(8)
) const_3_8 (
    .out(const_3_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_3_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_30_8_32_8 (
    input clk,
    input reset,
    output [29:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [29:0] Register_inst0_O;
wire [7:0] const_8_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq3 Register_inst0 (
    .I(config_data[29:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h08),
    .width(8)
) const_8_8 (
    .out(const_8_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_8_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_30_8_32_4 (
    input clk,
    input reset,
    output [29:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [29:0] Register_inst0_O;
wire [7:0] const_4_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq3 Register_inst0 (
    .I(config_data[29:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h04),
    .width(8)
) const_4_8 (
    .out(const_4_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_4_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_25_8_32_46 (
    input clk,
    input reset,
    output [24:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [24:0] Register_inst0_O;
wire [7:0] const_46_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq8 Register_inst0 (
    .I(config_data[24:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h2e),
    .width(8)
) const_46_8 (
    .out(const_46_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_46_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module ConfigRegister_24_8_32_0 (
    input clk,
    input reset,
    output [23:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [23:0] Register_inst0_O;
wire [7:0] const_0_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq9 Register_inst0 (
    .I(config_data[23:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_0_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module IOCoreReadyValid (
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    input [0:0] f2io_1,
    input [16:0] f2io_17,
    output [0:0] f2io_17_ready,
    input [0:0] f2io_17_valid,
    output [0:0] f2io_1_ready,
    input [0:0] f2io_1_valid,
    input [0:0] flush,
    input [0:0] flush_core,
    input [0:0] glb2io_1,
    input [16:0] glb2io_17,
    output [0:0] glb2io_17_ready,
    input [0:0] glb2io_17_valid,
    output [0:0] glb2io_1_ready,
    input [0:0] glb2io_1_valid,
    output [0:0] io2f_1,
    output [16:0] io2f_17,
    input [0:0] io2f_17_ready,
    output [0:0] io2f_17_valid,
    input [0:0] io2f_1_ready,
    output [0:0] io2f_1_valid,
    output [0:0] io2glb_1,
    output [16:0] io2glb_17,
    input [0:0] io2glb_17_ready,
    output [0:0] io2glb_17_valid,
    input [0:0] io2glb_1_ready,
    output [0:0] io2glb_1_valid,
    output [31:0] read_config_data,
    input reset,
    input [0:0] stall
);
wire [0:0] Invert1_inst0_out;
wire [0:0] Invert1_inst1_out;
wire ZextWrapper_24_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_24_32_inst0$self_O_in;
wire [23:0] config_reg_0_O;
wire coreir_wrapInAsyncReset_inst0_out;
wire coreir_wrapOutAsyncReset_inst0_out;
wire [0:0] f2io_17_valid_reg_sel_value_O;
wire [0:0] f2io_17_valid_reg_value_value_O;
wire [0:0] f2io_17_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] f2io_1_reg_sel_value_O;
wire [0:0] f2io_1_reg_value_value_O;
wire [0:0] f2io_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] f2io_1_valid_reg_sel_value_O;
wire [0:0] f2io_1_valid_reg_value_value_O;
wire [0:0] f2io_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] flush_mux_sel_value_O;
wire [0:0] flush_reg_sel_value_O;
wire [0:0] flush_reg_value_value_O;
wire [0:0] flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] glb2io_17_valid_reg_sel_value_O;
wire [0:0] glb2io_17_valid_reg_value_value_O;
wire [0:0] glb2io_17_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] glb2io_1_reg_sel_value_O;
wire [0:0] glb2io_1_reg_value_value_O;
wire [0:0] glb2io_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] glb2io_1_valid_reg_sel_value_O;
wire [0:0] glb2io_1_valid_reg_value_value_O;
wire [0:0] glb2io_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] io2f_17_ready_reg_sel_value_O;
wire [0:0] io2f_17_ready_reg_value_value_O;
wire [0:0] io2f_17_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] io2f_1_ready_reg_sel_value_O;
wire [0:0] io2f_1_ready_reg_value_value_O;
wire [0:0] io2f_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] io2glb_17_ready_reg_sel_value_O;
wire [0:0] io2glb_17_ready_reg_value_value_O;
wire [0:0] io2glb_17_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] io2glb_1_ready_reg_sel_value_O;
wire [0:0] io2glb_1_ready_reg_value_value_O;
wire [0:0] io2glb_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [16:0] io_core_W_inst0_io2glb_17;
wire [0:0] io_core_W_inst0_io2glb_17_valid;
wire [0:0] io_core_W_inst0_f2io_1_ready;
wire [0:0] io_core_W_inst0_glb2io_17_ready;
wire [16:0] io_core_W_inst0_io2f_17;
wire [0:0] io_core_W_inst0_io2glb_1;
wire [0:0] io_core_W_inst0_io2f_1_valid;
wire [0:0] io_core_W_inst0_io2glb_1_valid;
wire [0:0] io_core_W_inst0_glb2io_1_ready;
wire [0:0] io_core_W_inst0_f2io_17_ready;
wire [0:0] io_core_W_inst0_io2f_17_valid;
wire [0:0] io_core_W_inst0_io2f_1;
wire [0:0] tile_en_value_O;
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(coreir_wrapInAsyncReset_inst0_out),
    .out(Invert1_inst0_out)
);
coreir_not #(
    .width(1)
) Invert1_inst1 (
    .in(stall),
    .out(Invert1_inst1_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_24_32_inst0$bit_const_0_None (
    .out(ZextWrapper_24_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_24_32_inst0$self_O_out;
assign ZextWrapper_24_32_inst0$self_O_out = {ZextWrapper_24_32_inst0$bit_const_0_None_out,ZextWrapper_24_32_inst0$bit_const_0_None_out,ZextWrapper_24_32_inst0$bit_const_0_None_out,ZextWrapper_24_32_inst0$bit_const_0_None_out,ZextWrapper_24_32_inst0$bit_const_0_None_out,ZextWrapper_24_32_inst0$bit_const_0_None_out,ZextWrapper_24_32_inst0$bit_const_0_None_out,ZextWrapper_24_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_24_32_inst0$self_O (
    .in(ZextWrapper_24_32_inst0$self_O_in),
    .out(ZextWrapper_24_32_inst0$self_O_out)
);
ConfigRegister_24_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_wrap coreir_wrapInAsyncReset_inst0 (
    .in(reset),
    .out(coreir_wrapInAsyncReset_inst0_out)
);
coreir_wrap coreir_wrapOutAsyncReset_inst0 (
    .in(Invert1_inst0_out[0]),
    .out(coreir_wrapOutAsyncReset_inst0_out)
);
SliceWrapper_24_0_1 f2io_17_valid_reg_sel_value (
    .I(config_reg_0_O),
    .O(f2io_17_valid_reg_sel_value_O)
);
SliceWrapper_24_1_2 f2io_17_valid_reg_value_value (
    .I(config_reg_0_O),
    .O(f2io_17_valid_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) f2io_17_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(f2io_17_valid),
    .in1(f2io_17_valid_reg_value_value_O),
    .sel(f2io_17_valid_reg_sel_value_O[0]),
    .out(f2io_17_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_24_2_3 f2io_1_reg_sel_value (
    .I(config_reg_0_O),
    .O(f2io_1_reg_sel_value_O)
);
SliceWrapper_24_3_4 f2io_1_reg_value_value (
    .I(config_reg_0_O),
    .O(f2io_1_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) f2io_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(f2io_1),
    .in1(f2io_1_reg_value_value_O),
    .sel(f2io_1_reg_sel_value_O[0]),
    .out(f2io_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_24_4_5 f2io_1_valid_reg_sel_value (
    .I(config_reg_0_O),
    .O(f2io_1_valid_reg_sel_value_O)
);
SliceWrapper_24_5_6 f2io_1_valid_reg_value_value (
    .I(config_reg_0_O),
    .O(f2io_1_valid_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) f2io_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(f2io_1_valid),
    .in1(f2io_1_valid_reg_value_value_O),
    .sel(f2io_1_valid_reg_sel_value_O[0]),
    .out(f2io_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(flush_core),
    .in1(flush),
    .sel(flush_mux_sel_value_O[0]),
    .out(flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_24_6_7 flush_mux_sel_value (
    .I(config_reg_0_O),
    .O(flush_mux_sel_value_O)
);
SliceWrapper_24_7_8 flush_reg_sel_value (
    .I(config_reg_0_O),
    .O(flush_reg_sel_value_O)
);
SliceWrapper_24_8_9 flush_reg_value_value (
    .I(config_reg_0_O),
    .O(flush_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(flush),
    .in1(flush_reg_value_value_O),
    .sel(flush_reg_sel_value_O[0]),
    .out(flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_24_9_10 glb2io_17_valid_reg_sel_value (
    .I(config_reg_0_O),
    .O(glb2io_17_valid_reg_sel_value_O)
);
SliceWrapper_24_10_11 glb2io_17_valid_reg_value_value (
    .I(config_reg_0_O),
    .O(glb2io_17_valid_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) glb2io_17_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(glb2io_17_valid),
    .in1(glb2io_17_valid_reg_value_value_O),
    .sel(glb2io_17_valid_reg_sel_value_O[0]),
    .out(glb2io_17_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_24_11_12 glb2io_1_reg_sel_value (
    .I(config_reg_0_O),
    .O(glb2io_1_reg_sel_value_O)
);
SliceWrapper_24_12_13 glb2io_1_reg_value_value (
    .I(config_reg_0_O),
    .O(glb2io_1_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) glb2io_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(glb2io_1),
    .in1(glb2io_1_reg_value_value_O),
    .sel(glb2io_1_reg_sel_value_O[0]),
    .out(glb2io_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_24_13_14 glb2io_1_valid_reg_sel_value (
    .I(config_reg_0_O),
    .O(glb2io_1_valid_reg_sel_value_O)
);
SliceWrapper_24_14_15 glb2io_1_valid_reg_value_value (
    .I(config_reg_0_O),
    .O(glb2io_1_valid_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) glb2io_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(glb2io_1_valid),
    .in1(glb2io_1_valid_reg_value_value_O),
    .sel(glb2io_1_valid_reg_sel_value_O[0]),
    .out(glb2io_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_24_15_16 io2f_17_ready_reg_sel_value (
    .I(config_reg_0_O),
    .O(io2f_17_ready_reg_sel_value_O)
);
SliceWrapper_24_16_17 io2f_17_ready_reg_value_value (
    .I(config_reg_0_O),
    .O(io2f_17_ready_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) io2f_17_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(io2f_17_ready),
    .in1(io2f_17_ready_reg_value_value_O),
    .sel(io2f_17_ready_reg_sel_value_O[0]),
    .out(io2f_17_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_24_17_18 io2f_1_ready_reg_sel_value (
    .I(config_reg_0_O),
    .O(io2f_1_ready_reg_sel_value_O)
);
SliceWrapper_24_18_19 io2f_1_ready_reg_value_value (
    .I(config_reg_0_O),
    .O(io2f_1_ready_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) io2f_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(io2f_1_ready),
    .in1(io2f_1_ready_reg_value_value_O),
    .sel(io2f_1_ready_reg_sel_value_O[0]),
    .out(io2f_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_24_19_20 io2glb_17_ready_reg_sel_value (
    .I(config_reg_0_O),
    .O(io2glb_17_ready_reg_sel_value_O)
);
SliceWrapper_24_20_21 io2glb_17_ready_reg_value_value (
    .I(config_reg_0_O),
    .O(io2glb_17_ready_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) io2glb_17_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(io2glb_17_ready),
    .in1(io2glb_17_ready_reg_value_value_O),
    .sel(io2glb_17_ready_reg_sel_value_O[0]),
    .out(io2glb_17_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_24_21_22 io2glb_1_ready_reg_sel_value (
    .I(config_reg_0_O),
    .O(io2glb_1_ready_reg_sel_value_O)
);
SliceWrapper_24_22_23 io2glb_1_ready_reg_value_value (
    .I(config_reg_0_O),
    .O(io2glb_1_ready_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) io2glb_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(io2glb_1_ready),
    .in1(io2glb_1_ready_reg_value_value_O),
    .sel(io2glb_1_ready_reg_sel_value_O[0]),
    .out(io2glb_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
io_core_W io_core_W_inst0 (
    .io2glb_17(io_core_W_inst0_io2glb_17),
    .io2glb_17_valid(io_core_W_inst0_io2glb_17_valid),
    .f2io_17(f2io_17),
    .glb2io_1_valid(glb2io_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .f2io_1_ready(io_core_W_inst0_f2io_1_ready),
    .rst_n(coreir_wrapOutAsyncReset_inst0_out),
    .glb2io_17_valid(glb2io_17_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .tile_en(tile_en_value_O),
    .clk(clk),
    .glb2io_17_ready(io_core_W_inst0_glb2io_17_ready),
    .io2f_1_ready(io2f_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .io2glb_17_ready(io2glb_17_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .io2f_17(io_core_W_inst0_io2f_17),
    .io2glb_1(io_core_W_inst0_io2glb_1),
    .io2f_1_valid(io_core_W_inst0_io2f_1_valid),
    .f2io_17_valid(f2io_17_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .io2glb_1_valid(io_core_W_inst0_io2glb_1_valid),
    .glb2io_1_ready(io_core_W_inst0_glb2io_1_ready),
    .io2f_17_ready(io2f_17_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .io2glb_1_ready(io2glb_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .clk_en(Invert1_inst1_out),
    .f2io_17_ready(io_core_W_inst0_f2io_17_ready),
    .glb2io_1(glb2io_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .io2f_17_valid(io_core_W_inst0_io2f_17_valid),
    .f2io_1(f2io_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .io2f_1(io_core_W_inst0_io2f_1),
    .flush(flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .glb2io_17(glb2io_17),
    .f2io_1_valid(f2io_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_24_23_24 tile_en_value (
    .I(config_reg_0_O),
    .O(tile_en_value_O)
);
assign f2io_17_ready = io_core_W_inst0_f2io_17_ready;
assign f2io_1_ready = io_core_W_inst0_f2io_1_ready;
assign glb2io_17_ready = io_core_W_inst0_glb2io_17_ready;
assign glb2io_1_ready = io_core_W_inst0_glb2io_1_ready;
assign io2f_1 = io_core_W_inst0_io2f_1;
assign io2f_17 = io_core_W_inst0_io2f_17;
assign io2f_17_valid = io_core_W_inst0_io2f_17_valid;
assign io2f_1_valid = io_core_W_inst0_io2f_1_valid;
assign io2glb_1 = io_core_W_inst0_io2glb_1;
assign io2glb_17 = io_core_W_inst0_io2glb_17;
assign io2glb_17_valid = io_core_W_inst0_io2glb_17_valid;
assign io2glb_1_valid = io_core_W_inst0_io2glb_1_valid;
assign read_config_data = ZextWrapper_24_32_inst0$self_O_in;
endmodule

module ConfigRegister_23_8_32_5 (
    input clk,
    input reset,
    output [22:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [22:0] Register_inst0_O;
wire [7:0] const_5_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq6 Register_inst0 (
    .I(config_data[22:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h05),
    .width(8)
) const_5_8 (
    .out(const_5_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_5_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module SB_ID0_5TRACKS_B1_PE (
    input [0:0] PE_input_width_1_num_0_enable,
    input [31:0] PE_input_width_1_num_0_out_sel,
    input PE_input_width_1_num_0_ready,
    input [0:0] PE_input_width_1_num_1_enable,
    input [31:0] PE_input_width_1_num_1_out_sel,
    input PE_input_width_1_num_1_ready,
    input [0:0] PE_input_width_1_num_2_enable,
    input [31:0] PE_input_width_1_num_2_out_sel,
    input PE_input_width_1_num_2_ready,
    input [0:0] PE_output_width_1_num_0,
    output PE_output_width_1_num_0_ready_out,
    input PE_output_width_1_num_0_valid,
    input [0:0] PondTop_output_width_1_num_0,
    output PondTop_output_width_1_num_0_ready_out,
    input PondTop_output_width_1_num_0_valid,
    input [0:0] PondTop_output_width_1_num_1,
    output PondTop_output_width_1_num_1_ready_out,
    input PondTop_output_width_1_num_1_valid,
    input [0:0] SB_T0_EAST_SB_IN_B1,
    output SB_T0_EAST_SB_IN_B1_enable,
    output SB_T0_EAST_SB_IN_B1_ready_out,
    input SB_T0_EAST_SB_IN_B1_valid_in,
    output [0:0] SB_T0_EAST_SB_OUT_B1,
    output SB_T0_EAST_SB_OUT_B1_enable,
    input SB_T0_EAST_SB_OUT_B1_ready_in,
    output SB_T0_EAST_SB_OUT_B1_valid_out,
    input [0:0] SB_T0_NORTH_SB_IN_B1,
    output SB_T0_NORTH_SB_IN_B1_enable,
    output SB_T0_NORTH_SB_IN_B1_ready_out,
    input SB_T0_NORTH_SB_IN_B1_valid_in,
    output [0:0] SB_T0_NORTH_SB_OUT_B1,
    output SB_T0_NORTH_SB_OUT_B1_enable,
    input SB_T0_NORTH_SB_OUT_B1_ready_in,
    output SB_T0_NORTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T0_SOUTH_SB_IN_B1,
    output SB_T0_SOUTH_SB_IN_B1_enable,
    output SB_T0_SOUTH_SB_IN_B1_ready_out,
    input SB_T0_SOUTH_SB_IN_B1_valid_in,
    output [0:0] SB_T0_SOUTH_SB_OUT_B1,
    output SB_T0_SOUTH_SB_OUT_B1_enable,
    input SB_T0_SOUTH_SB_OUT_B1_ready_in,
    output SB_T0_SOUTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T0_WEST_SB_IN_B1,
    output SB_T0_WEST_SB_IN_B1_enable,
    output SB_T0_WEST_SB_IN_B1_ready_out,
    input SB_T0_WEST_SB_IN_B1_valid_in,
    output [0:0] SB_T0_WEST_SB_OUT_B1,
    output SB_T0_WEST_SB_OUT_B1_enable,
    input SB_T0_WEST_SB_OUT_B1_ready_in,
    output SB_T0_WEST_SB_OUT_B1_valid_out,
    input [0:0] SB_T1_EAST_SB_IN_B1,
    output SB_T1_EAST_SB_IN_B1_enable,
    output SB_T1_EAST_SB_IN_B1_ready_out,
    input SB_T1_EAST_SB_IN_B1_valid_in,
    output [0:0] SB_T1_EAST_SB_OUT_B1,
    output SB_T1_EAST_SB_OUT_B1_enable,
    input SB_T1_EAST_SB_OUT_B1_ready_in,
    output SB_T1_EAST_SB_OUT_B1_valid_out,
    input [0:0] SB_T1_NORTH_SB_IN_B1,
    output SB_T1_NORTH_SB_IN_B1_enable,
    output SB_T1_NORTH_SB_IN_B1_ready_out,
    input SB_T1_NORTH_SB_IN_B1_valid_in,
    output [0:0] SB_T1_NORTH_SB_OUT_B1,
    output SB_T1_NORTH_SB_OUT_B1_enable,
    input SB_T1_NORTH_SB_OUT_B1_ready_in,
    output SB_T1_NORTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T1_SOUTH_SB_IN_B1,
    output SB_T1_SOUTH_SB_IN_B1_enable,
    output SB_T1_SOUTH_SB_IN_B1_ready_out,
    input SB_T1_SOUTH_SB_IN_B1_valid_in,
    output [0:0] SB_T1_SOUTH_SB_OUT_B1,
    output SB_T1_SOUTH_SB_OUT_B1_enable,
    input SB_T1_SOUTH_SB_OUT_B1_ready_in,
    output SB_T1_SOUTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T1_WEST_SB_IN_B1,
    output SB_T1_WEST_SB_IN_B1_enable,
    output SB_T1_WEST_SB_IN_B1_ready_out,
    input SB_T1_WEST_SB_IN_B1_valid_in,
    output [0:0] SB_T1_WEST_SB_OUT_B1,
    output SB_T1_WEST_SB_OUT_B1_enable,
    input SB_T1_WEST_SB_OUT_B1_ready_in,
    output SB_T1_WEST_SB_OUT_B1_valid_out,
    input [0:0] SB_T2_EAST_SB_IN_B1,
    output SB_T2_EAST_SB_IN_B1_enable,
    output SB_T2_EAST_SB_IN_B1_ready_out,
    input SB_T2_EAST_SB_IN_B1_valid_in,
    output [0:0] SB_T2_EAST_SB_OUT_B1,
    output SB_T2_EAST_SB_OUT_B1_enable,
    input SB_T2_EAST_SB_OUT_B1_ready_in,
    output SB_T2_EAST_SB_OUT_B1_valid_out,
    input [0:0] SB_T2_NORTH_SB_IN_B1,
    output SB_T2_NORTH_SB_IN_B1_enable,
    output SB_T2_NORTH_SB_IN_B1_ready_out,
    input SB_T2_NORTH_SB_IN_B1_valid_in,
    output [0:0] SB_T2_NORTH_SB_OUT_B1,
    output SB_T2_NORTH_SB_OUT_B1_enable,
    input SB_T2_NORTH_SB_OUT_B1_ready_in,
    output SB_T2_NORTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T2_SOUTH_SB_IN_B1,
    output SB_T2_SOUTH_SB_IN_B1_enable,
    output SB_T2_SOUTH_SB_IN_B1_ready_out,
    input SB_T2_SOUTH_SB_IN_B1_valid_in,
    output [0:0] SB_T2_SOUTH_SB_OUT_B1,
    output SB_T2_SOUTH_SB_OUT_B1_enable,
    input SB_T2_SOUTH_SB_OUT_B1_ready_in,
    output SB_T2_SOUTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T2_WEST_SB_IN_B1,
    output SB_T2_WEST_SB_IN_B1_enable,
    output SB_T2_WEST_SB_IN_B1_ready_out,
    input SB_T2_WEST_SB_IN_B1_valid_in,
    output [0:0] SB_T2_WEST_SB_OUT_B1,
    output SB_T2_WEST_SB_OUT_B1_enable,
    input SB_T2_WEST_SB_OUT_B1_ready_in,
    output SB_T2_WEST_SB_OUT_B1_valid_out,
    input [0:0] SB_T3_EAST_SB_IN_B1,
    output SB_T3_EAST_SB_IN_B1_enable,
    output SB_T3_EAST_SB_IN_B1_ready_out,
    input SB_T3_EAST_SB_IN_B1_valid_in,
    output [0:0] SB_T3_EAST_SB_OUT_B1,
    output SB_T3_EAST_SB_OUT_B1_enable,
    input SB_T3_EAST_SB_OUT_B1_ready_in,
    output SB_T3_EAST_SB_OUT_B1_valid_out,
    input [0:0] SB_T3_NORTH_SB_IN_B1,
    output SB_T3_NORTH_SB_IN_B1_enable,
    output SB_T3_NORTH_SB_IN_B1_ready_out,
    input SB_T3_NORTH_SB_IN_B1_valid_in,
    output [0:0] SB_T3_NORTH_SB_OUT_B1,
    output SB_T3_NORTH_SB_OUT_B1_enable,
    input SB_T3_NORTH_SB_OUT_B1_ready_in,
    output SB_T3_NORTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T3_SOUTH_SB_IN_B1,
    output SB_T3_SOUTH_SB_IN_B1_enable,
    output SB_T3_SOUTH_SB_IN_B1_ready_out,
    input SB_T3_SOUTH_SB_IN_B1_valid_in,
    output [0:0] SB_T3_SOUTH_SB_OUT_B1,
    output SB_T3_SOUTH_SB_OUT_B1_enable,
    input SB_T3_SOUTH_SB_OUT_B1_ready_in,
    output SB_T3_SOUTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T3_WEST_SB_IN_B1,
    output SB_T3_WEST_SB_IN_B1_enable,
    output SB_T3_WEST_SB_IN_B1_ready_out,
    input SB_T3_WEST_SB_IN_B1_valid_in,
    output [0:0] SB_T3_WEST_SB_OUT_B1,
    output SB_T3_WEST_SB_OUT_B1_enable,
    input SB_T3_WEST_SB_OUT_B1_ready_in,
    output SB_T3_WEST_SB_OUT_B1_valid_out,
    input [0:0] SB_T4_EAST_SB_IN_B1,
    output SB_T4_EAST_SB_IN_B1_enable,
    output SB_T4_EAST_SB_IN_B1_ready_out,
    input SB_T4_EAST_SB_IN_B1_valid_in,
    output [0:0] SB_T4_EAST_SB_OUT_B1,
    output SB_T4_EAST_SB_OUT_B1_enable,
    input SB_T4_EAST_SB_OUT_B1_ready_in,
    output SB_T4_EAST_SB_OUT_B1_valid_out,
    input [0:0] SB_T4_NORTH_SB_IN_B1,
    output SB_T4_NORTH_SB_IN_B1_enable,
    output SB_T4_NORTH_SB_IN_B1_ready_out,
    input SB_T4_NORTH_SB_IN_B1_valid_in,
    output [0:0] SB_T4_NORTH_SB_OUT_B1,
    output SB_T4_NORTH_SB_OUT_B1_enable,
    input SB_T4_NORTH_SB_OUT_B1_ready_in,
    output SB_T4_NORTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T4_SOUTH_SB_IN_B1,
    output SB_T4_SOUTH_SB_IN_B1_enable,
    output SB_T4_SOUTH_SB_IN_B1_ready_out,
    input SB_T4_SOUTH_SB_IN_B1_valid_in,
    output [0:0] SB_T4_SOUTH_SB_OUT_B1,
    output SB_T4_SOUTH_SB_OUT_B1_enable,
    input SB_T4_SOUTH_SB_OUT_B1_ready_in,
    output SB_T4_SOUTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T4_WEST_SB_IN_B1,
    output SB_T4_WEST_SB_IN_B1_enable,
    output SB_T4_WEST_SB_IN_B1_ready_out,
    input SB_T4_WEST_SB_IN_B1_valid_in,
    output [0:0] SB_T4_WEST_SB_OUT_B1,
    output SB_T4_WEST_SB_OUT_B1_enable,
    input SB_T4_WEST_SB_OUT_B1_ready_in,
    output SB_T4_WEST_SB_OUT_B1_valid_out,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset,
    input [0:0] stall
);
wire [0:0] CB_PE_output_width_1_num_0_fan_in_O;
wire [0:0] CB_PondTop_output_width_1_num_0_fan_in_O;
wire [0:0] CB_PondTop_output_width_1_num_1_fan_in_O;
wire [0:0] Invert1_inst0_out;
wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1_O;
wire MUX_SB_T0_EAST_SB_OUT_B1_ready_out;
wire MUX_SB_T0_EAST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T0_EAST_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1_O;
wire MUX_SB_T0_NORTH_SB_OUT_B1_ready_out;
wire MUX_SB_T0_NORTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T0_NORTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1_O;
wire MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out;
wire MUX_SB_T0_SOUTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1_O;
wire MUX_SB_T0_WEST_SB_OUT_B1_ready_out;
wire MUX_SB_T0_WEST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T0_WEST_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1_O;
wire MUX_SB_T1_EAST_SB_OUT_B1_ready_out;
wire MUX_SB_T1_EAST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T1_EAST_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1_O;
wire MUX_SB_T1_NORTH_SB_OUT_B1_ready_out;
wire MUX_SB_T1_NORTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T1_NORTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1_O;
wire MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out;
wire MUX_SB_T1_SOUTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1_O;
wire MUX_SB_T1_WEST_SB_OUT_B1_ready_out;
wire MUX_SB_T1_WEST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T1_WEST_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1_O;
wire MUX_SB_T2_EAST_SB_OUT_B1_ready_out;
wire MUX_SB_T2_EAST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T2_EAST_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1_O;
wire MUX_SB_T2_NORTH_SB_OUT_B1_ready_out;
wire MUX_SB_T2_NORTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T2_NORTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1_O;
wire MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out;
wire MUX_SB_T2_SOUTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1_O;
wire MUX_SB_T2_WEST_SB_OUT_B1_ready_out;
wire MUX_SB_T2_WEST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T2_WEST_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1_O;
wire MUX_SB_T3_EAST_SB_OUT_B1_ready_out;
wire MUX_SB_T3_EAST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T3_EAST_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1_O;
wire MUX_SB_T3_NORTH_SB_OUT_B1_ready_out;
wire MUX_SB_T3_NORTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T3_NORTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1_O;
wire MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out;
wire MUX_SB_T3_SOUTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1_O;
wire MUX_SB_T3_WEST_SB_OUT_B1_ready_out;
wire MUX_SB_T3_WEST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T3_WEST_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1_O;
wire MUX_SB_T4_EAST_SB_OUT_B1_ready_out;
wire MUX_SB_T4_EAST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T4_EAST_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1_O;
wire MUX_SB_T4_NORTH_SB_OUT_B1_ready_out;
wire MUX_SB_T4_NORTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T4_NORTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1_O;
wire MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out;
wire MUX_SB_T4_SOUTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1_O;
wire MUX_SB_T4_WEST_SB_OUT_B1_ready_out;
wire MUX_SB_T4_WEST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T4_WEST_SB_OUT_B1_out_sel;
wire [0:0] REG_T0_EAST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T0_EAST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T0_EAST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T0_EAST_B1_end_value_O;
wire [0:0] REG_T0_EAST_B1_fifo_value_O;
wire [0:0] REG_T0_EAST_B1_start_value_O;
wire [0:0] REG_T0_NORTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T0_NORTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T0_NORTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T0_NORTH_B1_end_value_O;
wire [0:0] REG_T0_NORTH_B1_fifo_value_O;
wire [0:0] REG_T0_NORTH_B1_start_value_O;
wire [0:0] REG_T0_SOUTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T0_SOUTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T0_SOUTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T0_SOUTH_B1_end_value_O;
wire [0:0] REG_T0_SOUTH_B1_fifo_value_O;
wire [0:0] REG_T0_SOUTH_B1_start_value_O;
wire [0:0] REG_T0_WEST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T0_WEST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T0_WEST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T0_WEST_B1_end_value_O;
wire [0:0] REG_T0_WEST_B1_fifo_value_O;
wire [0:0] REG_T0_WEST_B1_start_value_O;
wire [0:0] REG_T1_EAST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T1_EAST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T1_EAST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T1_EAST_B1_end_value_O;
wire [0:0] REG_T1_EAST_B1_fifo_value_O;
wire [0:0] REG_T1_EAST_B1_start_value_O;
wire [0:0] REG_T1_NORTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T1_NORTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T1_NORTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T1_NORTH_B1_end_value_O;
wire [0:0] REG_T1_NORTH_B1_fifo_value_O;
wire [0:0] REG_T1_NORTH_B1_start_value_O;
wire [0:0] REG_T1_SOUTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T1_SOUTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T1_SOUTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T1_SOUTH_B1_end_value_O;
wire [0:0] REG_T1_SOUTH_B1_fifo_value_O;
wire [0:0] REG_T1_SOUTH_B1_start_value_O;
wire [0:0] REG_T1_WEST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T1_WEST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T1_WEST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T1_WEST_B1_end_value_O;
wire [0:0] REG_T1_WEST_B1_fifo_value_O;
wire [0:0] REG_T1_WEST_B1_start_value_O;
wire [0:0] REG_T2_EAST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T2_EAST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T2_EAST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T2_EAST_B1_end_value_O;
wire [0:0] REG_T2_EAST_B1_fifo_value_O;
wire [0:0] REG_T2_EAST_B1_start_value_O;
wire [0:0] REG_T2_NORTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T2_NORTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T2_NORTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T2_NORTH_B1_end_value_O;
wire [0:0] REG_T2_NORTH_B1_fifo_value_O;
wire [0:0] REG_T2_NORTH_B1_start_value_O;
wire [0:0] REG_T2_SOUTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T2_SOUTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T2_SOUTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T2_SOUTH_B1_end_value_O;
wire [0:0] REG_T2_SOUTH_B1_fifo_value_O;
wire [0:0] REG_T2_SOUTH_B1_start_value_O;
wire [0:0] REG_T2_WEST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T2_WEST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T2_WEST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T2_WEST_B1_end_value_O;
wire [0:0] REG_T2_WEST_B1_fifo_value_O;
wire [0:0] REG_T2_WEST_B1_start_value_O;
wire [0:0] REG_T3_EAST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T3_EAST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T3_EAST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T3_EAST_B1_end_value_O;
wire [0:0] REG_T3_EAST_B1_fifo_value_O;
wire [0:0] REG_T3_EAST_B1_start_value_O;
wire [0:0] REG_T3_NORTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T3_NORTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T3_NORTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T3_NORTH_B1_end_value_O;
wire [0:0] REG_T3_NORTH_B1_fifo_value_O;
wire [0:0] REG_T3_NORTH_B1_start_value_O;
wire [0:0] REG_T3_SOUTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T3_SOUTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T3_SOUTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T3_SOUTH_B1_end_value_O;
wire [0:0] REG_T3_SOUTH_B1_fifo_value_O;
wire [0:0] REG_T3_SOUTH_B1_start_value_O;
wire [0:0] REG_T3_WEST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T3_WEST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T3_WEST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T3_WEST_B1_end_value_O;
wire [0:0] REG_T3_WEST_B1_fifo_value_O;
wire [0:0] REG_T3_WEST_B1_start_value_O;
wire [0:0] REG_T4_EAST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T4_EAST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T4_EAST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T4_EAST_B1_end_value_O;
wire [0:0] REG_T4_EAST_B1_fifo_value_O;
wire [0:0] REG_T4_EAST_B1_start_value_O;
wire [0:0] REG_T4_NORTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T4_NORTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T4_NORTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T4_NORTH_B1_end_value_O;
wire [0:0] REG_T4_NORTH_B1_fifo_value_O;
wire [0:0] REG_T4_NORTH_B1_start_value_O;
wire [0:0] REG_T4_SOUTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T4_SOUTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T4_SOUTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T4_SOUTH_B1_end_value_O;
wire [0:0] REG_T4_SOUTH_B1_fifo_value_O;
wire [0:0] REG_T4_SOUTH_B1_start_value_O;
wire [0:0] REG_T4_WEST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T4_WEST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T4_WEST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T4_WEST_B1_end_value_O;
wire [0:0] REG_T4_WEST_B1_fifo_value_O;
wire [0:0] REG_T4_WEST_B1_start_value_O;
wire [0:0] RMUX_T0_EAST_B1_O;
wire RMUX_T0_EAST_B1_ready_out;
wire RMUX_T0_EAST_B1_valid_out;
wire [1:0] RMUX_T0_EAST_B1_out_sel;
wire [0:0] RMUX_T0_EAST_B1_sel_value_O;
wire [0:0] RMUX_T0_NORTH_B1_O;
wire RMUX_T0_NORTH_B1_ready_out;
wire RMUX_T0_NORTH_B1_valid_out;
wire [1:0] RMUX_T0_NORTH_B1_out_sel;
wire [0:0] RMUX_T0_NORTH_B1_sel_value_O;
wire [0:0] RMUX_T0_SOUTH_B1_O;
wire RMUX_T0_SOUTH_B1_ready_out;
wire RMUX_T0_SOUTH_B1_valid_out;
wire [1:0] RMUX_T0_SOUTH_B1_out_sel;
wire [0:0] RMUX_T0_SOUTH_B1_sel_value_O;
wire [0:0] RMUX_T0_WEST_B1_O;
wire RMUX_T0_WEST_B1_ready_out;
wire RMUX_T0_WEST_B1_valid_out;
wire [1:0] RMUX_T0_WEST_B1_out_sel;
wire [0:0] RMUX_T0_WEST_B1_sel_value_O;
wire [0:0] RMUX_T1_EAST_B1_O;
wire RMUX_T1_EAST_B1_ready_out;
wire RMUX_T1_EAST_B1_valid_out;
wire [1:0] RMUX_T1_EAST_B1_out_sel;
wire [0:0] RMUX_T1_EAST_B1_sel_value_O;
wire [0:0] RMUX_T1_NORTH_B1_O;
wire RMUX_T1_NORTH_B1_ready_out;
wire RMUX_T1_NORTH_B1_valid_out;
wire [1:0] RMUX_T1_NORTH_B1_out_sel;
wire [0:0] RMUX_T1_NORTH_B1_sel_value_O;
wire [0:0] RMUX_T1_SOUTH_B1_O;
wire RMUX_T1_SOUTH_B1_ready_out;
wire RMUX_T1_SOUTH_B1_valid_out;
wire [1:0] RMUX_T1_SOUTH_B1_out_sel;
wire [0:0] RMUX_T1_SOUTH_B1_sel_value_O;
wire [0:0] RMUX_T1_WEST_B1_O;
wire RMUX_T1_WEST_B1_ready_out;
wire RMUX_T1_WEST_B1_valid_out;
wire [1:0] RMUX_T1_WEST_B1_out_sel;
wire [0:0] RMUX_T1_WEST_B1_sel_value_O;
wire [0:0] RMUX_T2_EAST_B1_O;
wire RMUX_T2_EAST_B1_ready_out;
wire RMUX_T2_EAST_B1_valid_out;
wire [1:0] RMUX_T2_EAST_B1_out_sel;
wire [0:0] RMUX_T2_EAST_B1_sel_value_O;
wire [0:0] RMUX_T2_NORTH_B1_O;
wire RMUX_T2_NORTH_B1_ready_out;
wire RMUX_T2_NORTH_B1_valid_out;
wire [1:0] RMUX_T2_NORTH_B1_out_sel;
wire [0:0] RMUX_T2_NORTH_B1_sel_value_O;
wire [0:0] RMUX_T2_SOUTH_B1_O;
wire RMUX_T2_SOUTH_B1_ready_out;
wire RMUX_T2_SOUTH_B1_valid_out;
wire [1:0] RMUX_T2_SOUTH_B1_out_sel;
wire [0:0] RMUX_T2_SOUTH_B1_sel_value_O;
wire [0:0] RMUX_T2_WEST_B1_O;
wire RMUX_T2_WEST_B1_ready_out;
wire RMUX_T2_WEST_B1_valid_out;
wire [1:0] RMUX_T2_WEST_B1_out_sel;
wire [0:0] RMUX_T2_WEST_B1_sel_value_O;
wire [0:0] RMUX_T3_EAST_B1_O;
wire RMUX_T3_EAST_B1_ready_out;
wire RMUX_T3_EAST_B1_valid_out;
wire [1:0] RMUX_T3_EAST_B1_out_sel;
wire [0:0] RMUX_T3_EAST_B1_sel_value_O;
wire [0:0] RMUX_T3_NORTH_B1_O;
wire RMUX_T3_NORTH_B1_ready_out;
wire RMUX_T3_NORTH_B1_valid_out;
wire [1:0] RMUX_T3_NORTH_B1_out_sel;
wire [0:0] RMUX_T3_NORTH_B1_sel_value_O;
wire [0:0] RMUX_T3_SOUTH_B1_O;
wire RMUX_T3_SOUTH_B1_ready_out;
wire RMUX_T3_SOUTH_B1_valid_out;
wire [1:0] RMUX_T3_SOUTH_B1_out_sel;
wire [0:0] RMUX_T3_SOUTH_B1_sel_value_O;
wire [0:0] RMUX_T3_WEST_B1_O;
wire RMUX_T3_WEST_B1_ready_out;
wire RMUX_T3_WEST_B1_valid_out;
wire [1:0] RMUX_T3_WEST_B1_out_sel;
wire [0:0] RMUX_T3_WEST_B1_sel_value_O;
wire [0:0] RMUX_T4_EAST_B1_O;
wire RMUX_T4_EAST_B1_ready_out;
wire RMUX_T4_EAST_B1_valid_out;
wire [1:0] RMUX_T4_EAST_B1_out_sel;
wire [0:0] RMUX_T4_EAST_B1_sel_value_O;
wire [0:0] RMUX_T4_NORTH_B1_O;
wire RMUX_T4_NORTH_B1_ready_out;
wire RMUX_T4_NORTH_B1_valid_out;
wire [1:0] RMUX_T4_NORTH_B1_out_sel;
wire [0:0] RMUX_T4_NORTH_B1_sel_value_O;
wire [0:0] RMUX_T4_SOUTH_B1_O;
wire RMUX_T4_SOUTH_B1_ready_out;
wire RMUX_T4_SOUTH_B1_valid_out;
wire [1:0] RMUX_T4_SOUTH_B1_out_sel;
wire [0:0] RMUX_T4_SOUTH_B1_sel_value_O;
wire [0:0] RMUX_T4_WEST_B1_O;
wire RMUX_T4_WEST_B1_ready_out;
wire RMUX_T4_WEST_B1_valid_out;
wire [1:0] RMUX_T4_WEST_B1_out_sel;
wire [0:0] RMUX_T4_WEST_B1_sel_value_O;
wire [0:0] SB_T0_EAST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T0_EAST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T0_EAST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T0_EAST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T0_EAST_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T0_NORTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T0_NORTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T0_NORTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T0_NORTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T0_NORTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T0_SOUTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T0_SOUTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T0_SOUTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T0_SOUTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T0_SOUTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T0_WEST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T0_WEST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T0_WEST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T0_WEST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T0_WEST_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T1_EAST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T1_EAST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T1_EAST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T1_EAST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T1_EAST_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T1_NORTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T1_NORTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T1_NORTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T1_NORTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T1_NORTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T1_SOUTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T1_SOUTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T1_SOUTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T1_SOUTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T1_SOUTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T1_WEST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T1_WEST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T1_WEST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T1_WEST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T1_WEST_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T2_EAST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T2_EAST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T2_EAST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T2_EAST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T2_EAST_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T2_NORTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T2_NORTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T2_NORTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T2_NORTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T2_NORTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T2_SOUTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T2_SOUTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T2_SOUTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T2_SOUTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T2_SOUTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T2_WEST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T2_WEST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T2_WEST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T2_WEST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T2_WEST_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T3_EAST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T3_EAST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T3_EAST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T3_EAST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T3_EAST_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T3_NORTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T3_NORTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T3_NORTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T3_NORTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T3_NORTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T3_SOUTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T3_SOUTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T3_SOUTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T3_SOUTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T3_SOUTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T3_WEST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T3_WEST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T3_WEST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T3_WEST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T3_WEST_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T4_EAST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T4_EAST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T4_EAST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T4_EAST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T4_EAST_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T4_NORTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T4_NORTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T4_NORTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T4_NORTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T4_NORTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T4_SOUTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T4_SOUTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T4_SOUTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T4_SOUTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T4_SOUTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T4_WEST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T4_WEST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T4_WEST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T4_WEST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T4_WEST_SB_OUT_B1_sel_value_O;
wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1_O;
wire WIRE_SB_T0_EAST_SB_IN_B1_ready_out;
wire WIRE_SB_T0_EAST_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1_O;
wire WIRE_SB_T0_NORTH_SB_IN_B1_ready_out;
wire WIRE_SB_T0_NORTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1_O;
wire WIRE_SB_T0_SOUTH_SB_IN_B1_ready_out;
wire WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1_O;
wire WIRE_SB_T0_WEST_SB_IN_B1_ready_out;
wire WIRE_SB_T0_WEST_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1_O;
wire WIRE_SB_T1_EAST_SB_IN_B1_ready_out;
wire WIRE_SB_T1_EAST_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1_O;
wire WIRE_SB_T1_NORTH_SB_IN_B1_ready_out;
wire WIRE_SB_T1_NORTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1_O;
wire WIRE_SB_T1_SOUTH_SB_IN_B1_ready_out;
wire WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1_O;
wire WIRE_SB_T1_WEST_SB_IN_B1_ready_out;
wire WIRE_SB_T1_WEST_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1_O;
wire WIRE_SB_T2_EAST_SB_IN_B1_ready_out;
wire WIRE_SB_T2_EAST_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1_O;
wire WIRE_SB_T2_NORTH_SB_IN_B1_ready_out;
wire WIRE_SB_T2_NORTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1_O;
wire WIRE_SB_T2_SOUTH_SB_IN_B1_ready_out;
wire WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1_O;
wire WIRE_SB_T2_WEST_SB_IN_B1_ready_out;
wire WIRE_SB_T2_WEST_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1_O;
wire WIRE_SB_T3_EAST_SB_IN_B1_ready_out;
wire WIRE_SB_T3_EAST_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1_O;
wire WIRE_SB_T3_NORTH_SB_IN_B1_ready_out;
wire WIRE_SB_T3_NORTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1_O;
wire WIRE_SB_T3_SOUTH_SB_IN_B1_ready_out;
wire WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1_O;
wire WIRE_SB_T3_WEST_SB_IN_B1_ready_out;
wire WIRE_SB_T3_WEST_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1_O;
wire WIRE_SB_T4_EAST_SB_IN_B1_ready_out;
wire WIRE_SB_T4_EAST_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1_O;
wire WIRE_SB_T4_NORTH_SB_IN_B1_ready_out;
wire WIRE_SB_T4_NORTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1_O;
wire WIRE_SB_T4_SOUTH_SB_IN_B1_ready_out;
wire WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1_O;
wire WIRE_SB_T4_WEST_SB_IN_B1_ready_out;
wire WIRE_SB_T4_WEST_SB_IN_B1_valid_out;
wire ZextWrapper_23_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_23_32_inst0$self_O_in;
wire ZextWrapper_30_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_30_32_inst0$self_O_in;
wire ZextWrapper_31_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_31_32_inst0$self_O_in;
wire [0:0] and1_inst0_out;
wire [0:0] and1_inst1_out;
wire [0:0] and1_inst10_out;
wire [0:0] and1_inst11_out;
wire [0:0] and1_inst12_out;
wire [0:0] and1_inst13_out;
wire [0:0] and1_inst14_out;
wire [0:0] and1_inst15_out;
wire [0:0] and1_inst16_out;
wire [0:0] and1_inst17_out;
wire [0:0] and1_inst18_out;
wire [0:0] and1_inst19_out;
wire [0:0] and1_inst2_out;
wire [0:0] and1_inst3_out;
wire [0:0] and1_inst4_out;
wire [0:0] and1_inst5_out;
wire [0:0] and1_inst6_out;
wire [0:0] and1_inst7_out;
wire [0:0] and1_inst8_out;
wire [0:0] and1_inst9_out;
wire [31:0] config_reg_0_O;
wire [31:0] config_reg_1_O;
wire [31:0] config_reg_2_O;
wire [30:0] config_reg_3_O;
wire [29:0] config_reg_4_O;
wire [22:0] config_reg_5_O;
wire [0:0] const_0_1_out;
wire [31:0] const_0_32_out;
wire [0:0] const_1_1_out;
wire coreir_eq_1_inst0_out;
wire coreir_eq_1_inst1_out;
wire coreir_eq_1_inst10_out;
wire coreir_eq_1_inst11_out;
wire coreir_eq_1_inst12_out;
wire coreir_eq_1_inst13_out;
wire coreir_eq_1_inst14_out;
wire coreir_eq_1_inst15_out;
wire coreir_eq_1_inst16_out;
wire coreir_eq_1_inst17_out;
wire coreir_eq_1_inst18_out;
wire coreir_eq_1_inst19_out;
wire coreir_eq_1_inst2_out;
wire coreir_eq_1_inst3_out;
wire coreir_eq_1_inst4_out;
wire coreir_eq_1_inst5_out;
wire coreir_eq_1_inst6_out;
wire coreir_eq_1_inst7_out;
wire coreir_eq_1_inst8_out;
wire coreir_eq_1_inst9_out;
wire [31:0] mux_aoi_6_32_inst0_O;
wire [7:0] mux_aoi_6_32_inst0_out_sel;
wire [7:0] self_config_config_addr_out;
FanoutHash_E70AF988E4250F5 CB_PE_output_width_1_num_0_fan_in (
    .S13(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
    .E13(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
    .S6(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
    .E2(SB_T0_EAST_SB_OUT_B1_enable_value_O),
    .E12(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
    .E7(SB_T1_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
    .E18(SB_T4_EAST_SB_OUT_B1_enable_value_O),
    .I3(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
    .E19(SB_T4_WEST_SB_OUT_B1_enable_value_O),
    .I14(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
    .S14(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
    .I9(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
    .S12(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
    .S17(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
    .I13(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
    .S9(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
    .E10(SB_T2_EAST_SB_OUT_B1_enable_value_O),
    .E15(SB_T3_WEST_SB_OUT_B1_enable_value_O),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
    .E5(SB_T1_SOUTH_SB_OUT_B1_enable_value_O),
    .S10(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
    .E8(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
    .I11(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
    .I6(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
    .S15(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
    .I7(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
    .E14(SB_T3_EAST_SB_OUT_B1_enable_value_O),
    .I2(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
    .E11(SB_T2_WEST_SB_OUT_B1_enable_value_O),
    .S3(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
    .S8(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
    .I10(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
    .S16(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
    .E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
    .E16(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
    .E3(SB_T0_WEST_SB_OUT_B1_enable_value_O),
    .S18(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
    .S19(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
    .S2(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
    .S4(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
    .E9(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
    .I16(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
    .I12(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
    .S11(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
    .I17(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
    .I19(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
    .I18(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
    .S7(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
    .E4(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
    .E17(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
    .S5(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
    .I1(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
    .I5(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
    .E6(SB_T1_EAST_SB_OUT_B1_enable_value_O),
    .I4(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
    .I8(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
    .O(CB_PE_output_width_1_num_0_fan_in_O),
    .E1(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
    .I15(MUX_SB_T3_WEST_SB_OUT_B1_ready_out)
);
FanoutHash_F689C91787363AB CB_PondTop_output_width_1_num_0_fan_in (
    .S13(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
    .E13(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
    .S6(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
    .E2(SB_T0_EAST_SB_OUT_B1_enable_value_O),
    .E12(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
    .E7(SB_T1_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
    .E18(SB_T4_EAST_SB_OUT_B1_enable_value_O),
    .I3(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
    .E19(SB_T4_WEST_SB_OUT_B1_enable_value_O),
    .I14(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
    .S14(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
    .I9(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
    .S12(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
    .E20(PE_input_width_1_num_0_enable),
    .S17(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
    .I13(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
    .S9(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
    .E10(SB_T2_EAST_SB_OUT_B1_enable_value_O),
    .E15(SB_T3_WEST_SB_OUT_B1_enable_value_O),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
    .E5(SB_T1_SOUTH_SB_OUT_B1_enable_value_O),
    .S10(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
    .E8(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
    .I11(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
    .I6(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
    .S15(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
    .I20(PE_input_width_1_num_0_ready),
    .S20(PE_input_width_1_num_0_out_sel),
    .I7(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
    .E14(SB_T3_EAST_SB_OUT_B1_enable_value_O),
    .I2(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
    .E11(SB_T2_WEST_SB_OUT_B1_enable_value_O),
    .S3(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
    .S8(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
    .I10(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
    .S16(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
    .E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
    .E16(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
    .E3(SB_T0_WEST_SB_OUT_B1_enable_value_O),
    .S18(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
    .S19(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
    .S2(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
    .S4(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
    .E9(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
    .I16(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
    .I12(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
    .S11(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
    .I17(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
    .I19(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
    .I18(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
    .S7(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
    .E4(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
    .E17(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
    .S5(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
    .I1(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
    .I5(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
    .E6(SB_T1_EAST_SB_OUT_B1_enable_value_O),
    .I4(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
    .I8(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
    .O(CB_PondTop_output_width_1_num_0_fan_in_O),
    .E1(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
    .I15(MUX_SB_T3_WEST_SB_OUT_B1_ready_out)
);
FanoutHash_CE1AA874B742213 CB_PondTop_output_width_1_num_1_fan_in (
    .S13(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
    .E13(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
    .S6(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
    .E2(SB_T0_EAST_SB_OUT_B1_enable_value_O),
    .E12(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
    .E7(SB_T1_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
    .E18(SB_T4_EAST_SB_OUT_B1_enable_value_O),
    .I3(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
    .E19(SB_T4_WEST_SB_OUT_B1_enable_value_O),
    .I14(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
    .S14(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
    .I9(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
    .S12(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
    .S17(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
    .I13(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
    .S9(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
    .E10(SB_T2_EAST_SB_OUT_B1_enable_value_O),
    .E15(SB_T3_WEST_SB_OUT_B1_enable_value_O),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
    .E5(SB_T1_SOUTH_SB_OUT_B1_enable_value_O),
    .S10(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
    .E8(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
    .I11(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
    .I6(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
    .S15(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
    .I7(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
    .E14(SB_T3_EAST_SB_OUT_B1_enable_value_O),
    .I2(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
    .E11(SB_T2_WEST_SB_OUT_B1_enable_value_O),
    .S3(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
    .S8(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
    .I10(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
    .S16(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
    .E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
    .E16(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
    .E3(SB_T0_WEST_SB_OUT_B1_enable_value_O),
    .S18(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
    .S19(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
    .S2(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
    .S4(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
    .E9(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
    .I16(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
    .I12(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
    .S11(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
    .I17(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
    .I19(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
    .I18(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
    .S7(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
    .E4(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
    .E17(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
    .S5(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
    .I1(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
    .I5(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
    .E6(SB_T1_EAST_SB_OUT_B1_enable_value_O),
    .I4(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
    .I8(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
    .O(CB_PondTop_output_width_1_num_1_fan_in_O),
    .E1(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
    .I15(MUX_SB_T3_WEST_SB_OUT_B1_ready_out)
);
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(stall),
    .out(Invert1_inst0_out)
);
wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1_I [5:0];
assign MUX_SB_T0_EAST_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T0_EAST_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T0_EAST_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T0_EAST_SB_OUT_B1_I[2] = WIRE_SB_T4_NORTH_SB_IN_B1_O;
assign MUX_SB_T0_EAST_SB_OUT_B1_I[1] = WIRE_SB_T3_SOUTH_SB_IN_B1_O;
assign MUX_SB_T0_EAST_SB_OUT_B1_I[0] = WIRE_SB_T0_WEST_SB_IN_B1_O;
wire [5:0] MUX_SB_T0_EAST_SB_OUT_B1_valid_in;
assign MUX_SB_T0_EAST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T4_NORTH_SB_IN_B1_valid_out,WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T0_WEST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T0_EAST_SB_OUT_B1 (
    .I(MUX_SB_T0_EAST_SB_OUT_B1_I),
    .O(MUX_SB_T0_EAST_SB_OUT_B1_O),
    .ready_in(SB_T0_EAST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T0_EAST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T0_EAST_SB_OUT_B1_valid_out),
    .S(SB_T0_EAST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T0_EAST_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T0_NORTH_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T0_NORTH_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T0_NORTH_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T0_NORTH_SB_OUT_B1_I[2] = WIRE_SB_T0_SOUTH_SB_IN_B1_O;
assign MUX_SB_T0_NORTH_SB_OUT_B1_I[1] = WIRE_SB_T1_EAST_SB_IN_B1_O;
assign MUX_SB_T0_NORTH_SB_OUT_B1_I[0] = WIRE_SB_T0_WEST_SB_IN_B1_O;
wire [5:0] MUX_SB_T0_NORTH_SB_OUT_B1_valid_in;
assign MUX_SB_T0_NORTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T1_EAST_SB_IN_B1_valid_out,WIRE_SB_T0_WEST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T0_NORTH_SB_OUT_B1 (
    .I(MUX_SB_T0_NORTH_SB_OUT_B1_I),
    .O(MUX_SB_T0_NORTH_SB_OUT_B1_O),
    .ready_in(SB_T0_NORTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T0_NORTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T0_NORTH_SB_OUT_B1_valid_out),
    .S(SB_T0_NORTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[2] = WIRE_SB_T1_WEST_SB_IN_B1_O;
assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[1] = WIRE_SB_T0_NORTH_SB_IN_B1_O;
assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[0] = WIRE_SB_T3_EAST_SB_IN_B1_O;
wire [5:0] MUX_SB_T0_SOUTH_SB_OUT_B1_valid_in;
assign MUX_SB_T0_SOUTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T1_WEST_SB_IN_B1_valid_out,WIRE_SB_T0_NORTH_SB_IN_B1_valid_out,WIRE_SB_T3_EAST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T0_SOUTH_SB_OUT_B1 (
    .I(MUX_SB_T0_SOUTH_SB_OUT_B1_I),
    .O(MUX_SB_T0_SOUTH_SB_OUT_B1_O),
    .ready_in(SB_T0_SOUTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T0_SOUTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T0_SOUTH_SB_OUT_B1_valid_out),
    .S(SB_T0_SOUTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1_I [5:0];
assign MUX_SB_T0_WEST_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T0_WEST_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T0_WEST_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T0_WEST_SB_OUT_B1_I[2] = WIRE_SB_T0_EAST_SB_IN_B1_O;
assign MUX_SB_T0_WEST_SB_OUT_B1_I[1] = WIRE_SB_T4_SOUTH_SB_IN_B1_O;
assign MUX_SB_T0_WEST_SB_OUT_B1_I[0] = WIRE_SB_T0_NORTH_SB_IN_B1_O;
wire [5:0] MUX_SB_T0_WEST_SB_OUT_B1_valid_in;
assign MUX_SB_T0_WEST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T0_EAST_SB_IN_B1_valid_out,WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T0_NORTH_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T0_WEST_SB_OUT_B1 (
    .I(MUX_SB_T0_WEST_SB_OUT_B1_I),
    .O(MUX_SB_T0_WEST_SB_OUT_B1_O),
    .ready_in(SB_T0_WEST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T0_WEST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T0_WEST_SB_OUT_B1_valid_out),
    .S(SB_T0_WEST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T0_WEST_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1_I [5:0];
assign MUX_SB_T1_EAST_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T1_EAST_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T1_EAST_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T1_EAST_SB_OUT_B1_I[2] = WIRE_SB_T2_SOUTH_SB_IN_B1_O;
assign MUX_SB_T1_EAST_SB_OUT_B1_I[1] = WIRE_SB_T1_WEST_SB_IN_B1_O;
assign MUX_SB_T1_EAST_SB_OUT_B1_I[0] = WIRE_SB_T0_NORTH_SB_IN_B1_O;
wire [5:0] MUX_SB_T1_EAST_SB_OUT_B1_valid_in;
assign MUX_SB_T1_EAST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T1_WEST_SB_IN_B1_valid_out,WIRE_SB_T0_NORTH_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T1_EAST_SB_OUT_B1 (
    .I(MUX_SB_T1_EAST_SB_OUT_B1_I),
    .O(MUX_SB_T1_EAST_SB_OUT_B1_O),
    .ready_in(SB_T1_EAST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T1_EAST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T1_EAST_SB_OUT_B1_valid_out),
    .S(SB_T1_EAST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T1_EAST_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T1_NORTH_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T1_NORTH_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T1_NORTH_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T1_NORTH_SB_OUT_B1_I[2] = WIRE_SB_T4_WEST_SB_IN_B1_O;
assign MUX_SB_T1_NORTH_SB_OUT_B1_I[1] = WIRE_SB_T1_SOUTH_SB_IN_B1_O;
assign MUX_SB_T1_NORTH_SB_OUT_B1_I[0] = WIRE_SB_T2_EAST_SB_IN_B1_O;
wire [5:0] MUX_SB_T1_NORTH_SB_OUT_B1_valid_in;
assign MUX_SB_T1_NORTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T4_WEST_SB_IN_B1_valid_out,WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T2_EAST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T1_NORTH_SB_OUT_B1 (
    .I(MUX_SB_T1_NORTH_SB_OUT_B1_I),
    .O(MUX_SB_T1_NORTH_SB_OUT_B1_O),
    .ready_in(SB_T1_NORTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T1_NORTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T1_NORTH_SB_OUT_B1_valid_out),
    .S(SB_T1_NORTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[2] = WIRE_SB_T2_WEST_SB_IN_B1_O;
assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[1] = WIRE_SB_T1_NORTH_SB_IN_B1_O;
assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[0] = WIRE_SB_T2_EAST_SB_IN_B1_O;
wire [5:0] MUX_SB_T1_SOUTH_SB_OUT_B1_valid_in;
assign MUX_SB_T1_SOUTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T2_WEST_SB_IN_B1_valid_out,WIRE_SB_T1_NORTH_SB_IN_B1_valid_out,WIRE_SB_T2_EAST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T1_SOUTH_SB_OUT_B1 (
    .I(MUX_SB_T1_SOUTH_SB_OUT_B1_I),
    .O(MUX_SB_T1_SOUTH_SB_OUT_B1_O),
    .ready_in(SB_T1_SOUTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T1_SOUTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T1_SOUTH_SB_OUT_B1_valid_out),
    .S(SB_T1_SOUTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1_I [5:0];
assign MUX_SB_T1_WEST_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T1_WEST_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T1_WEST_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T1_WEST_SB_OUT_B1_I[2] = WIRE_SB_T1_EAST_SB_IN_B1_O;
assign MUX_SB_T1_WEST_SB_OUT_B1_I[1] = WIRE_SB_T0_SOUTH_SB_IN_B1_O;
assign MUX_SB_T1_WEST_SB_OUT_B1_I[0] = WIRE_SB_T4_NORTH_SB_IN_B1_O;
wire [5:0] MUX_SB_T1_WEST_SB_OUT_B1_valid_in;
assign MUX_SB_T1_WEST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T1_EAST_SB_IN_B1_valid_out,WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T4_NORTH_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T1_WEST_SB_OUT_B1 (
    .I(MUX_SB_T1_WEST_SB_OUT_B1_I),
    .O(MUX_SB_T1_WEST_SB_OUT_B1_O),
    .ready_in(SB_T1_WEST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T1_WEST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T1_WEST_SB_OUT_B1_valid_out),
    .S(SB_T1_WEST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T1_WEST_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1_I [5:0];
assign MUX_SB_T2_EAST_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T2_EAST_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T2_EAST_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T2_EAST_SB_OUT_B1_I[2] = WIRE_SB_T2_WEST_SB_IN_B1_O;
assign MUX_SB_T2_EAST_SB_OUT_B1_I[1] = WIRE_SB_T1_SOUTH_SB_IN_B1_O;
assign MUX_SB_T2_EAST_SB_OUT_B1_I[0] = WIRE_SB_T1_NORTH_SB_IN_B1_O;
wire [5:0] MUX_SB_T2_EAST_SB_OUT_B1_valid_in;
assign MUX_SB_T2_EAST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T2_WEST_SB_IN_B1_valid_out,WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T1_NORTH_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T2_EAST_SB_OUT_B1 (
    .I(MUX_SB_T2_EAST_SB_OUT_B1_I),
    .O(MUX_SB_T2_EAST_SB_OUT_B1_O),
    .ready_in(SB_T2_EAST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T2_EAST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T2_EAST_SB_OUT_B1_valid_out),
    .S(SB_T2_EAST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T2_EAST_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T2_NORTH_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T2_NORTH_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T2_NORTH_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T2_NORTH_SB_OUT_B1_I[2] = WIRE_SB_T3_WEST_SB_IN_B1_O;
assign MUX_SB_T2_NORTH_SB_OUT_B1_I[1] = WIRE_SB_T2_SOUTH_SB_IN_B1_O;
assign MUX_SB_T2_NORTH_SB_OUT_B1_I[0] = WIRE_SB_T3_EAST_SB_IN_B1_O;
wire [5:0] MUX_SB_T2_NORTH_SB_OUT_B1_valid_in;
assign MUX_SB_T2_NORTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T3_WEST_SB_IN_B1_valid_out,WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T3_EAST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T2_NORTH_SB_OUT_B1 (
    .I(MUX_SB_T2_NORTH_SB_OUT_B1_I),
    .O(MUX_SB_T2_NORTH_SB_OUT_B1_O),
    .ready_in(SB_T2_NORTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T2_NORTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T2_NORTH_SB_OUT_B1_valid_out),
    .S(SB_T2_NORTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[2] = WIRE_SB_T3_WEST_SB_IN_B1_O;
assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[1] = WIRE_SB_T2_NORTH_SB_IN_B1_O;
assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[0] = WIRE_SB_T1_EAST_SB_IN_B1_O;
wire [5:0] MUX_SB_T2_SOUTH_SB_OUT_B1_valid_in;
assign MUX_SB_T2_SOUTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T3_WEST_SB_IN_B1_valid_out,WIRE_SB_T2_NORTH_SB_IN_B1_valid_out,WIRE_SB_T1_EAST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T2_SOUTH_SB_OUT_B1 (
    .I(MUX_SB_T2_SOUTH_SB_OUT_B1_I),
    .O(MUX_SB_T2_SOUTH_SB_OUT_B1_O),
    .ready_in(SB_T2_SOUTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T2_SOUTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T2_SOUTH_SB_OUT_B1_valid_out),
    .S(SB_T2_SOUTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1_I [5:0];
assign MUX_SB_T2_WEST_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T2_WEST_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T2_WEST_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T2_WEST_SB_OUT_B1_I[2] = WIRE_SB_T2_EAST_SB_IN_B1_O;
assign MUX_SB_T2_WEST_SB_OUT_B1_I[1] = WIRE_SB_T1_SOUTH_SB_IN_B1_O;
assign MUX_SB_T2_WEST_SB_OUT_B1_I[0] = WIRE_SB_T3_NORTH_SB_IN_B1_O;
wire [5:0] MUX_SB_T2_WEST_SB_OUT_B1_valid_in;
assign MUX_SB_T2_WEST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T2_EAST_SB_IN_B1_valid_out,WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T3_NORTH_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T2_WEST_SB_OUT_B1 (
    .I(MUX_SB_T2_WEST_SB_OUT_B1_I),
    .O(MUX_SB_T2_WEST_SB_OUT_B1_O),
    .ready_in(SB_T2_WEST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T2_WEST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T2_WEST_SB_OUT_B1_valid_out),
    .S(SB_T2_WEST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T2_WEST_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1_I [5:0];
assign MUX_SB_T3_EAST_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T3_EAST_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T3_EAST_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T3_EAST_SB_OUT_B1_I[2] = WIRE_SB_T3_WEST_SB_IN_B1_O;
assign MUX_SB_T3_EAST_SB_OUT_B1_I[1] = WIRE_SB_T2_NORTH_SB_IN_B1_O;
assign MUX_SB_T3_EAST_SB_OUT_B1_I[0] = WIRE_SB_T0_SOUTH_SB_IN_B1_O;
wire [5:0] MUX_SB_T3_EAST_SB_OUT_B1_valid_in;
assign MUX_SB_T3_EAST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T3_WEST_SB_IN_B1_valid_out,WIRE_SB_T2_NORTH_SB_IN_B1_valid_out,WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T3_EAST_SB_OUT_B1 (
    .I(MUX_SB_T3_EAST_SB_OUT_B1_I),
    .O(MUX_SB_T3_EAST_SB_OUT_B1_O),
    .ready_in(SB_T3_EAST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T3_EAST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T3_EAST_SB_OUT_B1_valid_out),
    .S(SB_T3_EAST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T3_EAST_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T3_NORTH_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T3_NORTH_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T3_NORTH_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T3_NORTH_SB_OUT_B1_I[2] = WIRE_SB_T3_SOUTH_SB_IN_B1_O;
assign MUX_SB_T3_NORTH_SB_OUT_B1_I[1] = WIRE_SB_T4_EAST_SB_IN_B1_O;
assign MUX_SB_T3_NORTH_SB_OUT_B1_I[0] = WIRE_SB_T2_WEST_SB_IN_B1_O;
wire [5:0] MUX_SB_T3_NORTH_SB_OUT_B1_valid_in;
assign MUX_SB_T3_NORTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T4_EAST_SB_IN_B1_valid_out,WIRE_SB_T2_WEST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T3_NORTH_SB_OUT_B1 (
    .I(MUX_SB_T3_NORTH_SB_OUT_B1_I),
    .O(MUX_SB_T3_NORTH_SB_OUT_B1_O),
    .ready_in(SB_T3_NORTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T3_NORTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T3_NORTH_SB_OUT_B1_valid_out),
    .S(SB_T3_NORTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[2] = WIRE_SB_T4_WEST_SB_IN_B1_O;
assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[1] = WIRE_SB_T3_NORTH_SB_IN_B1_O;
assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[0] = WIRE_SB_T0_EAST_SB_IN_B1_O;
wire [5:0] MUX_SB_T3_SOUTH_SB_OUT_B1_valid_in;
assign MUX_SB_T3_SOUTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T4_WEST_SB_IN_B1_valid_out,WIRE_SB_T3_NORTH_SB_IN_B1_valid_out,WIRE_SB_T0_EAST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T3_SOUTH_SB_OUT_B1 (
    .I(MUX_SB_T3_SOUTH_SB_OUT_B1_I),
    .O(MUX_SB_T3_SOUTH_SB_OUT_B1_O),
    .ready_in(SB_T3_SOUTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T3_SOUTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T3_SOUTH_SB_OUT_B1_valid_out),
    .S(SB_T3_SOUTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1_I [5:0];
assign MUX_SB_T3_WEST_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T3_WEST_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T3_WEST_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T3_WEST_SB_OUT_B1_I[2] = WIRE_SB_T3_EAST_SB_IN_B1_O;
assign MUX_SB_T3_WEST_SB_OUT_B1_I[1] = WIRE_SB_T2_SOUTH_SB_IN_B1_O;
assign MUX_SB_T3_WEST_SB_OUT_B1_I[0] = WIRE_SB_T2_NORTH_SB_IN_B1_O;
wire [5:0] MUX_SB_T3_WEST_SB_OUT_B1_valid_in;
assign MUX_SB_T3_WEST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T3_EAST_SB_IN_B1_valid_out,WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T2_NORTH_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T3_WEST_SB_OUT_B1 (
    .I(MUX_SB_T3_WEST_SB_OUT_B1_I),
    .O(MUX_SB_T3_WEST_SB_OUT_B1_O),
    .ready_in(SB_T3_WEST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T3_WEST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T3_WEST_SB_OUT_B1_valid_out),
    .S(SB_T3_WEST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T3_WEST_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1_I [5:0];
assign MUX_SB_T4_EAST_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T4_EAST_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T4_EAST_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T4_EAST_SB_OUT_B1_I[2] = WIRE_SB_T4_WEST_SB_IN_B1_O;
assign MUX_SB_T4_EAST_SB_OUT_B1_I[1] = WIRE_SB_T4_SOUTH_SB_IN_B1_O;
assign MUX_SB_T4_EAST_SB_OUT_B1_I[0] = WIRE_SB_T3_NORTH_SB_IN_B1_O;
wire [5:0] MUX_SB_T4_EAST_SB_OUT_B1_valid_in;
assign MUX_SB_T4_EAST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T4_WEST_SB_IN_B1_valid_out,WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T3_NORTH_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T4_EAST_SB_OUT_B1 (
    .I(MUX_SB_T4_EAST_SB_OUT_B1_I),
    .O(MUX_SB_T4_EAST_SB_OUT_B1_O),
    .ready_in(SB_T4_EAST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T4_EAST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T4_EAST_SB_OUT_B1_valid_out),
    .S(SB_T4_EAST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T4_EAST_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T4_NORTH_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T4_NORTH_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T4_NORTH_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T4_NORTH_SB_OUT_B1_I[2] = WIRE_SB_T4_SOUTH_SB_IN_B1_O;
assign MUX_SB_T4_NORTH_SB_OUT_B1_I[1] = WIRE_SB_T0_EAST_SB_IN_B1_O;
assign MUX_SB_T4_NORTH_SB_OUT_B1_I[0] = WIRE_SB_T1_WEST_SB_IN_B1_O;
wire [5:0] MUX_SB_T4_NORTH_SB_OUT_B1_valid_in;
assign MUX_SB_T4_NORTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T0_EAST_SB_IN_B1_valid_out,WIRE_SB_T1_WEST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T4_NORTH_SB_OUT_B1 (
    .I(MUX_SB_T4_NORTH_SB_OUT_B1_I),
    .O(MUX_SB_T4_NORTH_SB_OUT_B1_O),
    .ready_in(SB_T4_NORTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T4_NORTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T4_NORTH_SB_OUT_B1_valid_out),
    .S(SB_T4_NORTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[2] = WIRE_SB_T4_NORTH_SB_IN_B1_O;
assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[1] = WIRE_SB_T4_EAST_SB_IN_B1_O;
assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[0] = WIRE_SB_T0_WEST_SB_IN_B1_O;
wire [5:0] MUX_SB_T4_SOUTH_SB_OUT_B1_valid_in;
assign MUX_SB_T4_SOUTH_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T4_NORTH_SB_IN_B1_valid_out,WIRE_SB_T4_EAST_SB_IN_B1_valid_out,WIRE_SB_T0_WEST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T4_SOUTH_SB_OUT_B1 (
    .I(MUX_SB_T4_SOUTH_SB_OUT_B1_I),
    .O(MUX_SB_T4_SOUTH_SB_OUT_B1_O),
    .ready_in(SB_T4_SOUTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T4_SOUTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T4_SOUTH_SB_OUT_B1_valid_out),
    .S(SB_T4_SOUTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1_I [5:0];
assign MUX_SB_T4_WEST_SB_OUT_B1_I[5] = PondTop_output_width_1_num_1;
assign MUX_SB_T4_WEST_SB_OUT_B1_I[4] = PondTop_output_width_1_num_0;
assign MUX_SB_T4_WEST_SB_OUT_B1_I[3] = PE_output_width_1_num_0;
assign MUX_SB_T4_WEST_SB_OUT_B1_I[2] = WIRE_SB_T4_EAST_SB_IN_B1_O;
assign MUX_SB_T4_WEST_SB_OUT_B1_I[1] = WIRE_SB_T3_SOUTH_SB_IN_B1_O;
assign MUX_SB_T4_WEST_SB_OUT_B1_I[0] = WIRE_SB_T1_NORTH_SB_IN_B1_O;
wire [5:0] MUX_SB_T4_WEST_SB_OUT_B1_valid_in;
assign MUX_SB_T4_WEST_SB_OUT_B1_valid_in = {PondTop_output_width_1_num_1_valid,PondTop_output_width_1_num_0_valid,PE_output_width_1_num_0_valid,WIRE_SB_T4_EAST_SB_IN_B1_valid_out,WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T1_NORTH_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T4_WEST_SB_OUT_B1 (
    .I(MUX_SB_T4_WEST_SB_OUT_B1_I),
    .O(MUX_SB_T4_WEST_SB_OUT_B1_O),
    .ready_in(SB_T4_WEST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T4_WEST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T4_WEST_SB_OUT_B1_valid_out),
    .S(SB_T4_WEST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T4_WEST_SB_OUT_B1_out_sel)
);
SplitFifo_1 REG_T0_EAST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T0_EAST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T0_EAST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T0_EAST_B1_fifo_value_O[0]),
    .end_fifo(REG_T0_EAST_B1_end_value_O[0]),
    .data_in(MUX_SB_T0_EAST_SB_OUT_B1_O),
    .ready1(RMUX_T0_EAST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T0_EAST_SB_OUT_B1_valid_out),
    .data_out(REG_T0_EAST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T0_EAST_B1_start_value_O[0]),
    .clk_en(and1_inst2_out[0])
);
SliceWrapper_32_0_1 REG_T0_EAST_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T0_EAST_B1_end_value_O)
);
SliceWrapper_32_1_2 REG_T0_EAST_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T0_EAST_B1_fifo_value_O)
);
SliceWrapper_32_2_3 REG_T0_EAST_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T0_EAST_B1_start_value_O)
);
SplitFifo_1 REG_T0_NORTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T0_NORTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T0_NORTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T0_NORTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T0_NORTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T0_NORTH_SB_OUT_B1_O),
    .ready1(RMUX_T0_NORTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T0_NORTH_SB_OUT_B1_valid_out),
    .data_out(REG_T0_NORTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T0_NORTH_B1_start_value_O[0]),
    .clk_en(and1_inst0_out[0])
);
SliceWrapper_32_3_4 REG_T0_NORTH_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T0_NORTH_B1_end_value_O)
);
SliceWrapper_32_4_5 REG_T0_NORTH_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T0_NORTH_B1_fifo_value_O)
);
SliceWrapper_32_5_6 REG_T0_NORTH_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T0_NORTH_B1_start_value_O)
);
SplitFifo_1 REG_T0_SOUTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T0_SOUTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T0_SOUTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T0_SOUTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T0_SOUTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T0_SOUTH_SB_OUT_B1_O),
    .ready1(RMUX_T0_SOUTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T0_SOUTH_SB_OUT_B1_valid_out),
    .data_out(REG_T0_SOUTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T0_SOUTH_B1_start_value_O[0]),
    .clk_en(and1_inst1_out[0])
);
SliceWrapper_32_6_7 REG_T0_SOUTH_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T0_SOUTH_B1_end_value_O)
);
SliceWrapper_32_7_8 REG_T0_SOUTH_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T0_SOUTH_B1_fifo_value_O)
);
SliceWrapper_32_8_9 REG_T0_SOUTH_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T0_SOUTH_B1_start_value_O)
);
SplitFifo_1 REG_T0_WEST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T0_WEST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T0_WEST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T0_WEST_B1_fifo_value_O[0]),
    .end_fifo(REG_T0_WEST_B1_end_value_O[0]),
    .data_in(MUX_SB_T0_WEST_SB_OUT_B1_O),
    .ready1(RMUX_T0_WEST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T0_WEST_SB_OUT_B1_valid_out),
    .data_out(REG_T0_WEST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T0_WEST_B1_start_value_O[0]),
    .clk_en(and1_inst3_out[0])
);
SliceWrapper_32_9_10 REG_T0_WEST_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T0_WEST_B1_end_value_O)
);
SliceWrapper_32_10_11 REG_T0_WEST_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T0_WEST_B1_fifo_value_O)
);
SliceWrapper_32_11_12 REG_T0_WEST_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T0_WEST_B1_start_value_O)
);
SplitFifo_1 REG_T1_EAST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T1_EAST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T1_EAST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T1_EAST_B1_fifo_value_O[0]),
    .end_fifo(REG_T1_EAST_B1_end_value_O[0]),
    .data_in(MUX_SB_T1_EAST_SB_OUT_B1_O),
    .ready1(RMUX_T1_EAST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T1_EAST_SB_OUT_B1_valid_out),
    .data_out(REG_T1_EAST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T1_EAST_B1_start_value_O[0]),
    .clk_en(and1_inst6_out[0])
);
SliceWrapper_32_12_13 REG_T1_EAST_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T1_EAST_B1_end_value_O)
);
SliceWrapper_32_13_14 REG_T1_EAST_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T1_EAST_B1_fifo_value_O)
);
SliceWrapper_32_14_15 REG_T1_EAST_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T1_EAST_B1_start_value_O)
);
SplitFifo_1 REG_T1_NORTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T1_NORTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T1_NORTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T1_NORTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T1_NORTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T1_NORTH_SB_OUT_B1_O),
    .ready1(RMUX_T1_NORTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T1_NORTH_SB_OUT_B1_valid_out),
    .data_out(REG_T1_NORTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T1_NORTH_B1_start_value_O[0]),
    .clk_en(and1_inst4_out[0])
);
SliceWrapper_32_15_16 REG_T1_NORTH_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T1_NORTH_B1_end_value_O)
);
SliceWrapper_32_16_17 REG_T1_NORTH_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T1_NORTH_B1_fifo_value_O)
);
SliceWrapper_32_17_18 REG_T1_NORTH_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T1_NORTH_B1_start_value_O)
);
SplitFifo_1 REG_T1_SOUTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T1_SOUTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T1_SOUTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T1_SOUTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T1_SOUTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T1_SOUTH_SB_OUT_B1_O),
    .ready1(RMUX_T1_SOUTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T1_SOUTH_SB_OUT_B1_valid_out),
    .data_out(REG_T1_SOUTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T1_SOUTH_B1_start_value_O[0]),
    .clk_en(and1_inst5_out[0])
);
SliceWrapper_32_18_19 REG_T1_SOUTH_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T1_SOUTH_B1_end_value_O)
);
SliceWrapper_32_19_20 REG_T1_SOUTH_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T1_SOUTH_B1_fifo_value_O)
);
SliceWrapper_32_20_21 REG_T1_SOUTH_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T1_SOUTH_B1_start_value_O)
);
SplitFifo_1 REG_T1_WEST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T1_WEST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T1_WEST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T1_WEST_B1_fifo_value_O[0]),
    .end_fifo(REG_T1_WEST_B1_end_value_O[0]),
    .data_in(MUX_SB_T1_WEST_SB_OUT_B1_O),
    .ready1(RMUX_T1_WEST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T1_WEST_SB_OUT_B1_valid_out),
    .data_out(REG_T1_WEST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T1_WEST_B1_start_value_O[0]),
    .clk_en(and1_inst7_out[0])
);
SliceWrapper_32_21_22 REG_T1_WEST_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T1_WEST_B1_end_value_O)
);
SliceWrapper_32_22_23 REG_T1_WEST_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T1_WEST_B1_fifo_value_O)
);
SliceWrapper_32_23_24 REG_T1_WEST_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T1_WEST_B1_start_value_O)
);
SplitFifo_1 REG_T2_EAST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T2_EAST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T2_EAST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T2_EAST_B1_fifo_value_O[0]),
    .end_fifo(REG_T2_EAST_B1_end_value_O[0]),
    .data_in(MUX_SB_T2_EAST_SB_OUT_B1_O),
    .ready1(RMUX_T2_EAST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T2_EAST_SB_OUT_B1_valid_out),
    .data_out(REG_T2_EAST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T2_EAST_B1_start_value_O[0]),
    .clk_en(and1_inst10_out[0])
);
SliceWrapper_32_24_25 REG_T2_EAST_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T2_EAST_B1_end_value_O)
);
SliceWrapper_32_25_26 REG_T2_EAST_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T2_EAST_B1_fifo_value_O)
);
SliceWrapper_32_26_27 REG_T2_EAST_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T2_EAST_B1_start_value_O)
);
SplitFifo_1 REG_T2_NORTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T2_NORTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T2_NORTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T2_NORTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T2_NORTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T2_NORTH_SB_OUT_B1_O),
    .ready1(RMUX_T2_NORTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T2_NORTH_SB_OUT_B1_valid_out),
    .data_out(REG_T2_NORTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T2_NORTH_B1_start_value_O[0]),
    .clk_en(and1_inst8_out[0])
);
SliceWrapper_32_27_28 REG_T2_NORTH_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T2_NORTH_B1_end_value_O)
);
SliceWrapper_32_28_29 REG_T2_NORTH_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T2_NORTH_B1_fifo_value_O)
);
SliceWrapper_32_29_30 REG_T2_NORTH_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T2_NORTH_B1_start_value_O)
);
SplitFifo_1 REG_T2_SOUTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T2_SOUTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T2_SOUTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T2_SOUTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T2_SOUTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T2_SOUTH_SB_OUT_B1_O),
    .ready1(RMUX_T2_SOUTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T2_SOUTH_SB_OUT_B1_valid_out),
    .data_out(REG_T2_SOUTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T2_SOUTH_B1_start_value_O[0]),
    .clk_en(and1_inst9_out[0])
);
SliceWrapper_32_30_31 REG_T2_SOUTH_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T2_SOUTH_B1_end_value_O)
);
SliceWrapper_32_31_32 REG_T2_SOUTH_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T2_SOUTH_B1_fifo_value_O)
);
SliceWrapper_32_0_1 REG_T2_SOUTH_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T2_SOUTH_B1_start_value_O)
);
SplitFifo_1 REG_T2_WEST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T2_WEST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T2_WEST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T2_WEST_B1_fifo_value_O[0]),
    .end_fifo(REG_T2_WEST_B1_end_value_O[0]),
    .data_in(MUX_SB_T2_WEST_SB_OUT_B1_O),
    .ready1(RMUX_T2_WEST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T2_WEST_SB_OUT_B1_valid_out),
    .data_out(REG_T2_WEST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T2_WEST_B1_start_value_O[0]),
    .clk_en(and1_inst11_out[0])
);
SliceWrapper_32_1_2 REG_T2_WEST_B1_end_value (
    .I(config_reg_1_O),
    .O(REG_T2_WEST_B1_end_value_O)
);
SliceWrapper_32_2_3 REG_T2_WEST_B1_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T2_WEST_B1_fifo_value_O)
);
SliceWrapper_32_3_4 REG_T2_WEST_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T2_WEST_B1_start_value_O)
);
SplitFifo_1 REG_T3_EAST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T3_EAST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T3_EAST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T3_EAST_B1_fifo_value_O[0]),
    .end_fifo(REG_T3_EAST_B1_end_value_O[0]),
    .data_in(MUX_SB_T3_EAST_SB_OUT_B1_O),
    .ready1(RMUX_T3_EAST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T3_EAST_SB_OUT_B1_valid_out),
    .data_out(REG_T3_EAST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T3_EAST_B1_start_value_O[0]),
    .clk_en(and1_inst14_out[0])
);
SliceWrapper_32_4_5 REG_T3_EAST_B1_end_value (
    .I(config_reg_1_O),
    .O(REG_T3_EAST_B1_end_value_O)
);
SliceWrapper_32_5_6 REG_T3_EAST_B1_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T3_EAST_B1_fifo_value_O)
);
SliceWrapper_32_6_7 REG_T3_EAST_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T3_EAST_B1_start_value_O)
);
SplitFifo_1 REG_T3_NORTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T3_NORTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T3_NORTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T3_NORTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T3_NORTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T3_NORTH_SB_OUT_B1_O),
    .ready1(RMUX_T3_NORTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T3_NORTH_SB_OUT_B1_valid_out),
    .data_out(REG_T3_NORTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T3_NORTH_B1_start_value_O[0]),
    .clk_en(and1_inst12_out[0])
);
SliceWrapper_32_7_8 REG_T3_NORTH_B1_end_value (
    .I(config_reg_1_O),
    .O(REG_T3_NORTH_B1_end_value_O)
);
SliceWrapper_32_8_9 REG_T3_NORTH_B1_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T3_NORTH_B1_fifo_value_O)
);
SliceWrapper_32_9_10 REG_T3_NORTH_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T3_NORTH_B1_start_value_O)
);
SplitFifo_1 REG_T3_SOUTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T3_SOUTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T3_SOUTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T3_SOUTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T3_SOUTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T3_SOUTH_SB_OUT_B1_O),
    .ready1(RMUX_T3_SOUTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T3_SOUTH_SB_OUT_B1_valid_out),
    .data_out(REG_T3_SOUTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T3_SOUTH_B1_start_value_O[0]),
    .clk_en(and1_inst13_out[0])
);
SliceWrapper_32_10_11 REG_T3_SOUTH_B1_end_value (
    .I(config_reg_1_O),
    .O(REG_T3_SOUTH_B1_end_value_O)
);
SliceWrapper_32_11_12 REG_T3_SOUTH_B1_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T3_SOUTH_B1_fifo_value_O)
);
SliceWrapper_32_12_13 REG_T3_SOUTH_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T3_SOUTH_B1_start_value_O)
);
SplitFifo_1 REG_T3_WEST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T3_WEST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T3_WEST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T3_WEST_B1_fifo_value_O[0]),
    .end_fifo(REG_T3_WEST_B1_end_value_O[0]),
    .data_in(MUX_SB_T3_WEST_SB_OUT_B1_O),
    .ready1(RMUX_T3_WEST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T3_WEST_SB_OUT_B1_valid_out),
    .data_out(REG_T3_WEST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T3_WEST_B1_start_value_O[0]),
    .clk_en(and1_inst15_out[0])
);
SliceWrapper_32_13_14 REG_T3_WEST_B1_end_value (
    .I(config_reg_1_O),
    .O(REG_T3_WEST_B1_end_value_O)
);
SliceWrapper_32_14_15 REG_T3_WEST_B1_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T3_WEST_B1_fifo_value_O)
);
SliceWrapper_32_15_16 REG_T3_WEST_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T3_WEST_B1_start_value_O)
);
SplitFifo_1 REG_T4_EAST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T4_EAST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T4_EAST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T4_EAST_B1_fifo_value_O[0]),
    .end_fifo(REG_T4_EAST_B1_end_value_O[0]),
    .data_in(MUX_SB_T4_EAST_SB_OUT_B1_O),
    .ready1(RMUX_T4_EAST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T4_EAST_SB_OUT_B1_valid_out),
    .data_out(REG_T4_EAST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T4_EAST_B1_start_value_O[0]),
    .clk_en(and1_inst18_out[0])
);
SliceWrapper_32_16_17 REG_T4_EAST_B1_end_value (
    .I(config_reg_1_O),
    .O(REG_T4_EAST_B1_end_value_O)
);
SliceWrapper_32_17_18 REG_T4_EAST_B1_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T4_EAST_B1_fifo_value_O)
);
SliceWrapper_32_18_19 REG_T4_EAST_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T4_EAST_B1_start_value_O)
);
SplitFifo_1 REG_T4_NORTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T4_NORTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T4_NORTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T4_NORTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T4_NORTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T4_NORTH_SB_OUT_B1_O),
    .ready1(RMUX_T4_NORTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T4_NORTH_SB_OUT_B1_valid_out),
    .data_out(REG_T4_NORTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T4_NORTH_B1_start_value_O[0]),
    .clk_en(and1_inst16_out[0])
);
SliceWrapper_32_19_20 REG_T4_NORTH_B1_end_value (
    .I(config_reg_1_O),
    .O(REG_T4_NORTH_B1_end_value_O)
);
SliceWrapper_32_20_21 REG_T4_NORTH_B1_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T4_NORTH_B1_fifo_value_O)
);
SliceWrapper_32_21_22 REG_T4_NORTH_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T4_NORTH_B1_start_value_O)
);
SplitFifo_1 REG_T4_SOUTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T4_SOUTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T4_SOUTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T4_SOUTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T4_SOUTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T4_SOUTH_SB_OUT_B1_O),
    .ready1(RMUX_T4_SOUTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T4_SOUTH_SB_OUT_B1_valid_out),
    .data_out(REG_T4_SOUTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T4_SOUTH_B1_start_value_O[0]),
    .clk_en(and1_inst17_out[0])
);
SliceWrapper_32_22_23 REG_T4_SOUTH_B1_end_value (
    .I(config_reg_1_O),
    .O(REG_T4_SOUTH_B1_end_value_O)
);
SliceWrapper_32_23_24 REG_T4_SOUTH_B1_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T4_SOUTH_B1_fifo_value_O)
);
SliceWrapper_32_24_25 REG_T4_SOUTH_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T4_SOUTH_B1_start_value_O)
);
SplitFifo_1 REG_T4_WEST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T4_WEST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T4_WEST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T4_WEST_B1_fifo_value_O[0]),
    .end_fifo(REG_T4_WEST_B1_end_value_O[0]),
    .data_in(MUX_SB_T4_WEST_SB_OUT_B1_O),
    .ready1(RMUX_T4_WEST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T4_WEST_SB_OUT_B1_valid_out),
    .data_out(REG_T4_WEST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T4_WEST_B1_start_value_O[0]),
    .clk_en(and1_inst19_out[0])
);
SliceWrapper_32_25_26 REG_T4_WEST_B1_end_value (
    .I(config_reg_1_O),
    .O(REG_T4_WEST_B1_end_value_O)
);
SliceWrapper_32_26_27 REG_T4_WEST_B1_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T4_WEST_B1_fifo_value_O)
);
SliceWrapper_32_27_28 REG_T4_WEST_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T4_WEST_B1_start_value_O)
);
wire [0:0] RMUX_T0_EAST_B1_I [1:0];
assign RMUX_T0_EAST_B1_I[1] = REG_T0_EAST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T0_EAST_B1_I[0] = MUX_SB_T0_EAST_SB_OUT_B1_O;
wire [1:0] RMUX_T0_EAST_B1_valid_in;
assign RMUX_T0_EAST_B1_valid_in = {REG_T0_EAST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T0_EAST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T0_EAST_B1 (
    .I(RMUX_T0_EAST_B1_I),
    .O(RMUX_T0_EAST_B1_O),
    .ready_in(SB_T0_EAST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T0_EAST_B1_ready_out),
    .valid_in(RMUX_T0_EAST_B1_valid_in),
    .valid_out(RMUX_T0_EAST_B1_valid_out),
    .S(RMUX_T0_EAST_B1_sel_value_O),
    .out_sel(RMUX_T0_EAST_B1_out_sel)
);
SliceWrapper_32_28_29 RMUX_T0_EAST_B1_sel_value (
    .I(config_reg_1_O),
    .O(RMUX_T0_EAST_B1_sel_value_O)
);
wire [0:0] RMUX_T0_NORTH_B1_I [1:0];
assign RMUX_T0_NORTH_B1_I[1] = REG_T0_NORTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T0_NORTH_B1_I[0] = MUX_SB_T0_NORTH_SB_OUT_B1_O;
wire [1:0] RMUX_T0_NORTH_B1_valid_in;
assign RMUX_T0_NORTH_B1_valid_in = {REG_T0_NORTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T0_NORTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T0_NORTH_B1 (
    .I(RMUX_T0_NORTH_B1_I),
    .O(RMUX_T0_NORTH_B1_O),
    .ready_in(SB_T0_NORTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T0_NORTH_B1_ready_out),
    .valid_in(RMUX_T0_NORTH_B1_valid_in),
    .valid_out(RMUX_T0_NORTH_B1_valid_out),
    .S(RMUX_T0_NORTH_B1_sel_value_O),
    .out_sel(RMUX_T0_NORTH_B1_out_sel)
);
SliceWrapper_32_29_30 RMUX_T0_NORTH_B1_sel_value (
    .I(config_reg_1_O),
    .O(RMUX_T0_NORTH_B1_sel_value_O)
);
wire [0:0] RMUX_T0_SOUTH_B1_I [1:0];
assign RMUX_T0_SOUTH_B1_I[1] = REG_T0_SOUTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T0_SOUTH_B1_I[0] = MUX_SB_T0_SOUTH_SB_OUT_B1_O;
wire [1:0] RMUX_T0_SOUTH_B1_valid_in;
assign RMUX_T0_SOUTH_B1_valid_in = {REG_T0_SOUTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T0_SOUTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T0_SOUTH_B1 (
    .I(RMUX_T0_SOUTH_B1_I),
    .O(RMUX_T0_SOUTH_B1_O),
    .ready_in(SB_T0_SOUTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T0_SOUTH_B1_ready_out),
    .valid_in(RMUX_T0_SOUTH_B1_valid_in),
    .valid_out(RMUX_T0_SOUTH_B1_valid_out),
    .S(RMUX_T0_SOUTH_B1_sel_value_O),
    .out_sel(RMUX_T0_SOUTH_B1_out_sel)
);
SliceWrapper_32_30_31 RMUX_T0_SOUTH_B1_sel_value (
    .I(config_reg_1_O),
    .O(RMUX_T0_SOUTH_B1_sel_value_O)
);
wire [0:0] RMUX_T0_WEST_B1_I [1:0];
assign RMUX_T0_WEST_B1_I[1] = REG_T0_WEST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T0_WEST_B1_I[0] = MUX_SB_T0_WEST_SB_OUT_B1_O;
wire [1:0] RMUX_T0_WEST_B1_valid_in;
assign RMUX_T0_WEST_B1_valid_in = {REG_T0_WEST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T0_WEST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T0_WEST_B1 (
    .I(RMUX_T0_WEST_B1_I),
    .O(RMUX_T0_WEST_B1_O),
    .ready_in(SB_T0_WEST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T0_WEST_B1_ready_out),
    .valid_in(RMUX_T0_WEST_B1_valid_in),
    .valid_out(RMUX_T0_WEST_B1_valid_out),
    .S(RMUX_T0_WEST_B1_sel_value_O),
    .out_sel(RMUX_T0_WEST_B1_out_sel)
);
SliceWrapper_32_31_32 RMUX_T0_WEST_B1_sel_value (
    .I(config_reg_1_O),
    .O(RMUX_T0_WEST_B1_sel_value_O)
);
wire [0:0] RMUX_T1_EAST_B1_I [1:0];
assign RMUX_T1_EAST_B1_I[1] = REG_T1_EAST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T1_EAST_B1_I[0] = MUX_SB_T1_EAST_SB_OUT_B1_O;
wire [1:0] RMUX_T1_EAST_B1_valid_in;
assign RMUX_T1_EAST_B1_valid_in = {REG_T1_EAST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T1_EAST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T1_EAST_B1 (
    .I(RMUX_T1_EAST_B1_I),
    .O(RMUX_T1_EAST_B1_O),
    .ready_in(SB_T1_EAST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T1_EAST_B1_ready_out),
    .valid_in(RMUX_T1_EAST_B1_valid_in),
    .valid_out(RMUX_T1_EAST_B1_valid_out),
    .S(RMUX_T1_EAST_B1_sel_value_O),
    .out_sel(RMUX_T1_EAST_B1_out_sel)
);
SliceWrapper_32_0_1 RMUX_T1_EAST_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T1_EAST_B1_sel_value_O)
);
wire [0:0] RMUX_T1_NORTH_B1_I [1:0];
assign RMUX_T1_NORTH_B1_I[1] = REG_T1_NORTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T1_NORTH_B1_I[0] = MUX_SB_T1_NORTH_SB_OUT_B1_O;
wire [1:0] RMUX_T1_NORTH_B1_valid_in;
assign RMUX_T1_NORTH_B1_valid_in = {REG_T1_NORTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T1_NORTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T1_NORTH_B1 (
    .I(RMUX_T1_NORTH_B1_I),
    .O(RMUX_T1_NORTH_B1_O),
    .ready_in(SB_T1_NORTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T1_NORTH_B1_ready_out),
    .valid_in(RMUX_T1_NORTH_B1_valid_in),
    .valid_out(RMUX_T1_NORTH_B1_valid_out),
    .S(RMUX_T1_NORTH_B1_sel_value_O),
    .out_sel(RMUX_T1_NORTH_B1_out_sel)
);
SliceWrapper_32_1_2 RMUX_T1_NORTH_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T1_NORTH_B1_sel_value_O)
);
wire [0:0] RMUX_T1_SOUTH_B1_I [1:0];
assign RMUX_T1_SOUTH_B1_I[1] = REG_T1_SOUTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T1_SOUTH_B1_I[0] = MUX_SB_T1_SOUTH_SB_OUT_B1_O;
wire [1:0] RMUX_T1_SOUTH_B1_valid_in;
assign RMUX_T1_SOUTH_B1_valid_in = {REG_T1_SOUTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T1_SOUTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T1_SOUTH_B1 (
    .I(RMUX_T1_SOUTH_B1_I),
    .O(RMUX_T1_SOUTH_B1_O),
    .ready_in(SB_T1_SOUTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T1_SOUTH_B1_ready_out),
    .valid_in(RMUX_T1_SOUTH_B1_valid_in),
    .valid_out(RMUX_T1_SOUTH_B1_valid_out),
    .S(RMUX_T1_SOUTH_B1_sel_value_O),
    .out_sel(RMUX_T1_SOUTH_B1_out_sel)
);
SliceWrapper_32_2_3 RMUX_T1_SOUTH_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T1_SOUTH_B1_sel_value_O)
);
wire [0:0] RMUX_T1_WEST_B1_I [1:0];
assign RMUX_T1_WEST_B1_I[1] = REG_T1_WEST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T1_WEST_B1_I[0] = MUX_SB_T1_WEST_SB_OUT_B1_O;
wire [1:0] RMUX_T1_WEST_B1_valid_in;
assign RMUX_T1_WEST_B1_valid_in = {REG_T1_WEST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T1_WEST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T1_WEST_B1 (
    .I(RMUX_T1_WEST_B1_I),
    .O(RMUX_T1_WEST_B1_O),
    .ready_in(SB_T1_WEST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T1_WEST_B1_ready_out),
    .valid_in(RMUX_T1_WEST_B1_valid_in),
    .valid_out(RMUX_T1_WEST_B1_valid_out),
    .S(RMUX_T1_WEST_B1_sel_value_O),
    .out_sel(RMUX_T1_WEST_B1_out_sel)
);
SliceWrapper_32_3_4 RMUX_T1_WEST_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T1_WEST_B1_sel_value_O)
);
wire [0:0] RMUX_T2_EAST_B1_I [1:0];
assign RMUX_T2_EAST_B1_I[1] = REG_T2_EAST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T2_EAST_B1_I[0] = MUX_SB_T2_EAST_SB_OUT_B1_O;
wire [1:0] RMUX_T2_EAST_B1_valid_in;
assign RMUX_T2_EAST_B1_valid_in = {REG_T2_EAST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T2_EAST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T2_EAST_B1 (
    .I(RMUX_T2_EAST_B1_I),
    .O(RMUX_T2_EAST_B1_O),
    .ready_in(SB_T2_EAST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T2_EAST_B1_ready_out),
    .valid_in(RMUX_T2_EAST_B1_valid_in),
    .valid_out(RMUX_T2_EAST_B1_valid_out),
    .S(RMUX_T2_EAST_B1_sel_value_O),
    .out_sel(RMUX_T2_EAST_B1_out_sel)
);
SliceWrapper_32_4_5 RMUX_T2_EAST_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T2_EAST_B1_sel_value_O)
);
wire [0:0] RMUX_T2_NORTH_B1_I [1:0];
assign RMUX_T2_NORTH_B1_I[1] = REG_T2_NORTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T2_NORTH_B1_I[0] = MUX_SB_T2_NORTH_SB_OUT_B1_O;
wire [1:0] RMUX_T2_NORTH_B1_valid_in;
assign RMUX_T2_NORTH_B1_valid_in = {REG_T2_NORTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T2_NORTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T2_NORTH_B1 (
    .I(RMUX_T2_NORTH_B1_I),
    .O(RMUX_T2_NORTH_B1_O),
    .ready_in(SB_T2_NORTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T2_NORTH_B1_ready_out),
    .valid_in(RMUX_T2_NORTH_B1_valid_in),
    .valid_out(RMUX_T2_NORTH_B1_valid_out),
    .S(RMUX_T2_NORTH_B1_sel_value_O),
    .out_sel(RMUX_T2_NORTH_B1_out_sel)
);
SliceWrapper_32_5_6 RMUX_T2_NORTH_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T2_NORTH_B1_sel_value_O)
);
wire [0:0] RMUX_T2_SOUTH_B1_I [1:0];
assign RMUX_T2_SOUTH_B1_I[1] = REG_T2_SOUTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T2_SOUTH_B1_I[0] = MUX_SB_T2_SOUTH_SB_OUT_B1_O;
wire [1:0] RMUX_T2_SOUTH_B1_valid_in;
assign RMUX_T2_SOUTH_B1_valid_in = {REG_T2_SOUTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T2_SOUTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T2_SOUTH_B1 (
    .I(RMUX_T2_SOUTH_B1_I),
    .O(RMUX_T2_SOUTH_B1_O),
    .ready_in(SB_T2_SOUTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T2_SOUTH_B1_ready_out),
    .valid_in(RMUX_T2_SOUTH_B1_valid_in),
    .valid_out(RMUX_T2_SOUTH_B1_valid_out),
    .S(RMUX_T2_SOUTH_B1_sel_value_O),
    .out_sel(RMUX_T2_SOUTH_B1_out_sel)
);
SliceWrapper_32_6_7 RMUX_T2_SOUTH_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T2_SOUTH_B1_sel_value_O)
);
wire [0:0] RMUX_T2_WEST_B1_I [1:0];
assign RMUX_T2_WEST_B1_I[1] = REG_T2_WEST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T2_WEST_B1_I[0] = MUX_SB_T2_WEST_SB_OUT_B1_O;
wire [1:0] RMUX_T2_WEST_B1_valid_in;
assign RMUX_T2_WEST_B1_valid_in = {REG_T2_WEST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T2_WEST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T2_WEST_B1 (
    .I(RMUX_T2_WEST_B1_I),
    .O(RMUX_T2_WEST_B1_O),
    .ready_in(SB_T2_WEST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T2_WEST_B1_ready_out),
    .valid_in(RMUX_T2_WEST_B1_valid_in),
    .valid_out(RMUX_T2_WEST_B1_valid_out),
    .S(RMUX_T2_WEST_B1_sel_value_O),
    .out_sel(RMUX_T2_WEST_B1_out_sel)
);
SliceWrapper_32_7_8 RMUX_T2_WEST_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T2_WEST_B1_sel_value_O)
);
wire [0:0] RMUX_T3_EAST_B1_I [1:0];
assign RMUX_T3_EAST_B1_I[1] = REG_T3_EAST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T3_EAST_B1_I[0] = MUX_SB_T3_EAST_SB_OUT_B1_O;
wire [1:0] RMUX_T3_EAST_B1_valid_in;
assign RMUX_T3_EAST_B1_valid_in = {REG_T3_EAST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T3_EAST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T3_EAST_B1 (
    .I(RMUX_T3_EAST_B1_I),
    .O(RMUX_T3_EAST_B1_O),
    .ready_in(SB_T3_EAST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T3_EAST_B1_ready_out),
    .valid_in(RMUX_T3_EAST_B1_valid_in),
    .valid_out(RMUX_T3_EAST_B1_valid_out),
    .S(RMUX_T3_EAST_B1_sel_value_O),
    .out_sel(RMUX_T3_EAST_B1_out_sel)
);
SliceWrapper_32_8_9 RMUX_T3_EAST_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T3_EAST_B1_sel_value_O)
);
wire [0:0] RMUX_T3_NORTH_B1_I [1:0];
assign RMUX_T3_NORTH_B1_I[1] = REG_T3_NORTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T3_NORTH_B1_I[0] = MUX_SB_T3_NORTH_SB_OUT_B1_O;
wire [1:0] RMUX_T3_NORTH_B1_valid_in;
assign RMUX_T3_NORTH_B1_valid_in = {REG_T3_NORTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T3_NORTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T3_NORTH_B1 (
    .I(RMUX_T3_NORTH_B1_I),
    .O(RMUX_T3_NORTH_B1_O),
    .ready_in(SB_T3_NORTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T3_NORTH_B1_ready_out),
    .valid_in(RMUX_T3_NORTH_B1_valid_in),
    .valid_out(RMUX_T3_NORTH_B1_valid_out),
    .S(RMUX_T3_NORTH_B1_sel_value_O),
    .out_sel(RMUX_T3_NORTH_B1_out_sel)
);
SliceWrapper_32_9_10 RMUX_T3_NORTH_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T3_NORTH_B1_sel_value_O)
);
wire [0:0] RMUX_T3_SOUTH_B1_I [1:0];
assign RMUX_T3_SOUTH_B1_I[1] = REG_T3_SOUTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T3_SOUTH_B1_I[0] = MUX_SB_T3_SOUTH_SB_OUT_B1_O;
wire [1:0] RMUX_T3_SOUTH_B1_valid_in;
assign RMUX_T3_SOUTH_B1_valid_in = {REG_T3_SOUTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T3_SOUTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T3_SOUTH_B1 (
    .I(RMUX_T3_SOUTH_B1_I),
    .O(RMUX_T3_SOUTH_B1_O),
    .ready_in(SB_T3_SOUTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T3_SOUTH_B1_ready_out),
    .valid_in(RMUX_T3_SOUTH_B1_valid_in),
    .valid_out(RMUX_T3_SOUTH_B1_valid_out),
    .S(RMUX_T3_SOUTH_B1_sel_value_O),
    .out_sel(RMUX_T3_SOUTH_B1_out_sel)
);
SliceWrapper_32_10_11 RMUX_T3_SOUTH_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T3_SOUTH_B1_sel_value_O)
);
wire [0:0] RMUX_T3_WEST_B1_I [1:0];
assign RMUX_T3_WEST_B1_I[1] = REG_T3_WEST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T3_WEST_B1_I[0] = MUX_SB_T3_WEST_SB_OUT_B1_O;
wire [1:0] RMUX_T3_WEST_B1_valid_in;
assign RMUX_T3_WEST_B1_valid_in = {REG_T3_WEST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T3_WEST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T3_WEST_B1 (
    .I(RMUX_T3_WEST_B1_I),
    .O(RMUX_T3_WEST_B1_O),
    .ready_in(SB_T3_WEST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T3_WEST_B1_ready_out),
    .valid_in(RMUX_T3_WEST_B1_valid_in),
    .valid_out(RMUX_T3_WEST_B1_valid_out),
    .S(RMUX_T3_WEST_B1_sel_value_O),
    .out_sel(RMUX_T3_WEST_B1_out_sel)
);
SliceWrapper_32_11_12 RMUX_T3_WEST_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T3_WEST_B1_sel_value_O)
);
wire [0:0] RMUX_T4_EAST_B1_I [1:0];
assign RMUX_T4_EAST_B1_I[1] = REG_T4_EAST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T4_EAST_B1_I[0] = MUX_SB_T4_EAST_SB_OUT_B1_O;
wire [1:0] RMUX_T4_EAST_B1_valid_in;
assign RMUX_T4_EAST_B1_valid_in = {REG_T4_EAST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T4_EAST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T4_EAST_B1 (
    .I(RMUX_T4_EAST_B1_I),
    .O(RMUX_T4_EAST_B1_O),
    .ready_in(SB_T4_EAST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T4_EAST_B1_ready_out),
    .valid_in(RMUX_T4_EAST_B1_valid_in),
    .valid_out(RMUX_T4_EAST_B1_valid_out),
    .S(RMUX_T4_EAST_B1_sel_value_O),
    .out_sel(RMUX_T4_EAST_B1_out_sel)
);
SliceWrapper_32_12_13 RMUX_T4_EAST_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T4_EAST_B1_sel_value_O)
);
wire [0:0] RMUX_T4_NORTH_B1_I [1:0];
assign RMUX_T4_NORTH_B1_I[1] = REG_T4_NORTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T4_NORTH_B1_I[0] = MUX_SB_T4_NORTH_SB_OUT_B1_O;
wire [1:0] RMUX_T4_NORTH_B1_valid_in;
assign RMUX_T4_NORTH_B1_valid_in = {REG_T4_NORTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T4_NORTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T4_NORTH_B1 (
    .I(RMUX_T4_NORTH_B1_I),
    .O(RMUX_T4_NORTH_B1_O),
    .ready_in(SB_T4_NORTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T4_NORTH_B1_ready_out),
    .valid_in(RMUX_T4_NORTH_B1_valid_in),
    .valid_out(RMUX_T4_NORTH_B1_valid_out),
    .S(RMUX_T4_NORTH_B1_sel_value_O),
    .out_sel(RMUX_T4_NORTH_B1_out_sel)
);
SliceWrapper_32_13_14 RMUX_T4_NORTH_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T4_NORTH_B1_sel_value_O)
);
wire [0:0] RMUX_T4_SOUTH_B1_I [1:0];
assign RMUX_T4_SOUTH_B1_I[1] = REG_T4_SOUTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T4_SOUTH_B1_I[0] = MUX_SB_T4_SOUTH_SB_OUT_B1_O;
wire [1:0] RMUX_T4_SOUTH_B1_valid_in;
assign RMUX_T4_SOUTH_B1_valid_in = {REG_T4_SOUTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T4_SOUTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T4_SOUTH_B1 (
    .I(RMUX_T4_SOUTH_B1_I),
    .O(RMUX_T4_SOUTH_B1_O),
    .ready_in(SB_T4_SOUTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T4_SOUTH_B1_ready_out),
    .valid_in(RMUX_T4_SOUTH_B1_valid_in),
    .valid_out(RMUX_T4_SOUTH_B1_valid_out),
    .S(RMUX_T4_SOUTH_B1_sel_value_O),
    .out_sel(RMUX_T4_SOUTH_B1_out_sel)
);
SliceWrapper_32_14_15 RMUX_T4_SOUTH_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T4_SOUTH_B1_sel_value_O)
);
wire [0:0] RMUX_T4_WEST_B1_I [1:0];
assign RMUX_T4_WEST_B1_I[1] = REG_T4_WEST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T4_WEST_B1_I[0] = MUX_SB_T4_WEST_SB_OUT_B1_O;
wire [1:0] RMUX_T4_WEST_B1_valid_in;
assign RMUX_T4_WEST_B1_valid_in = {REG_T4_WEST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T4_WEST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T4_WEST_B1 (
    .I(RMUX_T4_WEST_B1_I),
    .O(RMUX_T4_WEST_B1_O),
    .ready_in(SB_T4_WEST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T4_WEST_B1_ready_out),
    .valid_in(RMUX_T4_WEST_B1_valid_in),
    .valid_out(RMUX_T4_WEST_B1_valid_out),
    .S(RMUX_T4_WEST_B1_sel_value_O),
    .out_sel(RMUX_T4_WEST_B1_out_sel)
);
SliceWrapper_32_15_16 RMUX_T4_WEST_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T4_WEST_B1_sel_value_O)
);
SliceWrapper_32_16_17 SB_T0_EAST_SB_IN_B1_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_EAST_SB_IN_B1_enable_value_O)
);
FanoutHash_302974B49BE3F0C4 SB_T0_EAST_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T0_WEST_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T0_EAST_SB_IN_B1_fan_in_O),
    .E1(SB_T3_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T0_EAST_SB_OUT_B1_FANOUT_I;
assign SB_T0_EAST_SB_OUT_B1_FANOUT_I = {REG_T0_EAST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T0_EAST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T0_EAST_SB_OUT_B1_FANOUT (
    .S(RMUX_T0_EAST_B1_out_sel),
    .O(SB_T0_EAST_SB_OUT_B1_FANOUT_O),
    .I(SB_T0_EAST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_32_17_18 SB_T0_EAST_SB_OUT_B1_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_EAST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_32_18_21 SB_T0_EAST_SB_OUT_B1_sel_value (
    .I(config_reg_2_O),
    .O(SB_T0_EAST_SB_OUT_B1_sel_value_O)
);
SliceWrapper_32_21_22 SB_T0_NORTH_SB_IN_B1_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_NORTH_SB_IN_B1_enable_value_O)
);
FanoutHash_47712AAC902ADA2 SB_T0_NORTH_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T0_WEST_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T0_NORTH_SB_IN_B1_fan_in_O),
    .E1(SB_T1_EAST_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T0_NORTH_SB_OUT_B1_FANOUT_I;
assign SB_T0_NORTH_SB_OUT_B1_FANOUT_I = {REG_T0_NORTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T0_NORTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T0_NORTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T0_NORTH_B1_out_sel),
    .O(SB_T0_NORTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T0_NORTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_32_22_23 SB_T0_NORTH_SB_OUT_B1_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_NORTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_32_23_26 SB_T0_NORTH_SB_OUT_B1_sel_value (
    .I(config_reg_2_O),
    .O(SB_T0_NORTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_32_26_27 SB_T0_SOUTH_SB_IN_B1_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_SOUTH_SB_IN_B1_enable_value_O)
);
FanoutHash_2785CE916183C5C SB_T0_SOUTH_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T1_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T3_EAST_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T0_SOUTH_SB_IN_B1_fan_in_O),
    .E1(SB_T0_NORTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T0_SOUTH_SB_OUT_B1_FANOUT_I;
assign SB_T0_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T0_SOUTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T0_SOUTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T0_SOUTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T0_SOUTH_B1_out_sel),
    .O(SB_T0_SOUTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T0_SOUTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_32_27_28 SB_T0_SOUTH_SB_OUT_B1_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_SOUTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_32_28_31 SB_T0_SOUTH_SB_OUT_B1_sel_value (
    .I(config_reg_2_O),
    .O(SB_T0_SOUTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_32_31_32 SB_T0_WEST_SB_IN_B1_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_WEST_SB_IN_B1_enable_value_O)
);
FanoutHash_65A468071775C7BB SB_T0_WEST_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T0_EAST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T0_WEST_SB_IN_B1_fan_in_O),
    .E1(SB_T4_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T0_WEST_SB_OUT_B1_FANOUT_I;
assign SB_T0_WEST_SB_OUT_B1_FANOUT_I = {REG_T0_WEST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T0_WEST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T0_WEST_SB_OUT_B1_FANOUT (
    .S(RMUX_T0_WEST_B1_out_sel),
    .O(SB_T0_WEST_SB_OUT_B1_FANOUT_O),
    .I(SB_T0_WEST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_31_0_1 SB_T0_WEST_SB_OUT_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T0_WEST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_31_1_4 SB_T0_WEST_SB_OUT_B1_sel_value (
    .I(config_reg_3_O),
    .O(SB_T0_WEST_SB_OUT_B1_sel_value_O)
);
SliceWrapper_31_4_5 SB_T1_EAST_SB_IN_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_EAST_SB_IN_B1_enable_value_O)
);
FanoutHash_4F83851A40824F89 SB_T1_EAST_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T1_EAST_SB_IN_B1_fan_in_O),
    .E1(SB_T1_WEST_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T1_EAST_SB_OUT_B1_FANOUT_I;
assign SB_T1_EAST_SB_OUT_B1_FANOUT_I = {REG_T1_EAST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T1_EAST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T1_EAST_SB_OUT_B1_FANOUT (
    .S(RMUX_T1_EAST_B1_out_sel),
    .O(SB_T1_EAST_SB_OUT_B1_FANOUT_O),
    .I(SB_T1_EAST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_31_5_6 SB_T1_EAST_SB_OUT_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_EAST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_31_6_9 SB_T1_EAST_SB_OUT_B1_sel_value (
    .I(config_reg_3_O),
    .O(SB_T1_EAST_SB_OUT_B1_sel_value_O)
);
SliceWrapper_31_9_10 SB_T1_NORTH_SB_IN_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_NORTH_SB_IN_B1_enable_value_O)
);
FanoutHash_4FADDC8F90390680 SB_T1_NORTH_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T4_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T2_EAST_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T1_NORTH_SB_IN_B1_fan_in_O),
    .E1(SB_T1_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T1_NORTH_SB_OUT_B1_FANOUT_I;
assign SB_T1_NORTH_SB_OUT_B1_FANOUT_I = {REG_T1_NORTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T1_NORTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T1_NORTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T1_NORTH_B1_out_sel),
    .O(SB_T1_NORTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T1_NORTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_31_10_11 SB_T1_NORTH_SB_OUT_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_NORTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_31_11_14 SB_T1_NORTH_SB_OUT_B1_sel_value (
    .I(config_reg_3_O),
    .O(SB_T1_NORTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_31_14_15 SB_T1_SOUTH_SB_IN_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_SOUTH_SB_IN_B1_enable_value_O)
);
FanoutHash_466EB88CFD0CAD7B SB_T1_SOUTH_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T2_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T2_EAST_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T1_SOUTH_SB_IN_B1_fan_in_O),
    .E1(SB_T1_NORTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T1_SOUTH_SB_OUT_B1_FANOUT_I;
assign SB_T1_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T1_SOUTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T1_SOUTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T1_SOUTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T1_SOUTH_B1_out_sel),
    .O(SB_T1_SOUTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T1_SOUTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_31_15_16 SB_T1_SOUTH_SB_OUT_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_SOUTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_31_16_19 SB_T1_SOUTH_SB_OUT_B1_sel_value (
    .I(config_reg_3_O),
    .O(SB_T1_SOUTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_31_19_20 SB_T1_WEST_SB_IN_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_WEST_SB_IN_B1_enable_value_O)
);
FanoutHash_7ED1C80229B84786 SB_T1_WEST_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T1_EAST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T1_WEST_SB_IN_B1_fan_in_O),
    .E1(SB_T0_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T1_WEST_SB_OUT_B1_FANOUT_I;
assign SB_T1_WEST_SB_OUT_B1_FANOUT_I = {REG_T1_WEST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T1_WEST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T1_WEST_SB_OUT_B1_FANOUT (
    .S(RMUX_T1_WEST_B1_out_sel),
    .O(SB_T1_WEST_SB_OUT_B1_FANOUT_O),
    .I(SB_T1_WEST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_31_20_21 SB_T1_WEST_SB_OUT_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_WEST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_31_21_24 SB_T1_WEST_SB_OUT_B1_sel_value (
    .I(config_reg_3_O),
    .O(SB_T1_WEST_SB_OUT_B1_sel_value_O)
);
SliceWrapper_31_24_25 SB_T2_EAST_SB_IN_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T2_EAST_SB_IN_B1_enable_value_O)
);
FanoutHash_7F4660D1463D9234 SB_T2_EAST_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T2_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T2_EAST_SB_IN_B1_fan_in_O),
    .E1(SB_T1_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T2_EAST_SB_OUT_B1_FANOUT_I;
assign SB_T2_EAST_SB_OUT_B1_FANOUT_I = {REG_T2_EAST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T2_EAST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T2_EAST_SB_OUT_B1_FANOUT (
    .S(RMUX_T2_EAST_B1_out_sel),
    .O(SB_T2_EAST_SB_OUT_B1_FANOUT_O),
    .I(SB_T2_EAST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_31_25_26 SB_T2_EAST_SB_OUT_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T2_EAST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_31_26_29 SB_T2_EAST_SB_OUT_B1_sel_value (
    .I(config_reg_3_O),
    .O(SB_T2_EAST_SB_OUT_B1_sel_value_O)
);
SliceWrapper_31_29_30 SB_T2_NORTH_SB_IN_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T2_NORTH_SB_IN_B1_enable_value_O)
);
FanoutHash_3B67229CB02928BA SB_T2_NORTH_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T3_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T3_EAST_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T2_NORTH_SB_IN_B1_fan_in_O),
    .E1(SB_T2_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T2_NORTH_SB_OUT_B1_FANOUT_I;
assign SB_T2_NORTH_SB_OUT_B1_FANOUT_I = {REG_T2_NORTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T2_NORTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T2_NORTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T2_NORTH_B1_out_sel),
    .O(SB_T2_NORTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T2_NORTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_31_30_31 SB_T2_NORTH_SB_OUT_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T2_NORTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_30_0_3 SB_T2_NORTH_SB_OUT_B1_sel_value (
    .I(config_reg_4_O),
    .O(SB_T2_NORTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_30_3_4 SB_T2_SOUTH_SB_IN_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T2_SOUTH_SB_IN_B1_enable_value_O)
);
FanoutHash_28125A548B305607 SB_T2_SOUTH_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T3_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T1_EAST_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T2_SOUTH_SB_IN_B1_fan_in_O),
    .E1(SB_T2_NORTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T2_SOUTH_SB_OUT_B1_FANOUT_I;
assign SB_T2_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T2_SOUTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T2_SOUTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T2_SOUTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T2_SOUTH_B1_out_sel),
    .O(SB_T2_SOUTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T2_SOUTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_30_4_5 SB_T2_SOUTH_SB_OUT_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T2_SOUTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_30_5_8 SB_T2_SOUTH_SB_OUT_B1_sel_value (
    .I(config_reg_4_O),
    .O(SB_T2_SOUTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_30_8_9 SB_T2_WEST_SB_IN_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T2_WEST_SB_IN_B1_enable_value_O)
);
FanoutHash_752C11B748DD905C SB_T2_WEST_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T2_EAST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T2_WEST_SB_IN_B1_fan_in_O),
    .E1(SB_T1_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T2_WEST_SB_OUT_B1_FANOUT_I;
assign SB_T2_WEST_SB_OUT_B1_FANOUT_I = {REG_T2_WEST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T2_WEST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T2_WEST_SB_OUT_B1_FANOUT (
    .S(RMUX_T2_WEST_B1_out_sel),
    .O(SB_T2_WEST_SB_OUT_B1_FANOUT_O),
    .I(SB_T2_WEST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_30_9_10 SB_T2_WEST_SB_OUT_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T2_WEST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_30_10_13 SB_T2_WEST_SB_OUT_B1_sel_value (
    .I(config_reg_4_O),
    .O(SB_T2_WEST_SB_OUT_B1_sel_value_O)
);
SliceWrapper_30_13_14 SB_T3_EAST_SB_IN_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_EAST_SB_IN_B1_enable_value_O)
);
FanoutHash_43D5C80ABD816837 SB_T3_EAST_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T3_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T3_EAST_SB_IN_B1_fan_in_O),
    .E1(SB_T2_NORTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T3_EAST_SB_OUT_B1_FANOUT_I;
assign SB_T3_EAST_SB_OUT_B1_FANOUT_I = {REG_T3_EAST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T3_EAST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T3_EAST_SB_OUT_B1_FANOUT (
    .S(RMUX_T3_EAST_B1_out_sel),
    .O(SB_T3_EAST_SB_OUT_B1_FANOUT_O),
    .I(SB_T3_EAST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_30_14_15 SB_T3_EAST_SB_OUT_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_EAST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_30_15_18 SB_T3_EAST_SB_OUT_B1_sel_value (
    .I(config_reg_4_O),
    .O(SB_T3_EAST_SB_OUT_B1_sel_value_O)
);
SliceWrapper_30_18_19 SB_T3_NORTH_SB_IN_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_NORTH_SB_IN_B1_enable_value_O)
);
FanoutHash_69376833A2418E2 SB_T3_NORTH_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T2_WEST_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T3_NORTH_SB_IN_B1_fan_in_O),
    .E1(SB_T4_EAST_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T3_NORTH_SB_OUT_B1_FANOUT_I;
assign SB_T3_NORTH_SB_OUT_B1_FANOUT_I = {REG_T3_NORTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T3_NORTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T3_NORTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T3_NORTH_B1_out_sel),
    .O(SB_T3_NORTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T3_NORTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_30_19_20 SB_T3_NORTH_SB_OUT_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_NORTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_30_20_23 SB_T3_NORTH_SB_OUT_B1_sel_value (
    .I(config_reg_4_O),
    .O(SB_T3_NORTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_30_23_24 SB_T3_SOUTH_SB_IN_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_SOUTH_SB_IN_B1_enable_value_O)
);
FanoutHash_66A75CC8494A4D6B SB_T3_SOUTH_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T4_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T0_EAST_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T3_SOUTH_SB_IN_B1_fan_in_O),
    .E1(SB_T3_NORTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T3_SOUTH_SB_OUT_B1_FANOUT_I;
assign SB_T3_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T3_SOUTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T3_SOUTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T3_SOUTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T3_SOUTH_B1_out_sel),
    .O(SB_T3_SOUTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T3_SOUTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_30_24_25 SB_T3_SOUTH_SB_OUT_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_SOUTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_30_25_28 SB_T3_SOUTH_SB_OUT_B1_sel_value (
    .I(config_reg_4_O),
    .O(SB_T3_SOUTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_30_28_29 SB_T3_WEST_SB_IN_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_WEST_SB_IN_B1_enable_value_O)
);
FanoutHash_31AE65CCDD94603 SB_T3_WEST_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T3_EAST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T3_WEST_SB_IN_B1_fan_in_O),
    .E1(SB_T2_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T3_WEST_SB_OUT_B1_FANOUT_I;
assign SB_T3_WEST_SB_OUT_B1_FANOUT_I = {REG_T3_WEST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T3_WEST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T3_WEST_SB_OUT_B1_FANOUT (
    .S(RMUX_T3_WEST_B1_out_sel),
    .O(SB_T3_WEST_SB_OUT_B1_FANOUT_O),
    .I(SB_T3_WEST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_30_29_30 SB_T3_WEST_SB_OUT_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_WEST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_23_0_3 SB_T3_WEST_SB_OUT_B1_sel_value (
    .I(config_reg_5_O),
    .O(SB_T3_WEST_SB_OUT_B1_sel_value_O)
);
SliceWrapper_23_3_4 SB_T4_EAST_SB_IN_B1_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_EAST_SB_IN_B1_enable_value_O)
);
FanoutHash_5D7AEC1255CDC1CC SB_T4_EAST_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T4_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T4_EAST_SB_IN_B1_fan_in_O),
    .E1(SB_T4_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T4_EAST_SB_OUT_B1_FANOUT_I;
assign SB_T4_EAST_SB_OUT_B1_FANOUT_I = {REG_T4_EAST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T4_EAST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T4_EAST_SB_OUT_B1_FANOUT (
    .S(RMUX_T4_EAST_B1_out_sel),
    .O(SB_T4_EAST_SB_OUT_B1_FANOUT_O),
    .I(SB_T4_EAST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_23_4_5 SB_T4_EAST_SB_OUT_B1_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_EAST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_23_5_8 SB_T4_EAST_SB_OUT_B1_sel_value (
    .I(config_reg_5_O),
    .O(SB_T4_EAST_SB_OUT_B1_sel_value_O)
);
SliceWrapper_23_8_9 SB_T4_NORTH_SB_IN_B1_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_NORTH_SB_IN_B1_enable_value_O)
);
FanoutHash_184DFC10DAF19BE9 SB_T4_NORTH_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T1_WEST_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T4_NORTH_SB_IN_B1_fan_in_O),
    .E1(SB_T0_EAST_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T4_NORTH_SB_OUT_B1_FANOUT_I;
assign SB_T4_NORTH_SB_OUT_B1_FANOUT_I = {REG_T4_NORTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T4_NORTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T4_NORTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T4_NORTH_B1_out_sel),
    .O(SB_T4_NORTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T4_NORTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_23_9_10 SB_T4_NORTH_SB_OUT_B1_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_NORTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_23_10_13 SB_T4_NORTH_SB_OUT_B1_sel_value (
    .I(config_reg_5_O),
    .O(SB_T4_NORTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_23_13_14 SB_T4_SOUTH_SB_IN_B1_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_SOUTH_SB_IN_B1_enable_value_O)
);
FanoutHash_26B6474864379B6A SB_T4_SOUTH_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T0_WEST_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T4_SOUTH_SB_IN_B1_fan_in_O),
    .E1(SB_T4_EAST_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T4_SOUTH_SB_OUT_B1_FANOUT_I;
assign SB_T4_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T4_SOUTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T4_SOUTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T4_SOUTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T4_SOUTH_B1_out_sel),
    .O(SB_T4_SOUTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T4_SOUTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_23_14_15 SB_T4_SOUTH_SB_OUT_B1_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_SOUTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_23_15_18 SB_T4_SOUTH_SB_OUT_B1_sel_value (
    .I(config_reg_5_O),
    .O(SB_T4_SOUTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_23_18_19 SB_T4_WEST_SB_IN_B1_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_WEST_SB_IN_B1_enable_value_O)
);
FanoutHash_1816466D6957000 SB_T4_WEST_SB_IN_B1_fan_in (
    .S6(const_0_32_out),
    .E2(SB_T4_EAST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
    .I3(PE_input_width_1_num_0_ready),
    .S0(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
    .E5(PE_input_width_1_num_2_enable),
    .I6(const_0_1_out),
    .I2(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
    .S3(PE_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
    .E3(PE_input_width_1_num_0_enable),
    .E0(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
    .S4(PE_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
    .E4(PE_input_width_1_num_1_enable),
    .S5(PE_input_width_1_num_2_out_sel),
    .I1(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
    .I5(PE_input_width_1_num_2_ready),
    .E6(const_0_1_out),
    .I4(PE_input_width_1_num_1_ready),
    .O(SB_T4_WEST_SB_IN_B1_fan_in_O),
    .E1(SB_T3_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T4_WEST_SB_OUT_B1_FANOUT_I;
assign SB_T4_WEST_SB_OUT_B1_FANOUT_I = {REG_T4_WEST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T4_WEST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T4_WEST_SB_OUT_B1_FANOUT (
    .S(RMUX_T4_WEST_B1_out_sel),
    .O(SB_T4_WEST_SB_OUT_B1_FANOUT_O),
    .I(SB_T4_WEST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_23_19_20 SB_T4_WEST_SB_OUT_B1_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_WEST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_23_20_23 SB_T4_WEST_SB_OUT_B1_sel_value (
    .I(config_reg_5_O),
    .O(SB_T4_WEST_SB_OUT_B1_sel_value_O)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T0_EAST_SB_IN_B1 (
    .I(SB_T0_EAST_SB_IN_B1),
    .O(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .ready_in(SB_T0_EAST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T0_EAST_SB_IN_B1_ready_out),
    .valid_in(SB_T0_EAST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T0_EAST_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T0_NORTH_SB_IN_B1 (
    .I(SB_T0_NORTH_SB_IN_B1),
    .O(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .ready_in(SB_T0_NORTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T0_NORTH_SB_IN_B1_ready_out),
    .valid_in(SB_T0_NORTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T0_NORTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T0_SOUTH_SB_IN_B1 (
    .I(SB_T0_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .ready_in(SB_T0_SOUTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T0_SOUTH_SB_IN_B1_ready_out),
    .valid_in(SB_T0_SOUTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T0_WEST_SB_IN_B1 (
    .I(SB_T0_WEST_SB_IN_B1),
    .O(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .ready_in(SB_T0_WEST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T0_WEST_SB_IN_B1_ready_out),
    .valid_in(SB_T0_WEST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T0_WEST_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T1_EAST_SB_IN_B1 (
    .I(SB_T1_EAST_SB_IN_B1),
    .O(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .ready_in(SB_T1_EAST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T1_EAST_SB_IN_B1_ready_out),
    .valid_in(SB_T1_EAST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T1_EAST_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T1_NORTH_SB_IN_B1 (
    .I(SB_T1_NORTH_SB_IN_B1),
    .O(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .ready_in(SB_T1_NORTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T1_NORTH_SB_IN_B1_ready_out),
    .valid_in(SB_T1_NORTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T1_NORTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T1_SOUTH_SB_IN_B1 (
    .I(SB_T1_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .ready_in(SB_T1_SOUTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T1_SOUTH_SB_IN_B1_ready_out),
    .valid_in(SB_T1_SOUTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T1_WEST_SB_IN_B1 (
    .I(SB_T1_WEST_SB_IN_B1),
    .O(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .ready_in(SB_T1_WEST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T1_WEST_SB_IN_B1_ready_out),
    .valid_in(SB_T1_WEST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T1_WEST_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T2_EAST_SB_IN_B1 (
    .I(SB_T2_EAST_SB_IN_B1),
    .O(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .ready_in(SB_T2_EAST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T2_EAST_SB_IN_B1_ready_out),
    .valid_in(SB_T2_EAST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T2_EAST_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T2_NORTH_SB_IN_B1 (
    .I(SB_T2_NORTH_SB_IN_B1),
    .O(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .ready_in(SB_T2_NORTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T2_NORTH_SB_IN_B1_ready_out),
    .valid_in(SB_T2_NORTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T2_NORTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T2_SOUTH_SB_IN_B1 (
    .I(SB_T2_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .ready_in(SB_T2_SOUTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T2_SOUTH_SB_IN_B1_ready_out),
    .valid_in(SB_T2_SOUTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T2_WEST_SB_IN_B1 (
    .I(SB_T2_WEST_SB_IN_B1),
    .O(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .ready_in(SB_T2_WEST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T2_WEST_SB_IN_B1_ready_out),
    .valid_in(SB_T2_WEST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T2_WEST_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T3_EAST_SB_IN_B1 (
    .I(SB_T3_EAST_SB_IN_B1),
    .O(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .ready_in(SB_T3_EAST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T3_EAST_SB_IN_B1_ready_out),
    .valid_in(SB_T3_EAST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T3_EAST_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T3_NORTH_SB_IN_B1 (
    .I(SB_T3_NORTH_SB_IN_B1),
    .O(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .ready_in(SB_T3_NORTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T3_NORTH_SB_IN_B1_ready_out),
    .valid_in(SB_T3_NORTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T3_NORTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T3_SOUTH_SB_IN_B1 (
    .I(SB_T3_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .ready_in(SB_T3_SOUTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T3_SOUTH_SB_IN_B1_ready_out),
    .valid_in(SB_T3_SOUTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T3_WEST_SB_IN_B1 (
    .I(SB_T3_WEST_SB_IN_B1),
    .O(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .ready_in(SB_T3_WEST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T3_WEST_SB_IN_B1_ready_out),
    .valid_in(SB_T3_WEST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T3_WEST_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T4_EAST_SB_IN_B1 (
    .I(SB_T4_EAST_SB_IN_B1),
    .O(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .ready_in(SB_T4_EAST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T4_EAST_SB_IN_B1_ready_out),
    .valid_in(SB_T4_EAST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T4_EAST_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T4_NORTH_SB_IN_B1 (
    .I(SB_T4_NORTH_SB_IN_B1),
    .O(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .ready_in(SB_T4_NORTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T4_NORTH_SB_IN_B1_ready_out),
    .valid_in(SB_T4_NORTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T4_NORTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T4_SOUTH_SB_IN_B1 (
    .I(SB_T4_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .ready_in(SB_T4_SOUTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T4_SOUTH_SB_IN_B1_ready_out),
    .valid_in(SB_T4_SOUTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T4_WEST_SB_IN_B1 (
    .I(SB_T4_WEST_SB_IN_B1),
    .O(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .ready_in(SB_T4_WEST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T4_WEST_SB_IN_B1_ready_out),
    .valid_in(SB_T4_WEST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T4_WEST_SB_IN_B1_valid_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_23_32_inst0$bit_const_0_None (
    .out(ZextWrapper_23_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_23_32_inst0$self_O_out;
assign ZextWrapper_23_32_inst0$self_O_out = {ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,config_reg_5_O};
mantle_wire__typeBitIn32 ZextWrapper_23_32_inst0$self_O (
    .in(ZextWrapper_23_32_inst0$self_O_in),
    .out(ZextWrapper_23_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_30_32_inst0$bit_const_0_None (
    .out(ZextWrapper_30_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_30_32_inst0$self_O_out;
assign ZextWrapper_30_32_inst0$self_O_out = {ZextWrapper_30_32_inst0$bit_const_0_None_out,ZextWrapper_30_32_inst0$bit_const_0_None_out,config_reg_4_O};
mantle_wire__typeBitIn32 ZextWrapper_30_32_inst0$self_O (
    .in(ZextWrapper_30_32_inst0$self_O_in),
    .out(ZextWrapper_30_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_31_32_inst0$bit_const_0_None (
    .out(ZextWrapper_31_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_31_32_inst0$self_O_out;
assign ZextWrapper_31_32_inst0$self_O_out = {ZextWrapper_31_32_inst0$bit_const_0_None_out,config_reg_3_O};
mantle_wire__typeBitIn32 ZextWrapper_31_32_inst0$self_O (
    .in(ZextWrapper_31_32_inst0$self_O_in),
    .out(ZextWrapper_31_32_inst0$self_O_out)
);
coreir_and #(
    .width(1)
) and1_inst0 (
    .in0(coreir_eq_1_inst0_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst0_out)
);
coreir_and #(
    .width(1)
) and1_inst1 (
    .in0(coreir_eq_1_inst1_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst1_out)
);
coreir_and #(
    .width(1)
) and1_inst10 (
    .in0(coreir_eq_1_inst10_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst10_out)
);
coreir_and #(
    .width(1)
) and1_inst11 (
    .in0(coreir_eq_1_inst11_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst11_out)
);
coreir_and #(
    .width(1)
) and1_inst12 (
    .in0(coreir_eq_1_inst12_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst12_out)
);
coreir_and #(
    .width(1)
) and1_inst13 (
    .in0(coreir_eq_1_inst13_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst13_out)
);
coreir_and #(
    .width(1)
) and1_inst14 (
    .in0(coreir_eq_1_inst14_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst14_out)
);
coreir_and #(
    .width(1)
) and1_inst15 (
    .in0(coreir_eq_1_inst15_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst15_out)
);
coreir_and #(
    .width(1)
) and1_inst16 (
    .in0(coreir_eq_1_inst16_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst16_out)
);
coreir_and #(
    .width(1)
) and1_inst17 (
    .in0(coreir_eq_1_inst17_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst17_out)
);
coreir_and #(
    .width(1)
) and1_inst18 (
    .in0(coreir_eq_1_inst18_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst18_out)
);
coreir_and #(
    .width(1)
) and1_inst19 (
    .in0(coreir_eq_1_inst19_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst19_out)
);
coreir_and #(
    .width(1)
) and1_inst2 (
    .in0(coreir_eq_1_inst2_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst2_out)
);
coreir_and #(
    .width(1)
) and1_inst3 (
    .in0(coreir_eq_1_inst3_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst3_out)
);
coreir_and #(
    .width(1)
) and1_inst4 (
    .in0(coreir_eq_1_inst4_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst4_out)
);
coreir_and #(
    .width(1)
) and1_inst5 (
    .in0(coreir_eq_1_inst5_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst5_out)
);
coreir_and #(
    .width(1)
) and1_inst6 (
    .in0(coreir_eq_1_inst6_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst6_out)
);
coreir_and #(
    .width(1)
) and1_inst7 (
    .in0(coreir_eq_1_inst7_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst7_out)
);
coreir_and #(
    .width(1)
) and1_inst8 (
    .in0(coreir_eq_1_inst8_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst8_out)
);
coreir_and #(
    .width(1)
) and1_inst9 (
    .in0(coreir_eq_1_inst9_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst9_out)
);
wire [7:0] config_reg_0_config_addr;
assign config_reg_0_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_32_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_reg_0_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_1_config_addr;
assign config_reg_1_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_32_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_reg_1_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_2_config_addr;
assign config_reg_2_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_32_8_32_2 config_reg_2 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_2_O),
    .config_addr(config_reg_2_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_3_config_addr;
assign config_reg_3_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_31_8_32_3 config_reg_3 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_3_O),
    .config_addr(config_reg_3_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_4_config_addr;
assign config_reg_4_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_30_8_32_4 config_reg_4 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_4_O),
    .config_addr(config_reg_4_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_5_config_addr;
assign config_reg_5_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_23_8_32_5 config_reg_5 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_5_O),
    .config_addr(config_reg_5_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_const #(
    .value(1'h0),
    .width(1)
) const_0_1 (
    .out(const_0_1_out)
);
coreir_const #(
    .value(32'h00000000),
    .width(32)
) const_0_32 (
    .out(const_0_32_out)
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst0 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_NORTH_B1_sel_value_O),
    .out(coreir_eq_1_inst0_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst1 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_SOUTH_B1_sel_value_O),
    .out(coreir_eq_1_inst1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst10 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_EAST_B1_sel_value_O),
    .out(coreir_eq_1_inst10_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst11 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_WEST_B1_sel_value_O),
    .out(coreir_eq_1_inst11_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst12 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_NORTH_B1_sel_value_O),
    .out(coreir_eq_1_inst12_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst13 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_SOUTH_B1_sel_value_O),
    .out(coreir_eq_1_inst13_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst14 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_EAST_B1_sel_value_O),
    .out(coreir_eq_1_inst14_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst15 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_WEST_B1_sel_value_O),
    .out(coreir_eq_1_inst15_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst16 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_NORTH_B1_sel_value_O),
    .out(coreir_eq_1_inst16_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst17 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_SOUTH_B1_sel_value_O),
    .out(coreir_eq_1_inst17_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst18 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_EAST_B1_sel_value_O),
    .out(coreir_eq_1_inst18_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst19 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_WEST_B1_sel_value_O),
    .out(coreir_eq_1_inst19_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst2 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_EAST_B1_sel_value_O),
    .out(coreir_eq_1_inst2_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst3 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_WEST_B1_sel_value_O),
    .out(coreir_eq_1_inst3_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst4 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_NORTH_B1_sel_value_O),
    .out(coreir_eq_1_inst4_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst5 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_SOUTH_B1_sel_value_O),
    .out(coreir_eq_1_inst5_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst6 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_EAST_B1_sel_value_O),
    .out(coreir_eq_1_inst6_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst7 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_WEST_B1_sel_value_O),
    .out(coreir_eq_1_inst7_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst8 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_NORTH_B1_sel_value_O),
    .out(coreir_eq_1_inst8_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst9 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_SOUTH_B1_sel_value_O),
    .out(coreir_eq_1_inst9_out)
);
wire [31:0] mux_aoi_6_32_inst0_I [5:0];
assign mux_aoi_6_32_inst0_I[5] = ZextWrapper_23_32_inst0$self_O_in;
assign mux_aoi_6_32_inst0_I[4] = ZextWrapper_30_32_inst0$self_O_in;
assign mux_aoi_6_32_inst0_I[3] = ZextWrapper_31_32_inst0$self_O_in;
assign mux_aoi_6_32_inst0_I[2] = config_reg_2_O;
assign mux_aoi_6_32_inst0_I[1] = config_reg_1_O;
assign mux_aoi_6_32_inst0_I[0] = config_reg_0_O;
mux_aoi_6_32 mux_aoi_6_32_inst0 (
    .I(mux_aoi_6_32_inst0_I),
    .O(mux_aoi_6_32_inst0_O),
    .S(self_config_config_addr_out[2:0]),
    .out_sel(mux_aoi_6_32_inst0_out_sel)
);
mantle_wire__typeBit8 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
assign PE_output_width_1_num_0_ready_out = CB_PE_output_width_1_num_0_fan_in_O[0];
assign PondTop_output_width_1_num_0_ready_out = CB_PondTop_output_width_1_num_0_fan_in_O[0];
assign PondTop_output_width_1_num_1_ready_out = CB_PondTop_output_width_1_num_1_fan_in_O[0];
assign SB_T0_EAST_SB_IN_B1_enable = SB_T0_EAST_SB_IN_B1_enable_value_O[0];
assign SB_T0_EAST_SB_IN_B1_ready_out = WIRE_SB_T0_EAST_SB_IN_B1_ready_out;
assign SB_T0_EAST_SB_OUT_B1 = RMUX_T0_EAST_B1_O;
assign SB_T0_EAST_SB_OUT_B1_enable = SB_T0_EAST_SB_OUT_B1_enable_value_O[0];
assign SB_T0_EAST_SB_OUT_B1_valid_out = RMUX_T0_EAST_B1_valid_out;
assign SB_T0_NORTH_SB_IN_B1_enable = SB_T0_NORTH_SB_IN_B1_enable_value_O[0];
assign SB_T0_NORTH_SB_IN_B1_ready_out = WIRE_SB_T0_NORTH_SB_IN_B1_ready_out;
assign SB_T0_NORTH_SB_OUT_B1 = RMUX_T0_NORTH_B1_O;
assign SB_T0_NORTH_SB_OUT_B1_enable = SB_T0_NORTH_SB_OUT_B1_enable_value_O[0];
assign SB_T0_NORTH_SB_OUT_B1_valid_out = RMUX_T0_NORTH_B1_valid_out;
assign SB_T0_SOUTH_SB_IN_B1_enable = SB_T0_SOUTH_SB_IN_B1_enable_value_O[0];
assign SB_T0_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T0_SOUTH_SB_IN_B1_ready_out;
assign SB_T0_SOUTH_SB_OUT_B1 = RMUX_T0_SOUTH_B1_O;
assign SB_T0_SOUTH_SB_OUT_B1_enable = SB_T0_SOUTH_SB_OUT_B1_enable_value_O[0];
assign SB_T0_SOUTH_SB_OUT_B1_valid_out = RMUX_T0_SOUTH_B1_valid_out;
assign SB_T0_WEST_SB_IN_B1_enable = SB_T0_WEST_SB_IN_B1_enable_value_O[0];
assign SB_T0_WEST_SB_IN_B1_ready_out = WIRE_SB_T0_WEST_SB_IN_B1_ready_out;
assign SB_T0_WEST_SB_OUT_B1 = RMUX_T0_WEST_B1_O;
assign SB_T0_WEST_SB_OUT_B1_enable = SB_T0_WEST_SB_OUT_B1_enable_value_O[0];
assign SB_T0_WEST_SB_OUT_B1_valid_out = RMUX_T0_WEST_B1_valid_out;
assign SB_T1_EAST_SB_IN_B1_enable = SB_T1_EAST_SB_IN_B1_enable_value_O[0];
assign SB_T1_EAST_SB_IN_B1_ready_out = WIRE_SB_T1_EAST_SB_IN_B1_ready_out;
assign SB_T1_EAST_SB_OUT_B1 = RMUX_T1_EAST_B1_O;
assign SB_T1_EAST_SB_OUT_B1_enable = SB_T1_EAST_SB_OUT_B1_enable_value_O[0];
assign SB_T1_EAST_SB_OUT_B1_valid_out = RMUX_T1_EAST_B1_valid_out;
assign SB_T1_NORTH_SB_IN_B1_enable = SB_T1_NORTH_SB_IN_B1_enable_value_O[0];
assign SB_T1_NORTH_SB_IN_B1_ready_out = WIRE_SB_T1_NORTH_SB_IN_B1_ready_out;
assign SB_T1_NORTH_SB_OUT_B1 = RMUX_T1_NORTH_B1_O;
assign SB_T1_NORTH_SB_OUT_B1_enable = SB_T1_NORTH_SB_OUT_B1_enable_value_O[0];
assign SB_T1_NORTH_SB_OUT_B1_valid_out = RMUX_T1_NORTH_B1_valid_out;
assign SB_T1_SOUTH_SB_IN_B1_enable = SB_T1_SOUTH_SB_IN_B1_enable_value_O[0];
assign SB_T1_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T1_SOUTH_SB_IN_B1_ready_out;
assign SB_T1_SOUTH_SB_OUT_B1 = RMUX_T1_SOUTH_B1_O;
assign SB_T1_SOUTH_SB_OUT_B1_enable = SB_T1_SOUTH_SB_OUT_B1_enable_value_O[0];
assign SB_T1_SOUTH_SB_OUT_B1_valid_out = RMUX_T1_SOUTH_B1_valid_out;
assign SB_T1_WEST_SB_IN_B1_enable = SB_T1_WEST_SB_IN_B1_enable_value_O[0];
assign SB_T1_WEST_SB_IN_B1_ready_out = WIRE_SB_T1_WEST_SB_IN_B1_ready_out;
assign SB_T1_WEST_SB_OUT_B1 = RMUX_T1_WEST_B1_O;
assign SB_T1_WEST_SB_OUT_B1_enable = SB_T1_WEST_SB_OUT_B1_enable_value_O[0];
assign SB_T1_WEST_SB_OUT_B1_valid_out = RMUX_T1_WEST_B1_valid_out;
assign SB_T2_EAST_SB_IN_B1_enable = SB_T2_EAST_SB_IN_B1_enable_value_O[0];
assign SB_T2_EAST_SB_IN_B1_ready_out = WIRE_SB_T2_EAST_SB_IN_B1_ready_out;
assign SB_T2_EAST_SB_OUT_B1 = RMUX_T2_EAST_B1_O;
assign SB_T2_EAST_SB_OUT_B1_enable = SB_T2_EAST_SB_OUT_B1_enable_value_O[0];
assign SB_T2_EAST_SB_OUT_B1_valid_out = RMUX_T2_EAST_B1_valid_out;
assign SB_T2_NORTH_SB_IN_B1_enable = SB_T2_NORTH_SB_IN_B1_enable_value_O[0];
assign SB_T2_NORTH_SB_IN_B1_ready_out = WIRE_SB_T2_NORTH_SB_IN_B1_ready_out;
assign SB_T2_NORTH_SB_OUT_B1 = RMUX_T2_NORTH_B1_O;
assign SB_T2_NORTH_SB_OUT_B1_enable = SB_T2_NORTH_SB_OUT_B1_enable_value_O[0];
assign SB_T2_NORTH_SB_OUT_B1_valid_out = RMUX_T2_NORTH_B1_valid_out;
assign SB_T2_SOUTH_SB_IN_B1_enable = SB_T2_SOUTH_SB_IN_B1_enable_value_O[0];
assign SB_T2_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T2_SOUTH_SB_IN_B1_ready_out;
assign SB_T2_SOUTH_SB_OUT_B1 = RMUX_T2_SOUTH_B1_O;
assign SB_T2_SOUTH_SB_OUT_B1_enable = SB_T2_SOUTH_SB_OUT_B1_enable_value_O[0];
assign SB_T2_SOUTH_SB_OUT_B1_valid_out = RMUX_T2_SOUTH_B1_valid_out;
assign SB_T2_WEST_SB_IN_B1_enable = SB_T2_WEST_SB_IN_B1_enable_value_O[0];
assign SB_T2_WEST_SB_IN_B1_ready_out = WIRE_SB_T2_WEST_SB_IN_B1_ready_out;
assign SB_T2_WEST_SB_OUT_B1 = RMUX_T2_WEST_B1_O;
assign SB_T2_WEST_SB_OUT_B1_enable = SB_T2_WEST_SB_OUT_B1_enable_value_O[0];
assign SB_T2_WEST_SB_OUT_B1_valid_out = RMUX_T2_WEST_B1_valid_out;
assign SB_T3_EAST_SB_IN_B1_enable = SB_T3_EAST_SB_IN_B1_enable_value_O[0];
assign SB_T3_EAST_SB_IN_B1_ready_out = WIRE_SB_T3_EAST_SB_IN_B1_ready_out;
assign SB_T3_EAST_SB_OUT_B1 = RMUX_T3_EAST_B1_O;
assign SB_T3_EAST_SB_OUT_B1_enable = SB_T3_EAST_SB_OUT_B1_enable_value_O[0];
assign SB_T3_EAST_SB_OUT_B1_valid_out = RMUX_T3_EAST_B1_valid_out;
assign SB_T3_NORTH_SB_IN_B1_enable = SB_T3_NORTH_SB_IN_B1_enable_value_O[0];
assign SB_T3_NORTH_SB_IN_B1_ready_out = WIRE_SB_T3_NORTH_SB_IN_B1_ready_out;
assign SB_T3_NORTH_SB_OUT_B1 = RMUX_T3_NORTH_B1_O;
assign SB_T3_NORTH_SB_OUT_B1_enable = SB_T3_NORTH_SB_OUT_B1_enable_value_O[0];
assign SB_T3_NORTH_SB_OUT_B1_valid_out = RMUX_T3_NORTH_B1_valid_out;
assign SB_T3_SOUTH_SB_IN_B1_enable = SB_T3_SOUTH_SB_IN_B1_enable_value_O[0];
assign SB_T3_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T3_SOUTH_SB_IN_B1_ready_out;
assign SB_T3_SOUTH_SB_OUT_B1 = RMUX_T3_SOUTH_B1_O;
assign SB_T3_SOUTH_SB_OUT_B1_enable = SB_T3_SOUTH_SB_OUT_B1_enable_value_O[0];
assign SB_T3_SOUTH_SB_OUT_B1_valid_out = RMUX_T3_SOUTH_B1_valid_out;
assign SB_T3_WEST_SB_IN_B1_enable = SB_T3_WEST_SB_IN_B1_enable_value_O[0];
assign SB_T3_WEST_SB_IN_B1_ready_out = WIRE_SB_T3_WEST_SB_IN_B1_ready_out;
assign SB_T3_WEST_SB_OUT_B1 = RMUX_T3_WEST_B1_O;
assign SB_T3_WEST_SB_OUT_B1_enable = SB_T3_WEST_SB_OUT_B1_enable_value_O[0];
assign SB_T3_WEST_SB_OUT_B1_valid_out = RMUX_T3_WEST_B1_valid_out;
assign SB_T4_EAST_SB_IN_B1_enable = SB_T4_EAST_SB_IN_B1_enable_value_O[0];
assign SB_T4_EAST_SB_IN_B1_ready_out = WIRE_SB_T4_EAST_SB_IN_B1_ready_out;
assign SB_T4_EAST_SB_OUT_B1 = RMUX_T4_EAST_B1_O;
assign SB_T4_EAST_SB_OUT_B1_enable = SB_T4_EAST_SB_OUT_B1_enable_value_O[0];
assign SB_T4_EAST_SB_OUT_B1_valid_out = RMUX_T4_EAST_B1_valid_out;
assign SB_T4_NORTH_SB_IN_B1_enable = SB_T4_NORTH_SB_IN_B1_enable_value_O[0];
assign SB_T4_NORTH_SB_IN_B1_ready_out = WIRE_SB_T4_NORTH_SB_IN_B1_ready_out;
assign SB_T4_NORTH_SB_OUT_B1 = RMUX_T4_NORTH_B1_O;
assign SB_T4_NORTH_SB_OUT_B1_enable = SB_T4_NORTH_SB_OUT_B1_enable_value_O[0];
assign SB_T4_NORTH_SB_OUT_B1_valid_out = RMUX_T4_NORTH_B1_valid_out;
assign SB_T4_SOUTH_SB_IN_B1_enable = SB_T4_SOUTH_SB_IN_B1_enable_value_O[0];
assign SB_T4_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T4_SOUTH_SB_IN_B1_ready_out;
assign SB_T4_SOUTH_SB_OUT_B1 = RMUX_T4_SOUTH_B1_O;
assign SB_T4_SOUTH_SB_OUT_B1_enable = SB_T4_SOUTH_SB_OUT_B1_enable_value_O[0];
assign SB_T4_SOUTH_SB_OUT_B1_valid_out = RMUX_T4_SOUTH_B1_valid_out;
assign SB_T4_WEST_SB_IN_B1_enable = SB_T4_WEST_SB_IN_B1_enable_value_O[0];
assign SB_T4_WEST_SB_IN_B1_ready_out = WIRE_SB_T4_WEST_SB_IN_B1_ready_out;
assign SB_T4_WEST_SB_OUT_B1 = RMUX_T4_WEST_B1_O;
assign SB_T4_WEST_SB_OUT_B1_enable = SB_T4_WEST_SB_OUT_B1_enable_value_O[0];
assign SB_T4_WEST_SB_OUT_B1_valid_out = RMUX_T4_WEST_B1_valid_out;
assign read_config_data = mux_aoi_6_32_inst0_O;
endmodule

module SB_ID0_5TRACKS_B1_MemCore (
    input [0:0] MEM_input_width_1_num_0_enable,
    input [31:0] MEM_input_width_1_num_0_out_sel,
    input MEM_input_width_1_num_0_ready,
    input [0:0] MEM_input_width_1_num_1_enable,
    input [31:0] MEM_input_width_1_num_1_out_sel,
    input MEM_input_width_1_num_1_ready,
    input [0:0] MEM_output_width_1_num_0,
    output MEM_output_width_1_num_0_ready_out,
    input MEM_output_width_1_num_0_valid,
    input [0:0] MEM_output_width_1_num_1,
    output MEM_output_width_1_num_1_ready_out,
    input MEM_output_width_1_num_1_valid,
    input [0:0] MEM_output_width_1_num_2,
    output MEM_output_width_1_num_2_ready_out,
    input MEM_output_width_1_num_2_valid,
    input [0:0] SB_T0_EAST_SB_IN_B1,
    output SB_T0_EAST_SB_IN_B1_enable,
    output SB_T0_EAST_SB_IN_B1_ready_out,
    input SB_T0_EAST_SB_IN_B1_valid_in,
    output [0:0] SB_T0_EAST_SB_OUT_B1,
    output SB_T0_EAST_SB_OUT_B1_enable,
    input SB_T0_EAST_SB_OUT_B1_ready_in,
    output SB_T0_EAST_SB_OUT_B1_valid_out,
    input [0:0] SB_T0_NORTH_SB_IN_B1,
    output SB_T0_NORTH_SB_IN_B1_enable,
    output SB_T0_NORTH_SB_IN_B1_ready_out,
    input SB_T0_NORTH_SB_IN_B1_valid_in,
    output [0:0] SB_T0_NORTH_SB_OUT_B1,
    output SB_T0_NORTH_SB_OUT_B1_enable,
    input SB_T0_NORTH_SB_OUT_B1_ready_in,
    output SB_T0_NORTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T0_SOUTH_SB_IN_B1,
    output SB_T0_SOUTH_SB_IN_B1_enable,
    output SB_T0_SOUTH_SB_IN_B1_ready_out,
    input SB_T0_SOUTH_SB_IN_B1_valid_in,
    output [0:0] SB_T0_SOUTH_SB_OUT_B1,
    output SB_T0_SOUTH_SB_OUT_B1_enable,
    input SB_T0_SOUTH_SB_OUT_B1_ready_in,
    output SB_T0_SOUTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T0_WEST_SB_IN_B1,
    output SB_T0_WEST_SB_IN_B1_enable,
    output SB_T0_WEST_SB_IN_B1_ready_out,
    input SB_T0_WEST_SB_IN_B1_valid_in,
    output [0:0] SB_T0_WEST_SB_OUT_B1,
    output SB_T0_WEST_SB_OUT_B1_enable,
    input SB_T0_WEST_SB_OUT_B1_ready_in,
    output SB_T0_WEST_SB_OUT_B1_valid_out,
    input [0:0] SB_T1_EAST_SB_IN_B1,
    output SB_T1_EAST_SB_IN_B1_enable,
    output SB_T1_EAST_SB_IN_B1_ready_out,
    input SB_T1_EAST_SB_IN_B1_valid_in,
    output [0:0] SB_T1_EAST_SB_OUT_B1,
    output SB_T1_EAST_SB_OUT_B1_enable,
    input SB_T1_EAST_SB_OUT_B1_ready_in,
    output SB_T1_EAST_SB_OUT_B1_valid_out,
    input [0:0] SB_T1_NORTH_SB_IN_B1,
    output SB_T1_NORTH_SB_IN_B1_enable,
    output SB_T1_NORTH_SB_IN_B1_ready_out,
    input SB_T1_NORTH_SB_IN_B1_valid_in,
    output [0:0] SB_T1_NORTH_SB_OUT_B1,
    output SB_T1_NORTH_SB_OUT_B1_enable,
    input SB_T1_NORTH_SB_OUT_B1_ready_in,
    output SB_T1_NORTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T1_SOUTH_SB_IN_B1,
    output SB_T1_SOUTH_SB_IN_B1_enable,
    output SB_T1_SOUTH_SB_IN_B1_ready_out,
    input SB_T1_SOUTH_SB_IN_B1_valid_in,
    output [0:0] SB_T1_SOUTH_SB_OUT_B1,
    output SB_T1_SOUTH_SB_OUT_B1_enable,
    input SB_T1_SOUTH_SB_OUT_B1_ready_in,
    output SB_T1_SOUTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T1_WEST_SB_IN_B1,
    output SB_T1_WEST_SB_IN_B1_enable,
    output SB_T1_WEST_SB_IN_B1_ready_out,
    input SB_T1_WEST_SB_IN_B1_valid_in,
    output [0:0] SB_T1_WEST_SB_OUT_B1,
    output SB_T1_WEST_SB_OUT_B1_enable,
    input SB_T1_WEST_SB_OUT_B1_ready_in,
    output SB_T1_WEST_SB_OUT_B1_valid_out,
    input [0:0] SB_T2_EAST_SB_IN_B1,
    output SB_T2_EAST_SB_IN_B1_enable,
    output SB_T2_EAST_SB_IN_B1_ready_out,
    input SB_T2_EAST_SB_IN_B1_valid_in,
    output [0:0] SB_T2_EAST_SB_OUT_B1,
    output SB_T2_EAST_SB_OUT_B1_enable,
    input SB_T2_EAST_SB_OUT_B1_ready_in,
    output SB_T2_EAST_SB_OUT_B1_valid_out,
    input [0:0] SB_T2_NORTH_SB_IN_B1,
    output SB_T2_NORTH_SB_IN_B1_enable,
    output SB_T2_NORTH_SB_IN_B1_ready_out,
    input SB_T2_NORTH_SB_IN_B1_valid_in,
    output [0:0] SB_T2_NORTH_SB_OUT_B1,
    output SB_T2_NORTH_SB_OUT_B1_enable,
    input SB_T2_NORTH_SB_OUT_B1_ready_in,
    output SB_T2_NORTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T2_SOUTH_SB_IN_B1,
    output SB_T2_SOUTH_SB_IN_B1_enable,
    output SB_T2_SOUTH_SB_IN_B1_ready_out,
    input SB_T2_SOUTH_SB_IN_B1_valid_in,
    output [0:0] SB_T2_SOUTH_SB_OUT_B1,
    output SB_T2_SOUTH_SB_OUT_B1_enable,
    input SB_T2_SOUTH_SB_OUT_B1_ready_in,
    output SB_T2_SOUTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T2_WEST_SB_IN_B1,
    output SB_T2_WEST_SB_IN_B1_enable,
    output SB_T2_WEST_SB_IN_B1_ready_out,
    input SB_T2_WEST_SB_IN_B1_valid_in,
    output [0:0] SB_T2_WEST_SB_OUT_B1,
    output SB_T2_WEST_SB_OUT_B1_enable,
    input SB_T2_WEST_SB_OUT_B1_ready_in,
    output SB_T2_WEST_SB_OUT_B1_valid_out,
    input [0:0] SB_T3_EAST_SB_IN_B1,
    output SB_T3_EAST_SB_IN_B1_enable,
    output SB_T3_EAST_SB_IN_B1_ready_out,
    input SB_T3_EAST_SB_IN_B1_valid_in,
    output [0:0] SB_T3_EAST_SB_OUT_B1,
    output SB_T3_EAST_SB_OUT_B1_enable,
    input SB_T3_EAST_SB_OUT_B1_ready_in,
    output SB_T3_EAST_SB_OUT_B1_valid_out,
    input [0:0] SB_T3_NORTH_SB_IN_B1,
    output SB_T3_NORTH_SB_IN_B1_enable,
    output SB_T3_NORTH_SB_IN_B1_ready_out,
    input SB_T3_NORTH_SB_IN_B1_valid_in,
    output [0:0] SB_T3_NORTH_SB_OUT_B1,
    output SB_T3_NORTH_SB_OUT_B1_enable,
    input SB_T3_NORTH_SB_OUT_B1_ready_in,
    output SB_T3_NORTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T3_SOUTH_SB_IN_B1,
    output SB_T3_SOUTH_SB_IN_B1_enable,
    output SB_T3_SOUTH_SB_IN_B1_ready_out,
    input SB_T3_SOUTH_SB_IN_B1_valid_in,
    output [0:0] SB_T3_SOUTH_SB_OUT_B1,
    output SB_T3_SOUTH_SB_OUT_B1_enable,
    input SB_T3_SOUTH_SB_OUT_B1_ready_in,
    output SB_T3_SOUTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T3_WEST_SB_IN_B1,
    output SB_T3_WEST_SB_IN_B1_enable,
    output SB_T3_WEST_SB_IN_B1_ready_out,
    input SB_T3_WEST_SB_IN_B1_valid_in,
    output [0:0] SB_T3_WEST_SB_OUT_B1,
    output SB_T3_WEST_SB_OUT_B1_enable,
    input SB_T3_WEST_SB_OUT_B1_ready_in,
    output SB_T3_WEST_SB_OUT_B1_valid_out,
    input [0:0] SB_T4_EAST_SB_IN_B1,
    output SB_T4_EAST_SB_IN_B1_enable,
    output SB_T4_EAST_SB_IN_B1_ready_out,
    input SB_T4_EAST_SB_IN_B1_valid_in,
    output [0:0] SB_T4_EAST_SB_OUT_B1,
    output SB_T4_EAST_SB_OUT_B1_enable,
    input SB_T4_EAST_SB_OUT_B1_ready_in,
    output SB_T4_EAST_SB_OUT_B1_valid_out,
    input [0:0] SB_T4_NORTH_SB_IN_B1,
    output SB_T4_NORTH_SB_IN_B1_enable,
    output SB_T4_NORTH_SB_IN_B1_ready_out,
    input SB_T4_NORTH_SB_IN_B1_valid_in,
    output [0:0] SB_T4_NORTH_SB_OUT_B1,
    output SB_T4_NORTH_SB_OUT_B1_enable,
    input SB_T4_NORTH_SB_OUT_B1_ready_in,
    output SB_T4_NORTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T4_SOUTH_SB_IN_B1,
    output SB_T4_SOUTH_SB_IN_B1_enable,
    output SB_T4_SOUTH_SB_IN_B1_ready_out,
    input SB_T4_SOUTH_SB_IN_B1_valid_in,
    output [0:0] SB_T4_SOUTH_SB_OUT_B1,
    output SB_T4_SOUTH_SB_OUT_B1_enable,
    input SB_T4_SOUTH_SB_OUT_B1_ready_in,
    output SB_T4_SOUTH_SB_OUT_B1_valid_out,
    input [0:0] SB_T4_WEST_SB_IN_B1,
    output SB_T4_WEST_SB_IN_B1_enable,
    output SB_T4_WEST_SB_IN_B1_ready_out,
    input SB_T4_WEST_SB_IN_B1_valid_in,
    output [0:0] SB_T4_WEST_SB_OUT_B1,
    output SB_T4_WEST_SB_OUT_B1_enable,
    input SB_T4_WEST_SB_OUT_B1_ready_in,
    output SB_T4_WEST_SB_OUT_B1_valid_out,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset,
    input [0:0] stall
);
wire [0:0] CB_MEM_output_width_1_num_0_fan_in_O;
wire [0:0] CB_MEM_output_width_1_num_1_fan_in_O;
wire [0:0] CB_MEM_output_width_1_num_2_fan_in_O;
wire [0:0] Invert1_inst0_out;
wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1_O;
wire MUX_SB_T0_EAST_SB_OUT_B1_ready_out;
wire MUX_SB_T0_EAST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T0_EAST_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1_O;
wire MUX_SB_T0_NORTH_SB_OUT_B1_ready_out;
wire MUX_SB_T0_NORTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T0_NORTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1_O;
wire MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out;
wire MUX_SB_T0_SOUTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1_O;
wire MUX_SB_T0_WEST_SB_OUT_B1_ready_out;
wire MUX_SB_T0_WEST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T0_WEST_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1_O;
wire MUX_SB_T1_EAST_SB_OUT_B1_ready_out;
wire MUX_SB_T1_EAST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T1_EAST_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1_O;
wire MUX_SB_T1_NORTH_SB_OUT_B1_ready_out;
wire MUX_SB_T1_NORTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T1_NORTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1_O;
wire MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out;
wire MUX_SB_T1_SOUTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1_O;
wire MUX_SB_T1_WEST_SB_OUT_B1_ready_out;
wire MUX_SB_T1_WEST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T1_WEST_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1_O;
wire MUX_SB_T2_EAST_SB_OUT_B1_ready_out;
wire MUX_SB_T2_EAST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T2_EAST_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1_O;
wire MUX_SB_T2_NORTH_SB_OUT_B1_ready_out;
wire MUX_SB_T2_NORTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T2_NORTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1_O;
wire MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out;
wire MUX_SB_T2_SOUTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1_O;
wire MUX_SB_T2_WEST_SB_OUT_B1_ready_out;
wire MUX_SB_T2_WEST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T2_WEST_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1_O;
wire MUX_SB_T3_EAST_SB_OUT_B1_ready_out;
wire MUX_SB_T3_EAST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T3_EAST_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1_O;
wire MUX_SB_T3_NORTH_SB_OUT_B1_ready_out;
wire MUX_SB_T3_NORTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T3_NORTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1_O;
wire MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out;
wire MUX_SB_T3_SOUTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1_O;
wire MUX_SB_T3_WEST_SB_OUT_B1_ready_out;
wire MUX_SB_T3_WEST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T3_WEST_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1_O;
wire MUX_SB_T4_EAST_SB_OUT_B1_ready_out;
wire MUX_SB_T4_EAST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T4_EAST_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1_O;
wire MUX_SB_T4_NORTH_SB_OUT_B1_ready_out;
wire MUX_SB_T4_NORTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T4_NORTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1_O;
wire MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out;
wire MUX_SB_T4_SOUTH_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel;
wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1_O;
wire MUX_SB_T4_WEST_SB_OUT_B1_ready_out;
wire MUX_SB_T4_WEST_SB_OUT_B1_valid_out;
wire [7:0] MUX_SB_T4_WEST_SB_OUT_B1_out_sel;
wire [0:0] REG_T0_EAST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T0_EAST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T0_EAST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T0_EAST_B1_end_value_O;
wire [0:0] REG_T0_EAST_B1_fifo_value_O;
wire [0:0] REG_T0_EAST_B1_start_value_O;
wire [0:0] REG_T0_NORTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T0_NORTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T0_NORTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T0_NORTH_B1_end_value_O;
wire [0:0] REG_T0_NORTH_B1_fifo_value_O;
wire [0:0] REG_T0_NORTH_B1_start_value_O;
wire [0:0] REG_T0_SOUTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T0_SOUTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T0_SOUTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T0_SOUTH_B1_end_value_O;
wire [0:0] REG_T0_SOUTH_B1_fifo_value_O;
wire [0:0] REG_T0_SOUTH_B1_start_value_O;
wire [0:0] REG_T0_WEST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T0_WEST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T0_WEST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T0_WEST_B1_end_value_O;
wire [0:0] REG_T0_WEST_B1_fifo_value_O;
wire [0:0] REG_T0_WEST_B1_start_value_O;
wire [0:0] REG_T1_EAST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T1_EAST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T1_EAST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T1_EAST_B1_end_value_O;
wire [0:0] REG_T1_EAST_B1_fifo_value_O;
wire [0:0] REG_T1_EAST_B1_start_value_O;
wire [0:0] REG_T1_NORTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T1_NORTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T1_NORTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T1_NORTH_B1_end_value_O;
wire [0:0] REG_T1_NORTH_B1_fifo_value_O;
wire [0:0] REG_T1_NORTH_B1_start_value_O;
wire [0:0] REG_T1_SOUTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T1_SOUTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T1_SOUTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T1_SOUTH_B1_end_value_O;
wire [0:0] REG_T1_SOUTH_B1_fifo_value_O;
wire [0:0] REG_T1_SOUTH_B1_start_value_O;
wire [0:0] REG_T1_WEST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T1_WEST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T1_WEST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T1_WEST_B1_end_value_O;
wire [0:0] REG_T1_WEST_B1_fifo_value_O;
wire [0:0] REG_T1_WEST_B1_start_value_O;
wire [0:0] REG_T2_EAST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T2_EAST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T2_EAST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T2_EAST_B1_end_value_O;
wire [0:0] REG_T2_EAST_B1_fifo_value_O;
wire [0:0] REG_T2_EAST_B1_start_value_O;
wire [0:0] REG_T2_NORTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T2_NORTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T2_NORTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T2_NORTH_B1_end_value_O;
wire [0:0] REG_T2_NORTH_B1_fifo_value_O;
wire [0:0] REG_T2_NORTH_B1_start_value_O;
wire [0:0] REG_T2_SOUTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T2_SOUTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T2_SOUTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T2_SOUTH_B1_end_value_O;
wire [0:0] REG_T2_SOUTH_B1_fifo_value_O;
wire [0:0] REG_T2_SOUTH_B1_start_value_O;
wire [0:0] REG_T2_WEST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T2_WEST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T2_WEST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T2_WEST_B1_end_value_O;
wire [0:0] REG_T2_WEST_B1_fifo_value_O;
wire [0:0] REG_T2_WEST_B1_start_value_O;
wire [0:0] REG_T3_EAST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T3_EAST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T3_EAST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T3_EAST_B1_end_value_O;
wire [0:0] REG_T3_EAST_B1_fifo_value_O;
wire [0:0] REG_T3_EAST_B1_start_value_O;
wire [0:0] REG_T3_NORTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T3_NORTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T3_NORTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T3_NORTH_B1_end_value_O;
wire [0:0] REG_T3_NORTH_B1_fifo_value_O;
wire [0:0] REG_T3_NORTH_B1_start_value_O;
wire [0:0] REG_T3_SOUTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T3_SOUTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T3_SOUTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T3_SOUTH_B1_end_value_O;
wire [0:0] REG_T3_SOUTH_B1_fifo_value_O;
wire [0:0] REG_T3_SOUTH_B1_start_value_O;
wire [0:0] REG_T3_WEST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T3_WEST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T3_WEST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T3_WEST_B1_end_value_O;
wire [0:0] REG_T3_WEST_B1_fifo_value_O;
wire [0:0] REG_T3_WEST_B1_start_value_O;
wire [0:0] REG_T4_EAST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T4_EAST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T4_EAST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T4_EAST_B1_end_value_O;
wire [0:0] REG_T4_EAST_B1_fifo_value_O;
wire [0:0] REG_T4_EAST_B1_start_value_O;
wire [0:0] REG_T4_NORTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T4_NORTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T4_NORTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T4_NORTH_B1_end_value_O;
wire [0:0] REG_T4_NORTH_B1_fifo_value_O;
wire [0:0] REG_T4_NORTH_B1_start_value_O;
wire [0:0] REG_T4_SOUTH_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T4_SOUTH_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T4_SOUTH_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T4_SOUTH_B1_end_value_O;
wire [0:0] REG_T4_SOUTH_B1_fifo_value_O;
wire [0:0] REG_T4_SOUTH_B1_start_value_O;
wire [0:0] REG_T4_WEST_B1$SplitFifo_1_inst0_ready0;
wire [0:0] REG_T4_WEST_B1$SplitFifo_1_inst0_valid1;
wire [0:0] REG_T4_WEST_B1$SplitFifo_1_inst0_data_out;
wire [0:0] REG_T4_WEST_B1_end_value_O;
wire [0:0] REG_T4_WEST_B1_fifo_value_O;
wire [0:0] REG_T4_WEST_B1_start_value_O;
wire [0:0] RMUX_T0_EAST_B1_O;
wire RMUX_T0_EAST_B1_ready_out;
wire RMUX_T0_EAST_B1_valid_out;
wire [1:0] RMUX_T0_EAST_B1_out_sel;
wire [0:0] RMUX_T0_EAST_B1_sel_value_O;
wire [0:0] RMUX_T0_NORTH_B1_O;
wire RMUX_T0_NORTH_B1_ready_out;
wire RMUX_T0_NORTH_B1_valid_out;
wire [1:0] RMUX_T0_NORTH_B1_out_sel;
wire [0:0] RMUX_T0_NORTH_B1_sel_value_O;
wire [0:0] RMUX_T0_SOUTH_B1_O;
wire RMUX_T0_SOUTH_B1_ready_out;
wire RMUX_T0_SOUTH_B1_valid_out;
wire [1:0] RMUX_T0_SOUTH_B1_out_sel;
wire [0:0] RMUX_T0_SOUTH_B1_sel_value_O;
wire [0:0] RMUX_T0_WEST_B1_O;
wire RMUX_T0_WEST_B1_ready_out;
wire RMUX_T0_WEST_B1_valid_out;
wire [1:0] RMUX_T0_WEST_B1_out_sel;
wire [0:0] RMUX_T0_WEST_B1_sel_value_O;
wire [0:0] RMUX_T1_EAST_B1_O;
wire RMUX_T1_EAST_B1_ready_out;
wire RMUX_T1_EAST_B1_valid_out;
wire [1:0] RMUX_T1_EAST_B1_out_sel;
wire [0:0] RMUX_T1_EAST_B1_sel_value_O;
wire [0:0] RMUX_T1_NORTH_B1_O;
wire RMUX_T1_NORTH_B1_ready_out;
wire RMUX_T1_NORTH_B1_valid_out;
wire [1:0] RMUX_T1_NORTH_B1_out_sel;
wire [0:0] RMUX_T1_NORTH_B1_sel_value_O;
wire [0:0] RMUX_T1_SOUTH_B1_O;
wire RMUX_T1_SOUTH_B1_ready_out;
wire RMUX_T1_SOUTH_B1_valid_out;
wire [1:0] RMUX_T1_SOUTH_B1_out_sel;
wire [0:0] RMUX_T1_SOUTH_B1_sel_value_O;
wire [0:0] RMUX_T1_WEST_B1_O;
wire RMUX_T1_WEST_B1_ready_out;
wire RMUX_T1_WEST_B1_valid_out;
wire [1:0] RMUX_T1_WEST_B1_out_sel;
wire [0:0] RMUX_T1_WEST_B1_sel_value_O;
wire [0:0] RMUX_T2_EAST_B1_O;
wire RMUX_T2_EAST_B1_ready_out;
wire RMUX_T2_EAST_B1_valid_out;
wire [1:0] RMUX_T2_EAST_B1_out_sel;
wire [0:0] RMUX_T2_EAST_B1_sel_value_O;
wire [0:0] RMUX_T2_NORTH_B1_O;
wire RMUX_T2_NORTH_B1_ready_out;
wire RMUX_T2_NORTH_B1_valid_out;
wire [1:0] RMUX_T2_NORTH_B1_out_sel;
wire [0:0] RMUX_T2_NORTH_B1_sel_value_O;
wire [0:0] RMUX_T2_SOUTH_B1_O;
wire RMUX_T2_SOUTH_B1_ready_out;
wire RMUX_T2_SOUTH_B1_valid_out;
wire [1:0] RMUX_T2_SOUTH_B1_out_sel;
wire [0:0] RMUX_T2_SOUTH_B1_sel_value_O;
wire [0:0] RMUX_T2_WEST_B1_O;
wire RMUX_T2_WEST_B1_ready_out;
wire RMUX_T2_WEST_B1_valid_out;
wire [1:0] RMUX_T2_WEST_B1_out_sel;
wire [0:0] RMUX_T2_WEST_B1_sel_value_O;
wire [0:0] RMUX_T3_EAST_B1_O;
wire RMUX_T3_EAST_B1_ready_out;
wire RMUX_T3_EAST_B1_valid_out;
wire [1:0] RMUX_T3_EAST_B1_out_sel;
wire [0:0] RMUX_T3_EAST_B1_sel_value_O;
wire [0:0] RMUX_T3_NORTH_B1_O;
wire RMUX_T3_NORTH_B1_ready_out;
wire RMUX_T3_NORTH_B1_valid_out;
wire [1:0] RMUX_T3_NORTH_B1_out_sel;
wire [0:0] RMUX_T3_NORTH_B1_sel_value_O;
wire [0:0] RMUX_T3_SOUTH_B1_O;
wire RMUX_T3_SOUTH_B1_ready_out;
wire RMUX_T3_SOUTH_B1_valid_out;
wire [1:0] RMUX_T3_SOUTH_B1_out_sel;
wire [0:0] RMUX_T3_SOUTH_B1_sel_value_O;
wire [0:0] RMUX_T3_WEST_B1_O;
wire RMUX_T3_WEST_B1_ready_out;
wire RMUX_T3_WEST_B1_valid_out;
wire [1:0] RMUX_T3_WEST_B1_out_sel;
wire [0:0] RMUX_T3_WEST_B1_sel_value_O;
wire [0:0] RMUX_T4_EAST_B1_O;
wire RMUX_T4_EAST_B1_ready_out;
wire RMUX_T4_EAST_B1_valid_out;
wire [1:0] RMUX_T4_EAST_B1_out_sel;
wire [0:0] RMUX_T4_EAST_B1_sel_value_O;
wire [0:0] RMUX_T4_NORTH_B1_O;
wire RMUX_T4_NORTH_B1_ready_out;
wire RMUX_T4_NORTH_B1_valid_out;
wire [1:0] RMUX_T4_NORTH_B1_out_sel;
wire [0:0] RMUX_T4_NORTH_B1_sel_value_O;
wire [0:0] RMUX_T4_SOUTH_B1_O;
wire RMUX_T4_SOUTH_B1_ready_out;
wire RMUX_T4_SOUTH_B1_valid_out;
wire [1:0] RMUX_T4_SOUTH_B1_out_sel;
wire [0:0] RMUX_T4_SOUTH_B1_sel_value_O;
wire [0:0] RMUX_T4_WEST_B1_O;
wire RMUX_T4_WEST_B1_ready_out;
wire RMUX_T4_WEST_B1_valid_out;
wire [1:0] RMUX_T4_WEST_B1_out_sel;
wire [0:0] RMUX_T4_WEST_B1_sel_value_O;
wire [0:0] SB_T0_EAST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T0_EAST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T0_EAST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T0_EAST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T0_EAST_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T0_NORTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T0_NORTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T0_NORTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T0_NORTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T0_NORTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T0_SOUTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T0_SOUTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T0_SOUTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T0_SOUTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T0_SOUTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T0_WEST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T0_WEST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T0_WEST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T0_WEST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T0_WEST_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T1_EAST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T1_EAST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T1_EAST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T1_EAST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T1_EAST_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T1_NORTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T1_NORTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T1_NORTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T1_NORTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T1_NORTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T1_SOUTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T1_SOUTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T1_SOUTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T1_SOUTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T1_SOUTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T1_WEST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T1_WEST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T1_WEST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T1_WEST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T1_WEST_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T2_EAST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T2_EAST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T2_EAST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T2_EAST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T2_EAST_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T2_NORTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T2_NORTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T2_NORTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T2_NORTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T2_NORTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T2_SOUTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T2_SOUTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T2_SOUTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T2_SOUTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T2_SOUTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T2_WEST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T2_WEST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T2_WEST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T2_WEST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T2_WEST_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T3_EAST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T3_EAST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T3_EAST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T3_EAST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T3_EAST_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T3_NORTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T3_NORTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T3_NORTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T3_NORTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T3_NORTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T3_SOUTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T3_SOUTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T3_SOUTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T3_SOUTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T3_SOUTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T3_WEST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T3_WEST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T3_WEST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T3_WEST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T3_WEST_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T4_EAST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T4_EAST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T4_EAST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T4_EAST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T4_EAST_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T4_NORTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T4_NORTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T4_NORTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T4_NORTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T4_NORTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T4_SOUTH_SB_IN_B1_enable_value_O;
wire [0:0] SB_T4_SOUTH_SB_IN_B1_fan_in_O;
wire [0:0] SB_T4_SOUTH_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T4_SOUTH_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T4_SOUTH_SB_OUT_B1_sel_value_O;
wire [0:0] SB_T4_WEST_SB_IN_B1_enable_value_O;
wire [0:0] SB_T4_WEST_SB_IN_B1_fan_in_O;
wire [0:0] SB_T4_WEST_SB_OUT_B1_FANOUT_O;
wire [0:0] SB_T4_WEST_SB_OUT_B1_enable_value_O;
wire [2:0] SB_T4_WEST_SB_OUT_B1_sel_value_O;
wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1_O;
wire WIRE_SB_T0_EAST_SB_IN_B1_ready_out;
wire WIRE_SB_T0_EAST_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1_O;
wire WIRE_SB_T0_NORTH_SB_IN_B1_ready_out;
wire WIRE_SB_T0_NORTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1_O;
wire WIRE_SB_T0_SOUTH_SB_IN_B1_ready_out;
wire WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1_O;
wire WIRE_SB_T0_WEST_SB_IN_B1_ready_out;
wire WIRE_SB_T0_WEST_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1_O;
wire WIRE_SB_T1_EAST_SB_IN_B1_ready_out;
wire WIRE_SB_T1_EAST_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1_O;
wire WIRE_SB_T1_NORTH_SB_IN_B1_ready_out;
wire WIRE_SB_T1_NORTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1_O;
wire WIRE_SB_T1_SOUTH_SB_IN_B1_ready_out;
wire WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1_O;
wire WIRE_SB_T1_WEST_SB_IN_B1_ready_out;
wire WIRE_SB_T1_WEST_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1_O;
wire WIRE_SB_T2_EAST_SB_IN_B1_ready_out;
wire WIRE_SB_T2_EAST_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1_O;
wire WIRE_SB_T2_NORTH_SB_IN_B1_ready_out;
wire WIRE_SB_T2_NORTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1_O;
wire WIRE_SB_T2_SOUTH_SB_IN_B1_ready_out;
wire WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1_O;
wire WIRE_SB_T2_WEST_SB_IN_B1_ready_out;
wire WIRE_SB_T2_WEST_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1_O;
wire WIRE_SB_T3_EAST_SB_IN_B1_ready_out;
wire WIRE_SB_T3_EAST_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1_O;
wire WIRE_SB_T3_NORTH_SB_IN_B1_ready_out;
wire WIRE_SB_T3_NORTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1_O;
wire WIRE_SB_T3_SOUTH_SB_IN_B1_ready_out;
wire WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1_O;
wire WIRE_SB_T3_WEST_SB_IN_B1_ready_out;
wire WIRE_SB_T3_WEST_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1_O;
wire WIRE_SB_T4_EAST_SB_IN_B1_ready_out;
wire WIRE_SB_T4_EAST_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1_O;
wire WIRE_SB_T4_NORTH_SB_IN_B1_ready_out;
wire WIRE_SB_T4_NORTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1_O;
wire WIRE_SB_T4_SOUTH_SB_IN_B1_ready_out;
wire WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out;
wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1_O;
wire WIRE_SB_T4_WEST_SB_IN_B1_ready_out;
wire WIRE_SB_T4_WEST_SB_IN_B1_valid_out;
wire ZextWrapper_23_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_23_32_inst0$self_O_in;
wire ZextWrapper_30_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_30_32_inst0$self_O_in;
wire ZextWrapper_31_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_31_32_inst0$self_O_in;
wire [0:0] and1_inst0_out;
wire [0:0] and1_inst1_out;
wire [0:0] and1_inst10_out;
wire [0:0] and1_inst11_out;
wire [0:0] and1_inst12_out;
wire [0:0] and1_inst13_out;
wire [0:0] and1_inst14_out;
wire [0:0] and1_inst15_out;
wire [0:0] and1_inst16_out;
wire [0:0] and1_inst17_out;
wire [0:0] and1_inst18_out;
wire [0:0] and1_inst19_out;
wire [0:0] and1_inst2_out;
wire [0:0] and1_inst3_out;
wire [0:0] and1_inst4_out;
wire [0:0] and1_inst5_out;
wire [0:0] and1_inst6_out;
wire [0:0] and1_inst7_out;
wire [0:0] and1_inst8_out;
wire [0:0] and1_inst9_out;
wire [31:0] config_reg_0_O;
wire [31:0] config_reg_1_O;
wire [31:0] config_reg_2_O;
wire [30:0] config_reg_3_O;
wire [29:0] config_reg_4_O;
wire [22:0] config_reg_5_O;
wire [0:0] const_0_1_out;
wire [31:0] const_0_32_out;
wire [0:0] const_1_1_out;
wire coreir_eq_1_inst0_out;
wire coreir_eq_1_inst1_out;
wire coreir_eq_1_inst10_out;
wire coreir_eq_1_inst11_out;
wire coreir_eq_1_inst12_out;
wire coreir_eq_1_inst13_out;
wire coreir_eq_1_inst14_out;
wire coreir_eq_1_inst15_out;
wire coreir_eq_1_inst16_out;
wire coreir_eq_1_inst17_out;
wire coreir_eq_1_inst18_out;
wire coreir_eq_1_inst19_out;
wire coreir_eq_1_inst2_out;
wire coreir_eq_1_inst3_out;
wire coreir_eq_1_inst4_out;
wire coreir_eq_1_inst5_out;
wire coreir_eq_1_inst6_out;
wire coreir_eq_1_inst7_out;
wire coreir_eq_1_inst8_out;
wire coreir_eq_1_inst9_out;
wire [31:0] mux_aoi_6_32_inst0_O;
wire [7:0] mux_aoi_6_32_inst0_out_sel;
wire [7:0] self_config_config_addr_out;
FanoutHash_E70AF988E4250F5 CB_MEM_output_width_1_num_0_fan_in (
    .S13(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
    .E13(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
    .S6(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
    .E2(SB_T0_EAST_SB_OUT_B1_enable_value_O),
    .E12(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
    .E7(SB_T1_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
    .E18(SB_T4_EAST_SB_OUT_B1_enable_value_O),
    .I3(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
    .E19(SB_T4_WEST_SB_OUT_B1_enable_value_O),
    .I14(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
    .S14(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
    .I9(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
    .S12(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
    .S17(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
    .I13(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
    .S9(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
    .E10(SB_T2_EAST_SB_OUT_B1_enable_value_O),
    .E15(SB_T3_WEST_SB_OUT_B1_enable_value_O),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
    .E5(SB_T1_SOUTH_SB_OUT_B1_enable_value_O),
    .S10(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
    .E8(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
    .I11(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
    .I6(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
    .S15(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
    .I7(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
    .E14(SB_T3_EAST_SB_OUT_B1_enable_value_O),
    .I2(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
    .E11(SB_T2_WEST_SB_OUT_B1_enable_value_O),
    .S3(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
    .S8(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
    .I10(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
    .S16(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
    .E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
    .E16(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
    .E3(SB_T0_WEST_SB_OUT_B1_enable_value_O),
    .S18(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
    .S19(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
    .S2(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
    .S4(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
    .E9(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
    .I16(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
    .I12(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
    .S11(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
    .I17(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
    .I19(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
    .I18(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
    .S7(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
    .E4(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
    .E17(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
    .S5(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
    .I1(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
    .I5(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
    .E6(SB_T1_EAST_SB_OUT_B1_enable_value_O),
    .I4(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
    .I8(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
    .O(CB_MEM_output_width_1_num_0_fan_in_O),
    .E1(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
    .I15(MUX_SB_T3_WEST_SB_OUT_B1_ready_out)
);
FanoutHash_82899D6851EDC11 CB_MEM_output_width_1_num_1_fan_in (
    .S13(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
    .E13(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
    .S6(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
    .E2(SB_T0_EAST_SB_OUT_B1_enable_value_O),
    .E12(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
    .E7(SB_T1_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
    .E18(SB_T4_EAST_SB_OUT_B1_enable_value_O),
    .I3(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
    .E19(SB_T4_WEST_SB_OUT_B1_enable_value_O),
    .I14(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
    .S14(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
    .I9(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
    .S12(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
    .S17(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
    .I13(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
    .S9(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
    .E10(SB_T2_EAST_SB_OUT_B1_enable_value_O),
    .E15(SB_T3_WEST_SB_OUT_B1_enable_value_O),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
    .E5(SB_T1_SOUTH_SB_OUT_B1_enable_value_O),
    .S10(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
    .E8(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
    .I11(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
    .I6(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
    .S15(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
    .I7(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
    .E14(SB_T3_EAST_SB_OUT_B1_enable_value_O),
    .I2(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
    .E11(SB_T2_WEST_SB_OUT_B1_enable_value_O),
    .S3(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
    .S8(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
    .I10(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
    .S16(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
    .E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
    .E16(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
    .E3(SB_T0_WEST_SB_OUT_B1_enable_value_O),
    .S18(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
    .S19(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
    .S2(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
    .S4(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
    .E9(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
    .I16(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
    .I12(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
    .S11(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
    .I17(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
    .I19(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
    .I18(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
    .S7(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
    .E4(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
    .E17(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
    .S5(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
    .I1(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
    .I5(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
    .E6(SB_T1_EAST_SB_OUT_B1_enable_value_O),
    .I4(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
    .I8(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
    .O(CB_MEM_output_width_1_num_1_fan_in_O),
    .E1(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
    .I15(MUX_SB_T3_WEST_SB_OUT_B1_ready_out)
);
FanoutHash_CE1AA874B742213 CB_MEM_output_width_1_num_2_fan_in (
    .S13(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
    .E13(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
    .S6(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
    .E2(SB_T0_EAST_SB_OUT_B1_enable_value_O),
    .E12(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
    .E7(SB_T1_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
    .E18(SB_T4_EAST_SB_OUT_B1_enable_value_O),
    .I3(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
    .E19(SB_T4_WEST_SB_OUT_B1_enable_value_O),
    .I14(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
    .S14(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
    .I9(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
    .S12(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
    .S17(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
    .I13(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
    .S9(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
    .E10(SB_T2_EAST_SB_OUT_B1_enable_value_O),
    .E15(SB_T3_WEST_SB_OUT_B1_enable_value_O),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
    .E5(SB_T1_SOUTH_SB_OUT_B1_enable_value_O),
    .S10(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
    .E8(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
    .I11(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
    .I6(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
    .S15(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
    .I7(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
    .E14(SB_T3_EAST_SB_OUT_B1_enable_value_O),
    .I2(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
    .E11(SB_T2_WEST_SB_OUT_B1_enable_value_O),
    .S3(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
    .S8(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
    .I10(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
    .S16(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
    .E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
    .E16(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
    .E3(SB_T0_WEST_SB_OUT_B1_enable_value_O),
    .S18(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
    .S19(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
    .S2(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
    .S4(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
    .E9(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
    .I16(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
    .I12(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
    .S11(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
    .I17(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
    .I19(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
    .I18(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
    .S7(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
    .E4(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
    .E17(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
    .S5(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
    .I1(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
    .I5(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
    .E6(SB_T1_EAST_SB_OUT_B1_enable_value_O),
    .I4(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
    .I8(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
    .O(CB_MEM_output_width_1_num_2_fan_in_O),
    .E1(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
    .I15(MUX_SB_T3_WEST_SB_OUT_B1_ready_out)
);
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(stall),
    .out(Invert1_inst0_out)
);
wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1_I [5:0];
assign MUX_SB_T0_EAST_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T0_EAST_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T0_EAST_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T0_EAST_SB_OUT_B1_I[2] = WIRE_SB_T4_NORTH_SB_IN_B1_O;
assign MUX_SB_T0_EAST_SB_OUT_B1_I[1] = WIRE_SB_T3_SOUTH_SB_IN_B1_O;
assign MUX_SB_T0_EAST_SB_OUT_B1_I[0] = WIRE_SB_T0_WEST_SB_IN_B1_O;
wire [5:0] MUX_SB_T0_EAST_SB_OUT_B1_valid_in;
assign MUX_SB_T0_EAST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T4_NORTH_SB_IN_B1_valid_out,WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T0_WEST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T0_EAST_SB_OUT_B1 (
    .I(MUX_SB_T0_EAST_SB_OUT_B1_I),
    .O(MUX_SB_T0_EAST_SB_OUT_B1_O),
    .ready_in(SB_T0_EAST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T0_EAST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T0_EAST_SB_OUT_B1_valid_out),
    .S(SB_T0_EAST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T0_EAST_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T0_NORTH_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T0_NORTH_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T0_NORTH_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T0_NORTH_SB_OUT_B1_I[2] = WIRE_SB_T0_SOUTH_SB_IN_B1_O;
assign MUX_SB_T0_NORTH_SB_OUT_B1_I[1] = WIRE_SB_T1_EAST_SB_IN_B1_O;
assign MUX_SB_T0_NORTH_SB_OUT_B1_I[0] = WIRE_SB_T0_WEST_SB_IN_B1_O;
wire [5:0] MUX_SB_T0_NORTH_SB_OUT_B1_valid_in;
assign MUX_SB_T0_NORTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T1_EAST_SB_IN_B1_valid_out,WIRE_SB_T0_WEST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T0_NORTH_SB_OUT_B1 (
    .I(MUX_SB_T0_NORTH_SB_OUT_B1_I),
    .O(MUX_SB_T0_NORTH_SB_OUT_B1_O),
    .ready_in(SB_T0_NORTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T0_NORTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T0_NORTH_SB_OUT_B1_valid_out),
    .S(SB_T0_NORTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[2] = WIRE_SB_T1_WEST_SB_IN_B1_O;
assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[1] = WIRE_SB_T0_NORTH_SB_IN_B1_O;
assign MUX_SB_T0_SOUTH_SB_OUT_B1_I[0] = WIRE_SB_T3_EAST_SB_IN_B1_O;
wire [5:0] MUX_SB_T0_SOUTH_SB_OUT_B1_valid_in;
assign MUX_SB_T0_SOUTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T1_WEST_SB_IN_B1_valid_out,WIRE_SB_T0_NORTH_SB_IN_B1_valid_out,WIRE_SB_T3_EAST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T0_SOUTH_SB_OUT_B1 (
    .I(MUX_SB_T0_SOUTH_SB_OUT_B1_I),
    .O(MUX_SB_T0_SOUTH_SB_OUT_B1_O),
    .ready_in(SB_T0_SOUTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T0_SOUTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T0_SOUTH_SB_OUT_B1_valid_out),
    .S(SB_T0_SOUTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1_I [5:0];
assign MUX_SB_T0_WEST_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T0_WEST_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T0_WEST_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T0_WEST_SB_OUT_B1_I[2] = WIRE_SB_T0_EAST_SB_IN_B1_O;
assign MUX_SB_T0_WEST_SB_OUT_B1_I[1] = WIRE_SB_T4_SOUTH_SB_IN_B1_O;
assign MUX_SB_T0_WEST_SB_OUT_B1_I[0] = WIRE_SB_T0_NORTH_SB_IN_B1_O;
wire [5:0] MUX_SB_T0_WEST_SB_OUT_B1_valid_in;
assign MUX_SB_T0_WEST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T0_EAST_SB_IN_B1_valid_out,WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T0_NORTH_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T0_WEST_SB_OUT_B1 (
    .I(MUX_SB_T0_WEST_SB_OUT_B1_I),
    .O(MUX_SB_T0_WEST_SB_OUT_B1_O),
    .ready_in(SB_T0_WEST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T0_WEST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T0_WEST_SB_OUT_B1_valid_out),
    .S(SB_T0_WEST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T0_WEST_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1_I [5:0];
assign MUX_SB_T1_EAST_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T1_EAST_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T1_EAST_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T1_EAST_SB_OUT_B1_I[2] = WIRE_SB_T2_SOUTH_SB_IN_B1_O;
assign MUX_SB_T1_EAST_SB_OUT_B1_I[1] = WIRE_SB_T1_WEST_SB_IN_B1_O;
assign MUX_SB_T1_EAST_SB_OUT_B1_I[0] = WIRE_SB_T0_NORTH_SB_IN_B1_O;
wire [5:0] MUX_SB_T1_EAST_SB_OUT_B1_valid_in;
assign MUX_SB_T1_EAST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T1_WEST_SB_IN_B1_valid_out,WIRE_SB_T0_NORTH_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T1_EAST_SB_OUT_B1 (
    .I(MUX_SB_T1_EAST_SB_OUT_B1_I),
    .O(MUX_SB_T1_EAST_SB_OUT_B1_O),
    .ready_in(SB_T1_EAST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T1_EAST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T1_EAST_SB_OUT_B1_valid_out),
    .S(SB_T1_EAST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T1_EAST_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T1_NORTH_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T1_NORTH_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T1_NORTH_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T1_NORTH_SB_OUT_B1_I[2] = WIRE_SB_T4_WEST_SB_IN_B1_O;
assign MUX_SB_T1_NORTH_SB_OUT_B1_I[1] = WIRE_SB_T1_SOUTH_SB_IN_B1_O;
assign MUX_SB_T1_NORTH_SB_OUT_B1_I[0] = WIRE_SB_T2_EAST_SB_IN_B1_O;
wire [5:0] MUX_SB_T1_NORTH_SB_OUT_B1_valid_in;
assign MUX_SB_T1_NORTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T4_WEST_SB_IN_B1_valid_out,WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T2_EAST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T1_NORTH_SB_OUT_B1 (
    .I(MUX_SB_T1_NORTH_SB_OUT_B1_I),
    .O(MUX_SB_T1_NORTH_SB_OUT_B1_O),
    .ready_in(SB_T1_NORTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T1_NORTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T1_NORTH_SB_OUT_B1_valid_out),
    .S(SB_T1_NORTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[2] = WIRE_SB_T2_WEST_SB_IN_B1_O;
assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[1] = WIRE_SB_T1_NORTH_SB_IN_B1_O;
assign MUX_SB_T1_SOUTH_SB_OUT_B1_I[0] = WIRE_SB_T2_EAST_SB_IN_B1_O;
wire [5:0] MUX_SB_T1_SOUTH_SB_OUT_B1_valid_in;
assign MUX_SB_T1_SOUTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T2_WEST_SB_IN_B1_valid_out,WIRE_SB_T1_NORTH_SB_IN_B1_valid_out,WIRE_SB_T2_EAST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T1_SOUTH_SB_OUT_B1 (
    .I(MUX_SB_T1_SOUTH_SB_OUT_B1_I),
    .O(MUX_SB_T1_SOUTH_SB_OUT_B1_O),
    .ready_in(SB_T1_SOUTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T1_SOUTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T1_SOUTH_SB_OUT_B1_valid_out),
    .S(SB_T1_SOUTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1_I [5:0];
assign MUX_SB_T1_WEST_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T1_WEST_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T1_WEST_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T1_WEST_SB_OUT_B1_I[2] = WIRE_SB_T1_EAST_SB_IN_B1_O;
assign MUX_SB_T1_WEST_SB_OUT_B1_I[1] = WIRE_SB_T0_SOUTH_SB_IN_B1_O;
assign MUX_SB_T1_WEST_SB_OUT_B1_I[0] = WIRE_SB_T4_NORTH_SB_IN_B1_O;
wire [5:0] MUX_SB_T1_WEST_SB_OUT_B1_valid_in;
assign MUX_SB_T1_WEST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T1_EAST_SB_IN_B1_valid_out,WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T4_NORTH_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T1_WEST_SB_OUT_B1 (
    .I(MUX_SB_T1_WEST_SB_OUT_B1_I),
    .O(MUX_SB_T1_WEST_SB_OUT_B1_O),
    .ready_in(SB_T1_WEST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T1_WEST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T1_WEST_SB_OUT_B1_valid_out),
    .S(SB_T1_WEST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T1_WEST_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1_I [5:0];
assign MUX_SB_T2_EAST_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T2_EAST_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T2_EAST_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T2_EAST_SB_OUT_B1_I[2] = WIRE_SB_T2_WEST_SB_IN_B1_O;
assign MUX_SB_T2_EAST_SB_OUT_B1_I[1] = WIRE_SB_T1_SOUTH_SB_IN_B1_O;
assign MUX_SB_T2_EAST_SB_OUT_B1_I[0] = WIRE_SB_T1_NORTH_SB_IN_B1_O;
wire [5:0] MUX_SB_T2_EAST_SB_OUT_B1_valid_in;
assign MUX_SB_T2_EAST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T2_WEST_SB_IN_B1_valid_out,WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T1_NORTH_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T2_EAST_SB_OUT_B1 (
    .I(MUX_SB_T2_EAST_SB_OUT_B1_I),
    .O(MUX_SB_T2_EAST_SB_OUT_B1_O),
    .ready_in(SB_T2_EAST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T2_EAST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T2_EAST_SB_OUT_B1_valid_out),
    .S(SB_T2_EAST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T2_EAST_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T2_NORTH_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T2_NORTH_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T2_NORTH_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T2_NORTH_SB_OUT_B1_I[2] = WIRE_SB_T3_WEST_SB_IN_B1_O;
assign MUX_SB_T2_NORTH_SB_OUT_B1_I[1] = WIRE_SB_T2_SOUTH_SB_IN_B1_O;
assign MUX_SB_T2_NORTH_SB_OUT_B1_I[0] = WIRE_SB_T3_EAST_SB_IN_B1_O;
wire [5:0] MUX_SB_T2_NORTH_SB_OUT_B1_valid_in;
assign MUX_SB_T2_NORTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T3_WEST_SB_IN_B1_valid_out,WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T3_EAST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T2_NORTH_SB_OUT_B1 (
    .I(MUX_SB_T2_NORTH_SB_OUT_B1_I),
    .O(MUX_SB_T2_NORTH_SB_OUT_B1_O),
    .ready_in(SB_T2_NORTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T2_NORTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T2_NORTH_SB_OUT_B1_valid_out),
    .S(SB_T2_NORTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[2] = WIRE_SB_T3_WEST_SB_IN_B1_O;
assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[1] = WIRE_SB_T2_NORTH_SB_IN_B1_O;
assign MUX_SB_T2_SOUTH_SB_OUT_B1_I[0] = WIRE_SB_T1_EAST_SB_IN_B1_O;
wire [5:0] MUX_SB_T2_SOUTH_SB_OUT_B1_valid_in;
assign MUX_SB_T2_SOUTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T3_WEST_SB_IN_B1_valid_out,WIRE_SB_T2_NORTH_SB_IN_B1_valid_out,WIRE_SB_T1_EAST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T2_SOUTH_SB_OUT_B1 (
    .I(MUX_SB_T2_SOUTH_SB_OUT_B1_I),
    .O(MUX_SB_T2_SOUTH_SB_OUT_B1_O),
    .ready_in(SB_T2_SOUTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T2_SOUTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T2_SOUTH_SB_OUT_B1_valid_out),
    .S(SB_T2_SOUTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1_I [5:0];
assign MUX_SB_T2_WEST_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T2_WEST_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T2_WEST_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T2_WEST_SB_OUT_B1_I[2] = WIRE_SB_T2_EAST_SB_IN_B1_O;
assign MUX_SB_T2_WEST_SB_OUT_B1_I[1] = WIRE_SB_T1_SOUTH_SB_IN_B1_O;
assign MUX_SB_T2_WEST_SB_OUT_B1_I[0] = WIRE_SB_T3_NORTH_SB_IN_B1_O;
wire [5:0] MUX_SB_T2_WEST_SB_OUT_B1_valid_in;
assign MUX_SB_T2_WEST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T2_EAST_SB_IN_B1_valid_out,WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T3_NORTH_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T2_WEST_SB_OUT_B1 (
    .I(MUX_SB_T2_WEST_SB_OUT_B1_I),
    .O(MUX_SB_T2_WEST_SB_OUT_B1_O),
    .ready_in(SB_T2_WEST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T2_WEST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T2_WEST_SB_OUT_B1_valid_out),
    .S(SB_T2_WEST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T2_WEST_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1_I [5:0];
assign MUX_SB_T3_EAST_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T3_EAST_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T3_EAST_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T3_EAST_SB_OUT_B1_I[2] = WIRE_SB_T3_WEST_SB_IN_B1_O;
assign MUX_SB_T3_EAST_SB_OUT_B1_I[1] = WIRE_SB_T2_NORTH_SB_IN_B1_O;
assign MUX_SB_T3_EAST_SB_OUT_B1_I[0] = WIRE_SB_T0_SOUTH_SB_IN_B1_O;
wire [5:0] MUX_SB_T3_EAST_SB_OUT_B1_valid_in;
assign MUX_SB_T3_EAST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T3_WEST_SB_IN_B1_valid_out,WIRE_SB_T2_NORTH_SB_IN_B1_valid_out,WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T3_EAST_SB_OUT_B1 (
    .I(MUX_SB_T3_EAST_SB_OUT_B1_I),
    .O(MUX_SB_T3_EAST_SB_OUT_B1_O),
    .ready_in(SB_T3_EAST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T3_EAST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T3_EAST_SB_OUT_B1_valid_out),
    .S(SB_T3_EAST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T3_EAST_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T3_NORTH_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T3_NORTH_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T3_NORTH_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T3_NORTH_SB_OUT_B1_I[2] = WIRE_SB_T3_SOUTH_SB_IN_B1_O;
assign MUX_SB_T3_NORTH_SB_OUT_B1_I[1] = WIRE_SB_T4_EAST_SB_IN_B1_O;
assign MUX_SB_T3_NORTH_SB_OUT_B1_I[0] = WIRE_SB_T2_WEST_SB_IN_B1_O;
wire [5:0] MUX_SB_T3_NORTH_SB_OUT_B1_valid_in;
assign MUX_SB_T3_NORTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T4_EAST_SB_IN_B1_valid_out,WIRE_SB_T2_WEST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T3_NORTH_SB_OUT_B1 (
    .I(MUX_SB_T3_NORTH_SB_OUT_B1_I),
    .O(MUX_SB_T3_NORTH_SB_OUT_B1_O),
    .ready_in(SB_T3_NORTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T3_NORTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T3_NORTH_SB_OUT_B1_valid_out),
    .S(SB_T3_NORTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[2] = WIRE_SB_T4_WEST_SB_IN_B1_O;
assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[1] = WIRE_SB_T3_NORTH_SB_IN_B1_O;
assign MUX_SB_T3_SOUTH_SB_OUT_B1_I[0] = WIRE_SB_T0_EAST_SB_IN_B1_O;
wire [5:0] MUX_SB_T3_SOUTH_SB_OUT_B1_valid_in;
assign MUX_SB_T3_SOUTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T4_WEST_SB_IN_B1_valid_out,WIRE_SB_T3_NORTH_SB_IN_B1_valid_out,WIRE_SB_T0_EAST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T3_SOUTH_SB_OUT_B1 (
    .I(MUX_SB_T3_SOUTH_SB_OUT_B1_I),
    .O(MUX_SB_T3_SOUTH_SB_OUT_B1_O),
    .ready_in(SB_T3_SOUTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T3_SOUTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T3_SOUTH_SB_OUT_B1_valid_out),
    .S(SB_T3_SOUTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1_I [5:0];
assign MUX_SB_T3_WEST_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T3_WEST_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T3_WEST_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T3_WEST_SB_OUT_B1_I[2] = WIRE_SB_T3_EAST_SB_IN_B1_O;
assign MUX_SB_T3_WEST_SB_OUT_B1_I[1] = WIRE_SB_T2_SOUTH_SB_IN_B1_O;
assign MUX_SB_T3_WEST_SB_OUT_B1_I[0] = WIRE_SB_T2_NORTH_SB_IN_B1_O;
wire [5:0] MUX_SB_T3_WEST_SB_OUT_B1_valid_in;
assign MUX_SB_T3_WEST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T3_EAST_SB_IN_B1_valid_out,WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T2_NORTH_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T3_WEST_SB_OUT_B1 (
    .I(MUX_SB_T3_WEST_SB_OUT_B1_I),
    .O(MUX_SB_T3_WEST_SB_OUT_B1_O),
    .ready_in(SB_T3_WEST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T3_WEST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T3_WEST_SB_OUT_B1_valid_out),
    .S(SB_T3_WEST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T3_WEST_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1_I [5:0];
assign MUX_SB_T4_EAST_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T4_EAST_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T4_EAST_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T4_EAST_SB_OUT_B1_I[2] = WIRE_SB_T4_WEST_SB_IN_B1_O;
assign MUX_SB_T4_EAST_SB_OUT_B1_I[1] = WIRE_SB_T4_SOUTH_SB_IN_B1_O;
assign MUX_SB_T4_EAST_SB_OUT_B1_I[0] = WIRE_SB_T3_NORTH_SB_IN_B1_O;
wire [5:0] MUX_SB_T4_EAST_SB_OUT_B1_valid_in;
assign MUX_SB_T4_EAST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T4_WEST_SB_IN_B1_valid_out,WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T3_NORTH_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T4_EAST_SB_OUT_B1 (
    .I(MUX_SB_T4_EAST_SB_OUT_B1_I),
    .O(MUX_SB_T4_EAST_SB_OUT_B1_O),
    .ready_in(SB_T4_EAST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T4_EAST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T4_EAST_SB_OUT_B1_valid_out),
    .S(SB_T4_EAST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T4_EAST_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T4_NORTH_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T4_NORTH_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T4_NORTH_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T4_NORTH_SB_OUT_B1_I[2] = WIRE_SB_T4_SOUTH_SB_IN_B1_O;
assign MUX_SB_T4_NORTH_SB_OUT_B1_I[1] = WIRE_SB_T0_EAST_SB_IN_B1_O;
assign MUX_SB_T4_NORTH_SB_OUT_B1_I[0] = WIRE_SB_T1_WEST_SB_IN_B1_O;
wire [5:0] MUX_SB_T4_NORTH_SB_OUT_B1_valid_in;
assign MUX_SB_T4_NORTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T0_EAST_SB_IN_B1_valid_out,WIRE_SB_T1_WEST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T4_NORTH_SB_OUT_B1 (
    .I(MUX_SB_T4_NORTH_SB_OUT_B1_I),
    .O(MUX_SB_T4_NORTH_SB_OUT_B1_O),
    .ready_in(SB_T4_NORTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T4_NORTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T4_NORTH_SB_OUT_B1_valid_out),
    .S(SB_T4_NORTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1_I [5:0];
assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[2] = WIRE_SB_T4_NORTH_SB_IN_B1_O;
assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[1] = WIRE_SB_T4_EAST_SB_IN_B1_O;
assign MUX_SB_T4_SOUTH_SB_OUT_B1_I[0] = WIRE_SB_T0_WEST_SB_IN_B1_O;
wire [5:0] MUX_SB_T4_SOUTH_SB_OUT_B1_valid_in;
assign MUX_SB_T4_SOUTH_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T4_NORTH_SB_IN_B1_valid_out,WIRE_SB_T4_EAST_SB_IN_B1_valid_out,WIRE_SB_T0_WEST_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T4_SOUTH_SB_OUT_B1 (
    .I(MUX_SB_T4_SOUTH_SB_OUT_B1_I),
    .O(MUX_SB_T4_SOUTH_SB_OUT_B1_O),
    .ready_in(SB_T4_SOUTH_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T4_SOUTH_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T4_SOUTH_SB_OUT_B1_valid_out),
    .S(SB_T4_SOUTH_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel)
);
wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1_I [5:0];
assign MUX_SB_T4_WEST_SB_OUT_B1_I[5] = MEM_output_width_1_num_2;
assign MUX_SB_T4_WEST_SB_OUT_B1_I[4] = MEM_output_width_1_num_1;
assign MUX_SB_T4_WEST_SB_OUT_B1_I[3] = MEM_output_width_1_num_0;
assign MUX_SB_T4_WEST_SB_OUT_B1_I[2] = WIRE_SB_T4_EAST_SB_IN_B1_O;
assign MUX_SB_T4_WEST_SB_OUT_B1_I[1] = WIRE_SB_T3_SOUTH_SB_IN_B1_O;
assign MUX_SB_T4_WEST_SB_OUT_B1_I[0] = WIRE_SB_T1_NORTH_SB_IN_B1_O;
wire [5:0] MUX_SB_T4_WEST_SB_OUT_B1_valid_in;
assign MUX_SB_T4_WEST_SB_OUT_B1_valid_in = {MEM_output_width_1_num_2_valid,MEM_output_width_1_num_1_valid,MEM_output_width_1_num_0_valid,WIRE_SB_T4_EAST_SB_IN_B1_valid_out,WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out,WIRE_SB_T1_NORTH_SB_IN_B1_valid_out};
mux_aoi_ready_valid_6_1 MUX_SB_T4_WEST_SB_OUT_B1 (
    .I(MUX_SB_T4_WEST_SB_OUT_B1_I),
    .O(MUX_SB_T4_WEST_SB_OUT_B1_O),
    .ready_in(SB_T4_WEST_SB_OUT_B1_FANOUT_O[0]),
    .ready_out(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
    .valid_in(MUX_SB_T4_WEST_SB_OUT_B1_valid_in),
    .valid_out(MUX_SB_T4_WEST_SB_OUT_B1_valid_out),
    .S(SB_T4_WEST_SB_OUT_B1_sel_value_O),
    .out_sel(MUX_SB_T4_WEST_SB_OUT_B1_out_sel)
);
SplitFifo_1 REG_T0_EAST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T0_EAST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T0_EAST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T0_EAST_B1_fifo_value_O[0]),
    .end_fifo(REG_T0_EAST_B1_end_value_O[0]),
    .data_in(MUX_SB_T0_EAST_SB_OUT_B1_O),
    .ready1(RMUX_T0_EAST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T0_EAST_SB_OUT_B1_valid_out),
    .data_out(REG_T0_EAST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T0_EAST_B1_start_value_O[0]),
    .clk_en(and1_inst2_out[0])
);
SliceWrapper_32_0_1 REG_T0_EAST_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T0_EAST_B1_end_value_O)
);
SliceWrapper_32_1_2 REG_T0_EAST_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T0_EAST_B1_fifo_value_O)
);
SliceWrapper_32_2_3 REG_T0_EAST_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T0_EAST_B1_start_value_O)
);
SplitFifo_1 REG_T0_NORTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T0_NORTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T0_NORTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T0_NORTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T0_NORTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T0_NORTH_SB_OUT_B1_O),
    .ready1(RMUX_T0_NORTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T0_NORTH_SB_OUT_B1_valid_out),
    .data_out(REG_T0_NORTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T0_NORTH_B1_start_value_O[0]),
    .clk_en(and1_inst0_out[0])
);
SliceWrapper_32_3_4 REG_T0_NORTH_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T0_NORTH_B1_end_value_O)
);
SliceWrapper_32_4_5 REG_T0_NORTH_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T0_NORTH_B1_fifo_value_O)
);
SliceWrapper_32_5_6 REG_T0_NORTH_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T0_NORTH_B1_start_value_O)
);
SplitFifo_1 REG_T0_SOUTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T0_SOUTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T0_SOUTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T0_SOUTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T0_SOUTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T0_SOUTH_SB_OUT_B1_O),
    .ready1(RMUX_T0_SOUTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T0_SOUTH_SB_OUT_B1_valid_out),
    .data_out(REG_T0_SOUTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T0_SOUTH_B1_start_value_O[0]),
    .clk_en(and1_inst1_out[0])
);
SliceWrapper_32_6_7 REG_T0_SOUTH_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T0_SOUTH_B1_end_value_O)
);
SliceWrapper_32_7_8 REG_T0_SOUTH_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T0_SOUTH_B1_fifo_value_O)
);
SliceWrapper_32_8_9 REG_T0_SOUTH_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T0_SOUTH_B1_start_value_O)
);
SplitFifo_1 REG_T0_WEST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T0_WEST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T0_WEST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T0_WEST_B1_fifo_value_O[0]),
    .end_fifo(REG_T0_WEST_B1_end_value_O[0]),
    .data_in(MUX_SB_T0_WEST_SB_OUT_B1_O),
    .ready1(RMUX_T0_WEST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T0_WEST_SB_OUT_B1_valid_out),
    .data_out(REG_T0_WEST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T0_WEST_B1_start_value_O[0]),
    .clk_en(and1_inst3_out[0])
);
SliceWrapper_32_9_10 REG_T0_WEST_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T0_WEST_B1_end_value_O)
);
SliceWrapper_32_10_11 REG_T0_WEST_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T0_WEST_B1_fifo_value_O)
);
SliceWrapper_32_11_12 REG_T0_WEST_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T0_WEST_B1_start_value_O)
);
SplitFifo_1 REG_T1_EAST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T1_EAST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T1_EAST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T1_EAST_B1_fifo_value_O[0]),
    .end_fifo(REG_T1_EAST_B1_end_value_O[0]),
    .data_in(MUX_SB_T1_EAST_SB_OUT_B1_O),
    .ready1(RMUX_T1_EAST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T1_EAST_SB_OUT_B1_valid_out),
    .data_out(REG_T1_EAST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T1_EAST_B1_start_value_O[0]),
    .clk_en(and1_inst6_out[0])
);
SliceWrapper_32_12_13 REG_T1_EAST_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T1_EAST_B1_end_value_O)
);
SliceWrapper_32_13_14 REG_T1_EAST_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T1_EAST_B1_fifo_value_O)
);
SliceWrapper_32_14_15 REG_T1_EAST_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T1_EAST_B1_start_value_O)
);
SplitFifo_1 REG_T1_NORTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T1_NORTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T1_NORTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T1_NORTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T1_NORTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T1_NORTH_SB_OUT_B1_O),
    .ready1(RMUX_T1_NORTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T1_NORTH_SB_OUT_B1_valid_out),
    .data_out(REG_T1_NORTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T1_NORTH_B1_start_value_O[0]),
    .clk_en(and1_inst4_out[0])
);
SliceWrapper_32_15_16 REG_T1_NORTH_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T1_NORTH_B1_end_value_O)
);
SliceWrapper_32_16_17 REG_T1_NORTH_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T1_NORTH_B1_fifo_value_O)
);
SliceWrapper_32_17_18 REG_T1_NORTH_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T1_NORTH_B1_start_value_O)
);
SplitFifo_1 REG_T1_SOUTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T1_SOUTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T1_SOUTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T1_SOUTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T1_SOUTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T1_SOUTH_SB_OUT_B1_O),
    .ready1(RMUX_T1_SOUTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T1_SOUTH_SB_OUT_B1_valid_out),
    .data_out(REG_T1_SOUTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T1_SOUTH_B1_start_value_O[0]),
    .clk_en(and1_inst5_out[0])
);
SliceWrapper_32_18_19 REG_T1_SOUTH_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T1_SOUTH_B1_end_value_O)
);
SliceWrapper_32_19_20 REG_T1_SOUTH_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T1_SOUTH_B1_fifo_value_O)
);
SliceWrapper_32_20_21 REG_T1_SOUTH_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T1_SOUTH_B1_start_value_O)
);
SplitFifo_1 REG_T1_WEST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T1_WEST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T1_WEST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T1_WEST_B1_fifo_value_O[0]),
    .end_fifo(REG_T1_WEST_B1_end_value_O[0]),
    .data_in(MUX_SB_T1_WEST_SB_OUT_B1_O),
    .ready1(RMUX_T1_WEST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T1_WEST_SB_OUT_B1_valid_out),
    .data_out(REG_T1_WEST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T1_WEST_B1_start_value_O[0]),
    .clk_en(and1_inst7_out[0])
);
SliceWrapper_32_21_22 REG_T1_WEST_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T1_WEST_B1_end_value_O)
);
SliceWrapper_32_22_23 REG_T1_WEST_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T1_WEST_B1_fifo_value_O)
);
SliceWrapper_32_23_24 REG_T1_WEST_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T1_WEST_B1_start_value_O)
);
SplitFifo_1 REG_T2_EAST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T2_EAST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T2_EAST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T2_EAST_B1_fifo_value_O[0]),
    .end_fifo(REG_T2_EAST_B1_end_value_O[0]),
    .data_in(MUX_SB_T2_EAST_SB_OUT_B1_O),
    .ready1(RMUX_T2_EAST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T2_EAST_SB_OUT_B1_valid_out),
    .data_out(REG_T2_EAST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T2_EAST_B1_start_value_O[0]),
    .clk_en(and1_inst10_out[0])
);
SliceWrapper_32_24_25 REG_T2_EAST_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T2_EAST_B1_end_value_O)
);
SliceWrapper_32_25_26 REG_T2_EAST_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T2_EAST_B1_fifo_value_O)
);
SliceWrapper_32_26_27 REG_T2_EAST_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T2_EAST_B1_start_value_O)
);
SplitFifo_1 REG_T2_NORTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T2_NORTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T2_NORTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T2_NORTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T2_NORTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T2_NORTH_SB_OUT_B1_O),
    .ready1(RMUX_T2_NORTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T2_NORTH_SB_OUT_B1_valid_out),
    .data_out(REG_T2_NORTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T2_NORTH_B1_start_value_O[0]),
    .clk_en(and1_inst8_out[0])
);
SliceWrapper_32_27_28 REG_T2_NORTH_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T2_NORTH_B1_end_value_O)
);
SliceWrapper_32_28_29 REG_T2_NORTH_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T2_NORTH_B1_fifo_value_O)
);
SliceWrapper_32_29_30 REG_T2_NORTH_B1_start_value (
    .I(config_reg_0_O),
    .O(REG_T2_NORTH_B1_start_value_O)
);
SplitFifo_1 REG_T2_SOUTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T2_SOUTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T2_SOUTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T2_SOUTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T2_SOUTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T2_SOUTH_SB_OUT_B1_O),
    .ready1(RMUX_T2_SOUTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T2_SOUTH_SB_OUT_B1_valid_out),
    .data_out(REG_T2_SOUTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T2_SOUTH_B1_start_value_O[0]),
    .clk_en(and1_inst9_out[0])
);
SliceWrapper_32_30_31 REG_T2_SOUTH_B1_end_value (
    .I(config_reg_0_O),
    .O(REG_T2_SOUTH_B1_end_value_O)
);
SliceWrapper_32_31_32 REG_T2_SOUTH_B1_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T2_SOUTH_B1_fifo_value_O)
);
SliceWrapper_32_0_1 REG_T2_SOUTH_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T2_SOUTH_B1_start_value_O)
);
SplitFifo_1 REG_T2_WEST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T2_WEST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T2_WEST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T2_WEST_B1_fifo_value_O[0]),
    .end_fifo(REG_T2_WEST_B1_end_value_O[0]),
    .data_in(MUX_SB_T2_WEST_SB_OUT_B1_O),
    .ready1(RMUX_T2_WEST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T2_WEST_SB_OUT_B1_valid_out),
    .data_out(REG_T2_WEST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T2_WEST_B1_start_value_O[0]),
    .clk_en(and1_inst11_out[0])
);
SliceWrapper_32_1_2 REG_T2_WEST_B1_end_value (
    .I(config_reg_1_O),
    .O(REG_T2_WEST_B1_end_value_O)
);
SliceWrapper_32_2_3 REG_T2_WEST_B1_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T2_WEST_B1_fifo_value_O)
);
SliceWrapper_32_3_4 REG_T2_WEST_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T2_WEST_B1_start_value_O)
);
SplitFifo_1 REG_T3_EAST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T3_EAST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T3_EAST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T3_EAST_B1_fifo_value_O[0]),
    .end_fifo(REG_T3_EAST_B1_end_value_O[0]),
    .data_in(MUX_SB_T3_EAST_SB_OUT_B1_O),
    .ready1(RMUX_T3_EAST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T3_EAST_SB_OUT_B1_valid_out),
    .data_out(REG_T3_EAST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T3_EAST_B1_start_value_O[0]),
    .clk_en(and1_inst14_out[0])
);
SliceWrapper_32_4_5 REG_T3_EAST_B1_end_value (
    .I(config_reg_1_O),
    .O(REG_T3_EAST_B1_end_value_O)
);
SliceWrapper_32_5_6 REG_T3_EAST_B1_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T3_EAST_B1_fifo_value_O)
);
SliceWrapper_32_6_7 REG_T3_EAST_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T3_EAST_B1_start_value_O)
);
SplitFifo_1 REG_T3_NORTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T3_NORTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T3_NORTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T3_NORTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T3_NORTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T3_NORTH_SB_OUT_B1_O),
    .ready1(RMUX_T3_NORTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T3_NORTH_SB_OUT_B1_valid_out),
    .data_out(REG_T3_NORTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T3_NORTH_B1_start_value_O[0]),
    .clk_en(and1_inst12_out[0])
);
SliceWrapper_32_7_8 REG_T3_NORTH_B1_end_value (
    .I(config_reg_1_O),
    .O(REG_T3_NORTH_B1_end_value_O)
);
SliceWrapper_32_8_9 REG_T3_NORTH_B1_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T3_NORTH_B1_fifo_value_O)
);
SliceWrapper_32_9_10 REG_T3_NORTH_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T3_NORTH_B1_start_value_O)
);
SplitFifo_1 REG_T3_SOUTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T3_SOUTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T3_SOUTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T3_SOUTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T3_SOUTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T3_SOUTH_SB_OUT_B1_O),
    .ready1(RMUX_T3_SOUTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T3_SOUTH_SB_OUT_B1_valid_out),
    .data_out(REG_T3_SOUTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T3_SOUTH_B1_start_value_O[0]),
    .clk_en(and1_inst13_out[0])
);
SliceWrapper_32_10_11 REG_T3_SOUTH_B1_end_value (
    .I(config_reg_1_O),
    .O(REG_T3_SOUTH_B1_end_value_O)
);
SliceWrapper_32_11_12 REG_T3_SOUTH_B1_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T3_SOUTH_B1_fifo_value_O)
);
SliceWrapper_32_12_13 REG_T3_SOUTH_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T3_SOUTH_B1_start_value_O)
);
SplitFifo_1 REG_T3_WEST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T3_WEST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T3_WEST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T3_WEST_B1_fifo_value_O[0]),
    .end_fifo(REG_T3_WEST_B1_end_value_O[0]),
    .data_in(MUX_SB_T3_WEST_SB_OUT_B1_O),
    .ready1(RMUX_T3_WEST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T3_WEST_SB_OUT_B1_valid_out),
    .data_out(REG_T3_WEST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T3_WEST_B1_start_value_O[0]),
    .clk_en(and1_inst15_out[0])
);
SliceWrapper_32_13_14 REG_T3_WEST_B1_end_value (
    .I(config_reg_1_O),
    .O(REG_T3_WEST_B1_end_value_O)
);
SliceWrapper_32_14_15 REG_T3_WEST_B1_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T3_WEST_B1_fifo_value_O)
);
SliceWrapper_32_15_16 REG_T3_WEST_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T3_WEST_B1_start_value_O)
);
SplitFifo_1 REG_T4_EAST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T4_EAST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T4_EAST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T4_EAST_B1_fifo_value_O[0]),
    .end_fifo(REG_T4_EAST_B1_end_value_O[0]),
    .data_in(MUX_SB_T4_EAST_SB_OUT_B1_O),
    .ready1(RMUX_T4_EAST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T4_EAST_SB_OUT_B1_valid_out),
    .data_out(REG_T4_EAST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T4_EAST_B1_start_value_O[0]),
    .clk_en(and1_inst18_out[0])
);
SliceWrapper_32_16_17 REG_T4_EAST_B1_end_value (
    .I(config_reg_1_O),
    .O(REG_T4_EAST_B1_end_value_O)
);
SliceWrapper_32_17_18 REG_T4_EAST_B1_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T4_EAST_B1_fifo_value_O)
);
SliceWrapper_32_18_19 REG_T4_EAST_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T4_EAST_B1_start_value_O)
);
SplitFifo_1 REG_T4_NORTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T4_NORTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T4_NORTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T4_NORTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T4_NORTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T4_NORTH_SB_OUT_B1_O),
    .ready1(RMUX_T4_NORTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T4_NORTH_SB_OUT_B1_valid_out),
    .data_out(REG_T4_NORTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T4_NORTH_B1_start_value_O[0]),
    .clk_en(and1_inst16_out[0])
);
SliceWrapper_32_19_20 REG_T4_NORTH_B1_end_value (
    .I(config_reg_1_O),
    .O(REG_T4_NORTH_B1_end_value_O)
);
SliceWrapper_32_20_21 REG_T4_NORTH_B1_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T4_NORTH_B1_fifo_value_O)
);
SliceWrapper_32_21_22 REG_T4_NORTH_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T4_NORTH_B1_start_value_O)
);
SplitFifo_1 REG_T4_SOUTH_B1$SplitFifo_1_inst0 (
    .ready0(REG_T4_SOUTH_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T4_SOUTH_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T4_SOUTH_B1_fifo_value_O[0]),
    .end_fifo(REG_T4_SOUTH_B1_end_value_O[0]),
    .data_in(MUX_SB_T4_SOUTH_SB_OUT_B1_O),
    .ready1(RMUX_T4_SOUTH_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T4_SOUTH_SB_OUT_B1_valid_out),
    .data_out(REG_T4_SOUTH_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T4_SOUTH_B1_start_value_O[0]),
    .clk_en(and1_inst17_out[0])
);
SliceWrapper_32_22_23 REG_T4_SOUTH_B1_end_value (
    .I(config_reg_1_O),
    .O(REG_T4_SOUTH_B1_end_value_O)
);
SliceWrapper_32_23_24 REG_T4_SOUTH_B1_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T4_SOUTH_B1_fifo_value_O)
);
SliceWrapper_32_24_25 REG_T4_SOUTH_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T4_SOUTH_B1_start_value_O)
);
SplitFifo_1 REG_T4_WEST_B1$SplitFifo_1_inst0 (
    .ready0(REG_T4_WEST_B1$SplitFifo_1_inst0_ready0),
    .rst(reset),
    .valid1(REG_T4_WEST_B1$SplitFifo_1_inst0_valid1),
    .fifo_en(REG_T4_WEST_B1_fifo_value_O[0]),
    .end_fifo(REG_T4_WEST_B1_end_value_O[0]),
    .data_in(MUX_SB_T4_WEST_SB_OUT_B1_O),
    .ready1(RMUX_T4_WEST_B1_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T4_WEST_SB_OUT_B1_valid_out),
    .data_out(REG_T4_WEST_B1$SplitFifo_1_inst0_data_out),
    .start_fifo(REG_T4_WEST_B1_start_value_O[0]),
    .clk_en(and1_inst19_out[0])
);
SliceWrapper_32_25_26 REG_T4_WEST_B1_end_value (
    .I(config_reg_1_O),
    .O(REG_T4_WEST_B1_end_value_O)
);
SliceWrapper_32_26_27 REG_T4_WEST_B1_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T4_WEST_B1_fifo_value_O)
);
SliceWrapper_32_27_28 REG_T4_WEST_B1_start_value (
    .I(config_reg_1_O),
    .O(REG_T4_WEST_B1_start_value_O)
);
wire [0:0] RMUX_T0_EAST_B1_I [1:0];
assign RMUX_T0_EAST_B1_I[1] = REG_T0_EAST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T0_EAST_B1_I[0] = MUX_SB_T0_EAST_SB_OUT_B1_O;
wire [1:0] RMUX_T0_EAST_B1_valid_in;
assign RMUX_T0_EAST_B1_valid_in = {REG_T0_EAST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T0_EAST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T0_EAST_B1 (
    .I(RMUX_T0_EAST_B1_I),
    .O(RMUX_T0_EAST_B1_O),
    .ready_in(SB_T0_EAST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T0_EAST_B1_ready_out),
    .valid_in(RMUX_T0_EAST_B1_valid_in),
    .valid_out(RMUX_T0_EAST_B1_valid_out),
    .S(RMUX_T0_EAST_B1_sel_value_O),
    .out_sel(RMUX_T0_EAST_B1_out_sel)
);
SliceWrapper_32_28_29 RMUX_T0_EAST_B1_sel_value (
    .I(config_reg_1_O),
    .O(RMUX_T0_EAST_B1_sel_value_O)
);
wire [0:0] RMUX_T0_NORTH_B1_I [1:0];
assign RMUX_T0_NORTH_B1_I[1] = REG_T0_NORTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T0_NORTH_B1_I[0] = MUX_SB_T0_NORTH_SB_OUT_B1_O;
wire [1:0] RMUX_T0_NORTH_B1_valid_in;
assign RMUX_T0_NORTH_B1_valid_in = {REG_T0_NORTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T0_NORTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T0_NORTH_B1 (
    .I(RMUX_T0_NORTH_B1_I),
    .O(RMUX_T0_NORTH_B1_O),
    .ready_in(SB_T0_NORTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T0_NORTH_B1_ready_out),
    .valid_in(RMUX_T0_NORTH_B1_valid_in),
    .valid_out(RMUX_T0_NORTH_B1_valid_out),
    .S(RMUX_T0_NORTH_B1_sel_value_O),
    .out_sel(RMUX_T0_NORTH_B1_out_sel)
);
SliceWrapper_32_29_30 RMUX_T0_NORTH_B1_sel_value (
    .I(config_reg_1_O),
    .O(RMUX_T0_NORTH_B1_sel_value_O)
);
wire [0:0] RMUX_T0_SOUTH_B1_I [1:0];
assign RMUX_T0_SOUTH_B1_I[1] = REG_T0_SOUTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T0_SOUTH_B1_I[0] = MUX_SB_T0_SOUTH_SB_OUT_B1_O;
wire [1:0] RMUX_T0_SOUTH_B1_valid_in;
assign RMUX_T0_SOUTH_B1_valid_in = {REG_T0_SOUTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T0_SOUTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T0_SOUTH_B1 (
    .I(RMUX_T0_SOUTH_B1_I),
    .O(RMUX_T0_SOUTH_B1_O),
    .ready_in(SB_T0_SOUTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T0_SOUTH_B1_ready_out),
    .valid_in(RMUX_T0_SOUTH_B1_valid_in),
    .valid_out(RMUX_T0_SOUTH_B1_valid_out),
    .S(RMUX_T0_SOUTH_B1_sel_value_O),
    .out_sel(RMUX_T0_SOUTH_B1_out_sel)
);
SliceWrapper_32_30_31 RMUX_T0_SOUTH_B1_sel_value (
    .I(config_reg_1_O),
    .O(RMUX_T0_SOUTH_B1_sel_value_O)
);
wire [0:0] RMUX_T0_WEST_B1_I [1:0];
assign RMUX_T0_WEST_B1_I[1] = REG_T0_WEST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T0_WEST_B1_I[0] = MUX_SB_T0_WEST_SB_OUT_B1_O;
wire [1:0] RMUX_T0_WEST_B1_valid_in;
assign RMUX_T0_WEST_B1_valid_in = {REG_T0_WEST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T0_WEST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T0_WEST_B1 (
    .I(RMUX_T0_WEST_B1_I),
    .O(RMUX_T0_WEST_B1_O),
    .ready_in(SB_T0_WEST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T0_WEST_B1_ready_out),
    .valid_in(RMUX_T0_WEST_B1_valid_in),
    .valid_out(RMUX_T0_WEST_B1_valid_out),
    .S(RMUX_T0_WEST_B1_sel_value_O),
    .out_sel(RMUX_T0_WEST_B1_out_sel)
);
SliceWrapper_32_31_32 RMUX_T0_WEST_B1_sel_value (
    .I(config_reg_1_O),
    .O(RMUX_T0_WEST_B1_sel_value_O)
);
wire [0:0] RMUX_T1_EAST_B1_I [1:0];
assign RMUX_T1_EAST_B1_I[1] = REG_T1_EAST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T1_EAST_B1_I[0] = MUX_SB_T1_EAST_SB_OUT_B1_O;
wire [1:0] RMUX_T1_EAST_B1_valid_in;
assign RMUX_T1_EAST_B1_valid_in = {REG_T1_EAST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T1_EAST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T1_EAST_B1 (
    .I(RMUX_T1_EAST_B1_I),
    .O(RMUX_T1_EAST_B1_O),
    .ready_in(SB_T1_EAST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T1_EAST_B1_ready_out),
    .valid_in(RMUX_T1_EAST_B1_valid_in),
    .valid_out(RMUX_T1_EAST_B1_valid_out),
    .S(RMUX_T1_EAST_B1_sel_value_O),
    .out_sel(RMUX_T1_EAST_B1_out_sel)
);
SliceWrapper_32_0_1 RMUX_T1_EAST_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T1_EAST_B1_sel_value_O)
);
wire [0:0] RMUX_T1_NORTH_B1_I [1:0];
assign RMUX_T1_NORTH_B1_I[1] = REG_T1_NORTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T1_NORTH_B1_I[0] = MUX_SB_T1_NORTH_SB_OUT_B1_O;
wire [1:0] RMUX_T1_NORTH_B1_valid_in;
assign RMUX_T1_NORTH_B1_valid_in = {REG_T1_NORTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T1_NORTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T1_NORTH_B1 (
    .I(RMUX_T1_NORTH_B1_I),
    .O(RMUX_T1_NORTH_B1_O),
    .ready_in(SB_T1_NORTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T1_NORTH_B1_ready_out),
    .valid_in(RMUX_T1_NORTH_B1_valid_in),
    .valid_out(RMUX_T1_NORTH_B1_valid_out),
    .S(RMUX_T1_NORTH_B1_sel_value_O),
    .out_sel(RMUX_T1_NORTH_B1_out_sel)
);
SliceWrapper_32_1_2 RMUX_T1_NORTH_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T1_NORTH_B1_sel_value_O)
);
wire [0:0] RMUX_T1_SOUTH_B1_I [1:0];
assign RMUX_T1_SOUTH_B1_I[1] = REG_T1_SOUTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T1_SOUTH_B1_I[0] = MUX_SB_T1_SOUTH_SB_OUT_B1_O;
wire [1:0] RMUX_T1_SOUTH_B1_valid_in;
assign RMUX_T1_SOUTH_B1_valid_in = {REG_T1_SOUTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T1_SOUTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T1_SOUTH_B1 (
    .I(RMUX_T1_SOUTH_B1_I),
    .O(RMUX_T1_SOUTH_B1_O),
    .ready_in(SB_T1_SOUTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T1_SOUTH_B1_ready_out),
    .valid_in(RMUX_T1_SOUTH_B1_valid_in),
    .valid_out(RMUX_T1_SOUTH_B1_valid_out),
    .S(RMUX_T1_SOUTH_B1_sel_value_O),
    .out_sel(RMUX_T1_SOUTH_B1_out_sel)
);
SliceWrapper_32_2_3 RMUX_T1_SOUTH_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T1_SOUTH_B1_sel_value_O)
);
wire [0:0] RMUX_T1_WEST_B1_I [1:0];
assign RMUX_T1_WEST_B1_I[1] = REG_T1_WEST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T1_WEST_B1_I[0] = MUX_SB_T1_WEST_SB_OUT_B1_O;
wire [1:0] RMUX_T1_WEST_B1_valid_in;
assign RMUX_T1_WEST_B1_valid_in = {REG_T1_WEST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T1_WEST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T1_WEST_B1 (
    .I(RMUX_T1_WEST_B1_I),
    .O(RMUX_T1_WEST_B1_O),
    .ready_in(SB_T1_WEST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T1_WEST_B1_ready_out),
    .valid_in(RMUX_T1_WEST_B1_valid_in),
    .valid_out(RMUX_T1_WEST_B1_valid_out),
    .S(RMUX_T1_WEST_B1_sel_value_O),
    .out_sel(RMUX_T1_WEST_B1_out_sel)
);
SliceWrapper_32_3_4 RMUX_T1_WEST_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T1_WEST_B1_sel_value_O)
);
wire [0:0] RMUX_T2_EAST_B1_I [1:0];
assign RMUX_T2_EAST_B1_I[1] = REG_T2_EAST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T2_EAST_B1_I[0] = MUX_SB_T2_EAST_SB_OUT_B1_O;
wire [1:0] RMUX_T2_EAST_B1_valid_in;
assign RMUX_T2_EAST_B1_valid_in = {REG_T2_EAST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T2_EAST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T2_EAST_B1 (
    .I(RMUX_T2_EAST_B1_I),
    .O(RMUX_T2_EAST_B1_O),
    .ready_in(SB_T2_EAST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T2_EAST_B1_ready_out),
    .valid_in(RMUX_T2_EAST_B1_valid_in),
    .valid_out(RMUX_T2_EAST_B1_valid_out),
    .S(RMUX_T2_EAST_B1_sel_value_O),
    .out_sel(RMUX_T2_EAST_B1_out_sel)
);
SliceWrapper_32_4_5 RMUX_T2_EAST_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T2_EAST_B1_sel_value_O)
);
wire [0:0] RMUX_T2_NORTH_B1_I [1:0];
assign RMUX_T2_NORTH_B1_I[1] = REG_T2_NORTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T2_NORTH_B1_I[0] = MUX_SB_T2_NORTH_SB_OUT_B1_O;
wire [1:0] RMUX_T2_NORTH_B1_valid_in;
assign RMUX_T2_NORTH_B1_valid_in = {REG_T2_NORTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T2_NORTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T2_NORTH_B1 (
    .I(RMUX_T2_NORTH_B1_I),
    .O(RMUX_T2_NORTH_B1_O),
    .ready_in(SB_T2_NORTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T2_NORTH_B1_ready_out),
    .valid_in(RMUX_T2_NORTH_B1_valid_in),
    .valid_out(RMUX_T2_NORTH_B1_valid_out),
    .S(RMUX_T2_NORTH_B1_sel_value_O),
    .out_sel(RMUX_T2_NORTH_B1_out_sel)
);
SliceWrapper_32_5_6 RMUX_T2_NORTH_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T2_NORTH_B1_sel_value_O)
);
wire [0:0] RMUX_T2_SOUTH_B1_I [1:0];
assign RMUX_T2_SOUTH_B1_I[1] = REG_T2_SOUTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T2_SOUTH_B1_I[0] = MUX_SB_T2_SOUTH_SB_OUT_B1_O;
wire [1:0] RMUX_T2_SOUTH_B1_valid_in;
assign RMUX_T2_SOUTH_B1_valid_in = {REG_T2_SOUTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T2_SOUTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T2_SOUTH_B1 (
    .I(RMUX_T2_SOUTH_B1_I),
    .O(RMUX_T2_SOUTH_B1_O),
    .ready_in(SB_T2_SOUTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T2_SOUTH_B1_ready_out),
    .valid_in(RMUX_T2_SOUTH_B1_valid_in),
    .valid_out(RMUX_T2_SOUTH_B1_valid_out),
    .S(RMUX_T2_SOUTH_B1_sel_value_O),
    .out_sel(RMUX_T2_SOUTH_B1_out_sel)
);
SliceWrapper_32_6_7 RMUX_T2_SOUTH_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T2_SOUTH_B1_sel_value_O)
);
wire [0:0] RMUX_T2_WEST_B1_I [1:0];
assign RMUX_T2_WEST_B1_I[1] = REG_T2_WEST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T2_WEST_B1_I[0] = MUX_SB_T2_WEST_SB_OUT_B1_O;
wire [1:0] RMUX_T2_WEST_B1_valid_in;
assign RMUX_T2_WEST_B1_valid_in = {REG_T2_WEST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T2_WEST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T2_WEST_B1 (
    .I(RMUX_T2_WEST_B1_I),
    .O(RMUX_T2_WEST_B1_O),
    .ready_in(SB_T2_WEST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T2_WEST_B1_ready_out),
    .valid_in(RMUX_T2_WEST_B1_valid_in),
    .valid_out(RMUX_T2_WEST_B1_valid_out),
    .S(RMUX_T2_WEST_B1_sel_value_O),
    .out_sel(RMUX_T2_WEST_B1_out_sel)
);
SliceWrapper_32_7_8 RMUX_T2_WEST_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T2_WEST_B1_sel_value_O)
);
wire [0:0] RMUX_T3_EAST_B1_I [1:0];
assign RMUX_T3_EAST_B1_I[1] = REG_T3_EAST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T3_EAST_B1_I[0] = MUX_SB_T3_EAST_SB_OUT_B1_O;
wire [1:0] RMUX_T3_EAST_B1_valid_in;
assign RMUX_T3_EAST_B1_valid_in = {REG_T3_EAST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T3_EAST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T3_EAST_B1 (
    .I(RMUX_T3_EAST_B1_I),
    .O(RMUX_T3_EAST_B1_O),
    .ready_in(SB_T3_EAST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T3_EAST_B1_ready_out),
    .valid_in(RMUX_T3_EAST_B1_valid_in),
    .valid_out(RMUX_T3_EAST_B1_valid_out),
    .S(RMUX_T3_EAST_B1_sel_value_O),
    .out_sel(RMUX_T3_EAST_B1_out_sel)
);
SliceWrapper_32_8_9 RMUX_T3_EAST_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T3_EAST_B1_sel_value_O)
);
wire [0:0] RMUX_T3_NORTH_B1_I [1:0];
assign RMUX_T3_NORTH_B1_I[1] = REG_T3_NORTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T3_NORTH_B1_I[0] = MUX_SB_T3_NORTH_SB_OUT_B1_O;
wire [1:0] RMUX_T3_NORTH_B1_valid_in;
assign RMUX_T3_NORTH_B1_valid_in = {REG_T3_NORTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T3_NORTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T3_NORTH_B1 (
    .I(RMUX_T3_NORTH_B1_I),
    .O(RMUX_T3_NORTH_B1_O),
    .ready_in(SB_T3_NORTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T3_NORTH_B1_ready_out),
    .valid_in(RMUX_T3_NORTH_B1_valid_in),
    .valid_out(RMUX_T3_NORTH_B1_valid_out),
    .S(RMUX_T3_NORTH_B1_sel_value_O),
    .out_sel(RMUX_T3_NORTH_B1_out_sel)
);
SliceWrapper_32_9_10 RMUX_T3_NORTH_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T3_NORTH_B1_sel_value_O)
);
wire [0:0] RMUX_T3_SOUTH_B1_I [1:0];
assign RMUX_T3_SOUTH_B1_I[1] = REG_T3_SOUTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T3_SOUTH_B1_I[0] = MUX_SB_T3_SOUTH_SB_OUT_B1_O;
wire [1:0] RMUX_T3_SOUTH_B1_valid_in;
assign RMUX_T3_SOUTH_B1_valid_in = {REG_T3_SOUTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T3_SOUTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T3_SOUTH_B1 (
    .I(RMUX_T3_SOUTH_B1_I),
    .O(RMUX_T3_SOUTH_B1_O),
    .ready_in(SB_T3_SOUTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T3_SOUTH_B1_ready_out),
    .valid_in(RMUX_T3_SOUTH_B1_valid_in),
    .valid_out(RMUX_T3_SOUTH_B1_valid_out),
    .S(RMUX_T3_SOUTH_B1_sel_value_O),
    .out_sel(RMUX_T3_SOUTH_B1_out_sel)
);
SliceWrapper_32_10_11 RMUX_T3_SOUTH_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T3_SOUTH_B1_sel_value_O)
);
wire [0:0] RMUX_T3_WEST_B1_I [1:0];
assign RMUX_T3_WEST_B1_I[1] = REG_T3_WEST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T3_WEST_B1_I[0] = MUX_SB_T3_WEST_SB_OUT_B1_O;
wire [1:0] RMUX_T3_WEST_B1_valid_in;
assign RMUX_T3_WEST_B1_valid_in = {REG_T3_WEST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T3_WEST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T3_WEST_B1 (
    .I(RMUX_T3_WEST_B1_I),
    .O(RMUX_T3_WEST_B1_O),
    .ready_in(SB_T3_WEST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T3_WEST_B1_ready_out),
    .valid_in(RMUX_T3_WEST_B1_valid_in),
    .valid_out(RMUX_T3_WEST_B1_valid_out),
    .S(RMUX_T3_WEST_B1_sel_value_O),
    .out_sel(RMUX_T3_WEST_B1_out_sel)
);
SliceWrapper_32_11_12 RMUX_T3_WEST_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T3_WEST_B1_sel_value_O)
);
wire [0:0] RMUX_T4_EAST_B1_I [1:0];
assign RMUX_T4_EAST_B1_I[1] = REG_T4_EAST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T4_EAST_B1_I[0] = MUX_SB_T4_EAST_SB_OUT_B1_O;
wire [1:0] RMUX_T4_EAST_B1_valid_in;
assign RMUX_T4_EAST_B1_valid_in = {REG_T4_EAST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T4_EAST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T4_EAST_B1 (
    .I(RMUX_T4_EAST_B1_I),
    .O(RMUX_T4_EAST_B1_O),
    .ready_in(SB_T4_EAST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T4_EAST_B1_ready_out),
    .valid_in(RMUX_T4_EAST_B1_valid_in),
    .valid_out(RMUX_T4_EAST_B1_valid_out),
    .S(RMUX_T4_EAST_B1_sel_value_O),
    .out_sel(RMUX_T4_EAST_B1_out_sel)
);
SliceWrapper_32_12_13 RMUX_T4_EAST_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T4_EAST_B1_sel_value_O)
);
wire [0:0] RMUX_T4_NORTH_B1_I [1:0];
assign RMUX_T4_NORTH_B1_I[1] = REG_T4_NORTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T4_NORTH_B1_I[0] = MUX_SB_T4_NORTH_SB_OUT_B1_O;
wire [1:0] RMUX_T4_NORTH_B1_valid_in;
assign RMUX_T4_NORTH_B1_valid_in = {REG_T4_NORTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T4_NORTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T4_NORTH_B1 (
    .I(RMUX_T4_NORTH_B1_I),
    .O(RMUX_T4_NORTH_B1_O),
    .ready_in(SB_T4_NORTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T4_NORTH_B1_ready_out),
    .valid_in(RMUX_T4_NORTH_B1_valid_in),
    .valid_out(RMUX_T4_NORTH_B1_valid_out),
    .S(RMUX_T4_NORTH_B1_sel_value_O),
    .out_sel(RMUX_T4_NORTH_B1_out_sel)
);
SliceWrapper_32_13_14 RMUX_T4_NORTH_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T4_NORTH_B1_sel_value_O)
);
wire [0:0] RMUX_T4_SOUTH_B1_I [1:0];
assign RMUX_T4_SOUTH_B1_I[1] = REG_T4_SOUTH_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T4_SOUTH_B1_I[0] = MUX_SB_T4_SOUTH_SB_OUT_B1_O;
wire [1:0] RMUX_T4_SOUTH_B1_valid_in;
assign RMUX_T4_SOUTH_B1_valid_in = {REG_T4_SOUTH_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T4_SOUTH_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T4_SOUTH_B1 (
    .I(RMUX_T4_SOUTH_B1_I),
    .O(RMUX_T4_SOUTH_B1_O),
    .ready_in(SB_T4_SOUTH_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T4_SOUTH_B1_ready_out),
    .valid_in(RMUX_T4_SOUTH_B1_valid_in),
    .valid_out(RMUX_T4_SOUTH_B1_valid_out),
    .S(RMUX_T4_SOUTH_B1_sel_value_O),
    .out_sel(RMUX_T4_SOUTH_B1_out_sel)
);
SliceWrapper_32_14_15 RMUX_T4_SOUTH_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T4_SOUTH_B1_sel_value_O)
);
wire [0:0] RMUX_T4_WEST_B1_I [1:0];
assign RMUX_T4_WEST_B1_I[1] = REG_T4_WEST_B1$SplitFifo_1_inst0_data_out;
assign RMUX_T4_WEST_B1_I[0] = MUX_SB_T4_WEST_SB_OUT_B1_O;
wire [1:0] RMUX_T4_WEST_B1_valid_in;
assign RMUX_T4_WEST_B1_valid_in = {REG_T4_WEST_B1$SplitFifo_1_inst0_valid1[0],MUX_SB_T4_WEST_SB_OUT_B1_valid_out};
mux_aoi_ready_valid_2_1 RMUX_T4_WEST_B1 (
    .I(RMUX_T4_WEST_B1_I),
    .O(RMUX_T4_WEST_B1_O),
    .ready_in(SB_T4_WEST_SB_OUT_B1_ready_in),
    .ready_out(RMUX_T4_WEST_B1_ready_out),
    .valid_in(RMUX_T4_WEST_B1_valid_in),
    .valid_out(RMUX_T4_WEST_B1_valid_out),
    .S(RMUX_T4_WEST_B1_sel_value_O),
    .out_sel(RMUX_T4_WEST_B1_out_sel)
);
SliceWrapper_32_15_16 RMUX_T4_WEST_B1_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T4_WEST_B1_sel_value_O)
);
SliceWrapper_32_16_17 SB_T0_EAST_SB_IN_B1_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_EAST_SB_IN_B1_enable_value_O)
);
FanoutHash_4678C6877F96240E SB_T0_EAST_SB_IN_B1_fan_in (
    .E2(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T0_WEST_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T0_EAST_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T3_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T0_EAST_SB_OUT_B1_FANOUT_I;
assign SB_T0_EAST_SB_OUT_B1_FANOUT_I = {REG_T0_EAST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T0_EAST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T0_EAST_SB_OUT_B1_FANOUT (
    .S(RMUX_T0_EAST_B1_out_sel),
    .O(SB_T0_EAST_SB_OUT_B1_FANOUT_O),
    .I(SB_T0_EAST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_32_17_18 SB_T0_EAST_SB_OUT_B1_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_EAST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_32_18_21 SB_T0_EAST_SB_OUT_B1_sel_value (
    .I(config_reg_2_O),
    .O(SB_T0_EAST_SB_OUT_B1_sel_value_O)
);
SliceWrapper_32_21_22 SB_T0_NORTH_SB_IN_B1_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_NORTH_SB_IN_B1_enable_value_O)
);
FanoutHash_F95D10B01D02012 SB_T0_NORTH_SB_IN_B1_fan_in (
    .E2(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T0_WEST_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T0_NORTH_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T1_EAST_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T0_NORTH_SB_OUT_B1_FANOUT_I;
assign SB_T0_NORTH_SB_OUT_B1_FANOUT_I = {REG_T0_NORTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T0_NORTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T0_NORTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T0_NORTH_B1_out_sel),
    .O(SB_T0_NORTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T0_NORTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_32_22_23 SB_T0_NORTH_SB_OUT_B1_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_NORTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_32_23_26 SB_T0_NORTH_SB_OUT_B1_sel_value (
    .I(config_reg_2_O),
    .O(SB_T0_NORTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_32_26_27 SB_T0_SOUTH_SB_IN_B1_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_SOUTH_SB_IN_B1_enable_value_O)
);
FanoutHash_99D793215CEDDD5 SB_T0_SOUTH_SB_IN_B1_fan_in (
    .E2(SB_T1_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T3_EAST_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T0_SOUTH_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T0_NORTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T0_SOUTH_SB_OUT_B1_FANOUT_I;
assign SB_T0_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T0_SOUTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T0_SOUTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T0_SOUTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T0_SOUTH_B1_out_sel),
    .O(SB_T0_SOUTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T0_SOUTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_32_27_28 SB_T0_SOUTH_SB_OUT_B1_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_SOUTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_32_28_31 SB_T0_SOUTH_SB_OUT_B1_sel_value (
    .I(config_reg_2_O),
    .O(SB_T0_SOUTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_32_31_32 SB_T0_WEST_SB_IN_B1_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_WEST_SB_IN_B1_enable_value_O)
);
FanoutHash_3A0064632A577CF5 SB_T0_WEST_SB_IN_B1_fan_in (
    .E2(SB_T0_EAST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T0_WEST_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T4_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T0_WEST_SB_OUT_B1_FANOUT_I;
assign SB_T0_WEST_SB_OUT_B1_FANOUT_I = {REG_T0_WEST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T0_WEST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T0_WEST_SB_OUT_B1_FANOUT (
    .S(RMUX_T0_WEST_B1_out_sel),
    .O(SB_T0_WEST_SB_OUT_B1_FANOUT_O),
    .I(SB_T0_WEST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_31_0_1 SB_T0_WEST_SB_OUT_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T0_WEST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_31_1_4 SB_T0_WEST_SB_OUT_B1_sel_value (
    .I(config_reg_3_O),
    .O(SB_T0_WEST_SB_OUT_B1_sel_value_O)
);
SliceWrapper_31_4_5 SB_T1_EAST_SB_IN_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_EAST_SB_IN_B1_enable_value_O)
);
FanoutHash_1130FCC7DFE98006 SB_T1_EAST_SB_IN_B1_fan_in (
    .E2(SB_T2_SOUTH_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T0_NORTH_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T1_EAST_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T1_WEST_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T1_EAST_SB_OUT_B1_FANOUT_I;
assign SB_T1_EAST_SB_OUT_B1_FANOUT_I = {REG_T1_EAST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T1_EAST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T1_EAST_SB_OUT_B1_FANOUT (
    .S(RMUX_T1_EAST_B1_out_sel),
    .O(SB_T1_EAST_SB_OUT_B1_FANOUT_O),
    .I(SB_T1_EAST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_31_5_6 SB_T1_EAST_SB_OUT_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_EAST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_31_6_9 SB_T1_EAST_SB_OUT_B1_sel_value (
    .I(config_reg_3_O),
    .O(SB_T1_EAST_SB_OUT_B1_sel_value_O)
);
SliceWrapper_31_9_10 SB_T1_NORTH_SB_IN_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_NORTH_SB_IN_B1_enable_value_O)
);
FanoutHash_31555E0CDC460B97 SB_T1_NORTH_SB_IN_B1_fan_in (
    .E2(SB_T4_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T2_EAST_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T1_NORTH_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T1_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T1_NORTH_SB_OUT_B1_FANOUT_I;
assign SB_T1_NORTH_SB_OUT_B1_FANOUT_I = {REG_T1_NORTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T1_NORTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T1_NORTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T1_NORTH_B1_out_sel),
    .O(SB_T1_NORTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T1_NORTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_31_10_11 SB_T1_NORTH_SB_OUT_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_NORTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_31_11_14 SB_T1_NORTH_SB_OUT_B1_sel_value (
    .I(config_reg_3_O),
    .O(SB_T1_NORTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_31_14_15 SB_T1_SOUTH_SB_IN_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_SOUTH_SB_IN_B1_enable_value_O)
);
FanoutHash_4FF010386DB0B737 SB_T1_SOUTH_SB_IN_B1_fan_in (
    .E2(SB_T2_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T2_EAST_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T1_SOUTH_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T1_NORTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T1_SOUTH_SB_OUT_B1_FANOUT_I;
assign SB_T1_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T1_SOUTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T1_SOUTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T1_SOUTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T1_SOUTH_B1_out_sel),
    .O(SB_T1_SOUTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T1_SOUTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_31_15_16 SB_T1_SOUTH_SB_OUT_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_SOUTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_31_16_19 SB_T1_SOUTH_SB_OUT_B1_sel_value (
    .I(config_reg_3_O),
    .O(SB_T1_SOUTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_31_19_20 SB_T1_WEST_SB_IN_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_WEST_SB_IN_B1_enable_value_O)
);
FanoutHash_1A568579D8E9714B SB_T1_WEST_SB_IN_B1_fan_in (
    .E2(SB_T1_EAST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T1_WEST_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T0_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T1_WEST_SB_OUT_B1_FANOUT_I;
assign SB_T1_WEST_SB_OUT_B1_FANOUT_I = {REG_T1_WEST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T1_WEST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T1_WEST_SB_OUT_B1_FANOUT (
    .S(RMUX_T1_WEST_B1_out_sel),
    .O(SB_T1_WEST_SB_OUT_B1_FANOUT_O),
    .I(SB_T1_WEST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_31_20_21 SB_T1_WEST_SB_OUT_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_WEST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_31_21_24 SB_T1_WEST_SB_OUT_B1_sel_value (
    .I(config_reg_3_O),
    .O(SB_T1_WEST_SB_OUT_B1_sel_value_O)
);
SliceWrapper_31_24_25 SB_T2_EAST_SB_IN_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T2_EAST_SB_IN_B1_enable_value_O)
);
FanoutHash_278348DB702230E6 SB_T2_EAST_SB_IN_B1_fan_in (
    .E2(SB_T2_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T2_EAST_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T1_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T2_EAST_SB_OUT_B1_FANOUT_I;
assign SB_T2_EAST_SB_OUT_B1_FANOUT_I = {REG_T2_EAST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T2_EAST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T2_EAST_SB_OUT_B1_FANOUT (
    .S(RMUX_T2_EAST_B1_out_sel),
    .O(SB_T2_EAST_SB_OUT_B1_FANOUT_O),
    .I(SB_T2_EAST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_31_25_26 SB_T2_EAST_SB_OUT_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T2_EAST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_31_26_29 SB_T2_EAST_SB_OUT_B1_sel_value (
    .I(config_reg_3_O),
    .O(SB_T2_EAST_SB_OUT_B1_sel_value_O)
);
SliceWrapper_31_29_30 SB_T2_NORTH_SB_IN_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T2_NORTH_SB_IN_B1_enable_value_O)
);
FanoutHash_6EB42FA08A9B7B5B SB_T2_NORTH_SB_IN_B1_fan_in (
    .E2(SB_T3_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T3_EAST_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T2_NORTH_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T2_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T2_NORTH_SB_OUT_B1_FANOUT_I;
assign SB_T2_NORTH_SB_OUT_B1_FANOUT_I = {REG_T2_NORTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T2_NORTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T2_NORTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T2_NORTH_B1_out_sel),
    .O(SB_T2_NORTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T2_NORTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_31_30_31 SB_T2_NORTH_SB_OUT_B1_enable_value (
    .I(config_reg_3_O),
    .O(SB_T2_NORTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_30_0_3 SB_T2_NORTH_SB_OUT_B1_sel_value (
    .I(config_reg_4_O),
    .O(SB_T2_NORTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_30_3_4 SB_T2_SOUTH_SB_IN_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T2_SOUTH_SB_IN_B1_enable_value_O)
);
FanoutHash_308BAC760F688049 SB_T2_SOUTH_SB_IN_B1_fan_in (
    .E2(SB_T3_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T1_EAST_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T1_EAST_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T1_EAST_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T2_SOUTH_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T2_NORTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T2_SOUTH_SB_OUT_B1_FANOUT_I;
assign SB_T2_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T2_SOUTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T2_SOUTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T2_SOUTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T2_SOUTH_B1_out_sel),
    .O(SB_T2_SOUTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T2_SOUTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_30_4_5 SB_T2_SOUTH_SB_OUT_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T2_SOUTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_30_5_8 SB_T2_SOUTH_SB_OUT_B1_sel_value (
    .I(config_reg_4_O),
    .O(SB_T2_SOUTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_30_8_9 SB_T2_WEST_SB_IN_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T2_WEST_SB_IN_B1_enable_value_O)
);
FanoutHash_F8E7A0823DC8CDD SB_T2_WEST_SB_IN_B1_fan_in (
    .E2(SB_T2_EAST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T1_SOUTH_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T2_EAST_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T2_EAST_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T1_SOUTH_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T2_WEST_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T1_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T2_WEST_SB_OUT_B1_FANOUT_I;
assign SB_T2_WEST_SB_OUT_B1_FANOUT_I = {REG_T2_WEST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T2_WEST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T2_WEST_SB_OUT_B1_FANOUT (
    .S(RMUX_T2_WEST_B1_out_sel),
    .O(SB_T2_WEST_SB_OUT_B1_FANOUT_O),
    .I(SB_T2_WEST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_30_9_10 SB_T2_WEST_SB_OUT_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T2_WEST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_30_10_13 SB_T2_WEST_SB_OUT_B1_sel_value (
    .I(config_reg_4_O),
    .O(SB_T2_WEST_SB_OUT_B1_sel_value_O)
);
SliceWrapper_30_13_14 SB_T3_EAST_SB_IN_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_EAST_SB_IN_B1_enable_value_O)
);
FanoutHash_D70CFBE8EA3CE7F SB_T3_EAST_SB_IN_B1_fan_in (
    .E2(SB_T3_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T0_SOUTH_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T3_WEST_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T3_WEST_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T0_SOUTH_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T0_SOUTH_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T3_EAST_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T2_NORTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T3_EAST_SB_OUT_B1_FANOUT_I;
assign SB_T3_EAST_SB_OUT_B1_FANOUT_I = {REG_T3_EAST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T3_EAST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T3_EAST_SB_OUT_B1_FANOUT (
    .S(RMUX_T3_EAST_B1_out_sel),
    .O(SB_T3_EAST_SB_OUT_B1_FANOUT_O),
    .I(SB_T3_EAST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_30_14_15 SB_T3_EAST_SB_OUT_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_EAST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_30_15_18 SB_T3_EAST_SB_OUT_B1_sel_value (
    .I(config_reg_4_O),
    .O(SB_T3_EAST_SB_OUT_B1_sel_value_O)
);
SliceWrapper_30_18_19 SB_T3_NORTH_SB_IN_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_NORTH_SB_IN_B1_enable_value_O)
);
FanoutHash_5DE101F5B6936D07 SB_T3_NORTH_SB_IN_B1_fan_in (
    .E2(SB_T3_SOUTH_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T2_WEST_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T2_WEST_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T2_WEST_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T3_NORTH_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T4_EAST_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T3_NORTH_SB_OUT_B1_FANOUT_I;
assign SB_T3_NORTH_SB_OUT_B1_FANOUT_I = {REG_T3_NORTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T3_NORTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T3_NORTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T3_NORTH_B1_out_sel),
    .O(SB_T3_NORTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T3_NORTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_30_19_20 SB_T3_NORTH_SB_OUT_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_NORTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_30_20_23 SB_T3_NORTH_SB_OUT_B1_sel_value (
    .I(config_reg_4_O),
    .O(SB_T3_NORTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_30_23_24 SB_T3_SOUTH_SB_IN_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_SOUTH_SB_IN_B1_enable_value_O)
);
FanoutHash_13B77C2790BDE4E2 SB_T3_SOUTH_SB_IN_B1_fan_in (
    .E2(SB_T4_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T0_EAST_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T3_SOUTH_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T3_NORTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T3_SOUTH_SB_OUT_B1_FANOUT_I;
assign SB_T3_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T3_SOUTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T3_SOUTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T3_SOUTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T3_SOUTH_B1_out_sel),
    .O(SB_T3_SOUTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T3_SOUTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_30_24_25 SB_T3_SOUTH_SB_OUT_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_SOUTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_30_25_28 SB_T3_SOUTH_SB_OUT_B1_sel_value (
    .I(config_reg_4_O),
    .O(SB_T3_SOUTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_30_28_29 SB_T3_WEST_SB_IN_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_WEST_SB_IN_B1_enable_value_O)
);
FanoutHash_7FDF2D3240D4A947 SB_T3_WEST_SB_IN_B1_fan_in (
    .E2(SB_T3_EAST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T2_SOUTH_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T2_NORTH_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T3_EAST_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T3_EAST_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T2_NORTH_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T2_NORTH_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T2_SOUTH_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T3_WEST_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T2_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T3_WEST_SB_OUT_B1_FANOUT_I;
assign SB_T3_WEST_SB_OUT_B1_FANOUT_I = {REG_T3_WEST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T3_WEST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T3_WEST_SB_OUT_B1_FANOUT (
    .S(RMUX_T3_WEST_B1_out_sel),
    .O(SB_T3_WEST_SB_OUT_B1_FANOUT_O),
    .I(SB_T3_WEST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_30_29_30 SB_T3_WEST_SB_OUT_B1_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_WEST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_23_0_3 SB_T3_WEST_SB_OUT_B1_sel_value (
    .I(config_reg_5_O),
    .O(SB_T3_WEST_SB_OUT_B1_sel_value_O)
);
SliceWrapper_23_3_4 SB_T4_EAST_SB_IN_B1_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_EAST_SB_IN_B1_enable_value_O)
);
FanoutHash_11B554A18790BBBC SB_T4_EAST_SB_IN_B1_fan_in (
    .E2(SB_T4_WEST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T3_NORTH_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T4_WEST_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T4_WEST_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T3_NORTH_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T3_NORTH_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T4_EAST_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T4_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T4_EAST_SB_OUT_B1_FANOUT_I;
assign SB_T4_EAST_SB_OUT_B1_FANOUT_I = {REG_T4_EAST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T4_EAST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T4_EAST_SB_OUT_B1_FANOUT (
    .S(RMUX_T4_EAST_B1_out_sel),
    .O(SB_T4_EAST_SB_OUT_B1_FANOUT_O),
    .I(SB_T4_EAST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_23_4_5 SB_T4_EAST_SB_OUT_B1_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_EAST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_23_5_8 SB_T4_EAST_SB_OUT_B1_sel_value (
    .I(config_reg_5_O),
    .O(SB_T4_EAST_SB_OUT_B1_sel_value_O)
);
SliceWrapper_23_8_9 SB_T4_NORTH_SB_IN_B1_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_NORTH_SB_IN_B1_enable_value_O)
);
FanoutHash_37B926A0CDF82FCC SB_T4_NORTH_SB_IN_B1_fan_in (
    .E2(SB_T4_SOUTH_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T0_EAST_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T1_WEST_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T4_SOUTH_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T4_SOUTH_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T1_WEST_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T1_WEST_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T0_EAST_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T4_NORTH_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T0_EAST_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T4_NORTH_SB_OUT_B1_FANOUT_I;
assign SB_T4_NORTH_SB_OUT_B1_FANOUT_I = {REG_T4_NORTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T4_NORTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T4_NORTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T4_NORTH_B1_out_sel),
    .O(SB_T4_NORTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T4_NORTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_23_9_10 SB_T4_NORTH_SB_OUT_B1_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_NORTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_23_10_13 SB_T4_NORTH_SB_OUT_B1_sel_value (
    .I(config_reg_5_O),
    .O(SB_T4_NORTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_23_13_14 SB_T4_SOUTH_SB_IN_B1_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_SOUTH_SB_IN_B1_enable_value_O)
);
FanoutHash_1B10C32F008C11AC SB_T4_SOUTH_SB_IN_B1_fan_in (
    .E2(SB_T4_NORTH_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T0_WEST_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T4_NORTH_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T4_NORTH_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T0_WEST_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T0_WEST_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T4_SOUTH_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T4_EAST_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T4_SOUTH_SB_OUT_B1_FANOUT_I;
assign SB_T4_SOUTH_SB_OUT_B1_FANOUT_I = {REG_T4_SOUTH_B1$SplitFifo_1_inst0_ready0[0],RMUX_T4_SOUTH_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T4_SOUTH_SB_OUT_B1_FANOUT (
    .S(RMUX_T4_SOUTH_B1_out_sel),
    .O(SB_T4_SOUTH_SB_OUT_B1_FANOUT_O),
    .I(SB_T4_SOUTH_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_23_14_15 SB_T4_SOUTH_SB_OUT_B1_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_SOUTH_SB_OUT_B1_enable_value_O)
);
SliceWrapper_23_15_18 SB_T4_SOUTH_SB_OUT_B1_sel_value (
    .I(config_reg_5_O),
    .O(SB_T4_SOUTH_SB_OUT_B1_sel_value_O)
);
SliceWrapper_23_18_19 SB_T4_WEST_SB_IN_B1_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_WEST_SB_IN_B1_enable_value_O)
);
FanoutHash_660E59B0DDACF452 SB_T4_WEST_SB_IN_B1_fan_in (
    .E2(SB_T4_EAST_SB_OUT_B1_enable_value_O),
    .S1(MUX_SB_T3_SOUTH_SB_OUT_B1_out_sel),
    .I3(MEM_input_width_1_num_0_ready),
    .S0(MUX_SB_T1_NORTH_SB_OUT_B1_out_sel),
    .E5(const_0_1_out),
    .I2(MUX_SB_T4_EAST_SB_OUT_B1_ready_out),
    .S3(MEM_input_width_1_num_0_out_sel),
    .S2(MUX_SB_T4_EAST_SB_OUT_B1_out_sel),
    .E3(MEM_input_width_1_num_0_enable),
    .E0(SB_T1_NORTH_SB_OUT_B1_enable_value_O),
    .S4(MEM_input_width_1_num_1_out_sel),
    .I0(MUX_SB_T1_NORTH_SB_OUT_B1_ready_out),
    .E4(MEM_input_width_1_num_1_enable),
    .S5(const_0_32_out),
    .I1(MUX_SB_T3_SOUTH_SB_OUT_B1_ready_out),
    .I5(const_0_1_out),
    .O(SB_T4_WEST_SB_IN_B1_fan_in_O),
    .I4(MEM_input_width_1_num_1_ready),
    .E1(SB_T3_SOUTH_SB_OUT_B1_enable_value_O)
);
wire [1:0] SB_T4_WEST_SB_OUT_B1_FANOUT_I;
assign SB_T4_WEST_SB_OUT_B1_FANOUT_I = {REG_T4_WEST_B1$SplitFifo_1_inst0_ready0[0],RMUX_T4_WEST_B1_ready_out};
ExclusiveNodeFanout_H2 SB_T4_WEST_SB_OUT_B1_FANOUT (
    .S(RMUX_T4_WEST_B1_out_sel),
    .O(SB_T4_WEST_SB_OUT_B1_FANOUT_O),
    .I(SB_T4_WEST_SB_OUT_B1_FANOUT_I)
);
SliceWrapper_23_19_20 SB_T4_WEST_SB_OUT_B1_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_WEST_SB_OUT_B1_enable_value_O)
);
SliceWrapper_23_20_23 SB_T4_WEST_SB_OUT_B1_sel_value (
    .I(config_reg_5_O),
    .O(SB_T4_WEST_SB_OUT_B1_sel_value_O)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T0_EAST_SB_IN_B1 (
    .I(SB_T0_EAST_SB_IN_B1),
    .O(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .ready_in(SB_T0_EAST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T0_EAST_SB_IN_B1_ready_out),
    .valid_in(SB_T0_EAST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T0_EAST_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T0_NORTH_SB_IN_B1 (
    .I(SB_T0_NORTH_SB_IN_B1),
    .O(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .ready_in(SB_T0_NORTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T0_NORTH_SB_IN_B1_ready_out),
    .valid_in(SB_T0_NORTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T0_NORTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T0_SOUTH_SB_IN_B1 (
    .I(SB_T0_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .ready_in(SB_T0_SOUTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T0_SOUTH_SB_IN_B1_ready_out),
    .valid_in(SB_T0_SOUTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T0_SOUTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T0_WEST_SB_IN_B1 (
    .I(SB_T0_WEST_SB_IN_B1),
    .O(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .ready_in(SB_T0_WEST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T0_WEST_SB_IN_B1_ready_out),
    .valid_in(SB_T0_WEST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T0_WEST_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T1_EAST_SB_IN_B1 (
    .I(SB_T1_EAST_SB_IN_B1),
    .O(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .ready_in(SB_T1_EAST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T1_EAST_SB_IN_B1_ready_out),
    .valid_in(SB_T1_EAST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T1_EAST_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T1_NORTH_SB_IN_B1 (
    .I(SB_T1_NORTH_SB_IN_B1),
    .O(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .ready_in(SB_T1_NORTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T1_NORTH_SB_IN_B1_ready_out),
    .valid_in(SB_T1_NORTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T1_NORTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T1_SOUTH_SB_IN_B1 (
    .I(SB_T1_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .ready_in(SB_T1_SOUTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T1_SOUTH_SB_IN_B1_ready_out),
    .valid_in(SB_T1_SOUTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T1_SOUTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T1_WEST_SB_IN_B1 (
    .I(SB_T1_WEST_SB_IN_B1),
    .O(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .ready_in(SB_T1_WEST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T1_WEST_SB_IN_B1_ready_out),
    .valid_in(SB_T1_WEST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T1_WEST_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T2_EAST_SB_IN_B1 (
    .I(SB_T2_EAST_SB_IN_B1),
    .O(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .ready_in(SB_T2_EAST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T2_EAST_SB_IN_B1_ready_out),
    .valid_in(SB_T2_EAST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T2_EAST_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T2_NORTH_SB_IN_B1 (
    .I(SB_T2_NORTH_SB_IN_B1),
    .O(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .ready_in(SB_T2_NORTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T2_NORTH_SB_IN_B1_ready_out),
    .valid_in(SB_T2_NORTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T2_NORTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T2_SOUTH_SB_IN_B1 (
    .I(SB_T2_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .ready_in(SB_T2_SOUTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T2_SOUTH_SB_IN_B1_ready_out),
    .valid_in(SB_T2_SOUTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T2_SOUTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T2_WEST_SB_IN_B1 (
    .I(SB_T2_WEST_SB_IN_B1),
    .O(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .ready_in(SB_T2_WEST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T2_WEST_SB_IN_B1_ready_out),
    .valid_in(SB_T2_WEST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T2_WEST_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T3_EAST_SB_IN_B1 (
    .I(SB_T3_EAST_SB_IN_B1),
    .O(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .ready_in(SB_T3_EAST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T3_EAST_SB_IN_B1_ready_out),
    .valid_in(SB_T3_EAST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T3_EAST_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T3_NORTH_SB_IN_B1 (
    .I(SB_T3_NORTH_SB_IN_B1),
    .O(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .ready_in(SB_T3_NORTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T3_NORTH_SB_IN_B1_ready_out),
    .valid_in(SB_T3_NORTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T3_NORTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T3_SOUTH_SB_IN_B1 (
    .I(SB_T3_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .ready_in(SB_T3_SOUTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T3_SOUTH_SB_IN_B1_ready_out),
    .valid_in(SB_T3_SOUTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T3_SOUTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T3_WEST_SB_IN_B1 (
    .I(SB_T3_WEST_SB_IN_B1),
    .O(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .ready_in(SB_T3_WEST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T3_WEST_SB_IN_B1_ready_out),
    .valid_in(SB_T3_WEST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T3_WEST_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T4_EAST_SB_IN_B1 (
    .I(SB_T4_EAST_SB_IN_B1),
    .O(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .ready_in(SB_T4_EAST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T4_EAST_SB_IN_B1_ready_out),
    .valid_in(SB_T4_EAST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T4_EAST_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T4_NORTH_SB_IN_B1 (
    .I(SB_T4_NORTH_SB_IN_B1),
    .O(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .ready_in(SB_T4_NORTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T4_NORTH_SB_IN_B1_ready_out),
    .valid_in(SB_T4_NORTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T4_NORTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T4_SOUTH_SB_IN_B1 (
    .I(SB_T4_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .ready_in(SB_T4_SOUTH_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T4_SOUTH_SB_IN_B1_ready_out),
    .valid_in(SB_T4_SOUTH_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T4_SOUTH_SB_IN_B1_valid_out)
);
MuxWrapperAOI_1_1_RegularReadyValid WIRE_SB_T4_WEST_SB_IN_B1 (
    .I(SB_T4_WEST_SB_IN_B1),
    .O(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .ready_in(SB_T4_WEST_SB_IN_B1_fan_in_O[0]),
    .ready_out(WIRE_SB_T4_WEST_SB_IN_B1_ready_out),
    .valid_in(SB_T4_WEST_SB_IN_B1_valid_in),
    .valid_out(WIRE_SB_T4_WEST_SB_IN_B1_valid_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_23_32_inst0$bit_const_0_None (
    .out(ZextWrapper_23_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_23_32_inst0$self_O_out;
assign ZextWrapper_23_32_inst0$self_O_out = {ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,config_reg_5_O};
mantle_wire__typeBitIn32 ZextWrapper_23_32_inst0$self_O (
    .in(ZextWrapper_23_32_inst0$self_O_in),
    .out(ZextWrapper_23_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_30_32_inst0$bit_const_0_None (
    .out(ZextWrapper_30_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_30_32_inst0$self_O_out;
assign ZextWrapper_30_32_inst0$self_O_out = {ZextWrapper_30_32_inst0$bit_const_0_None_out,ZextWrapper_30_32_inst0$bit_const_0_None_out,config_reg_4_O};
mantle_wire__typeBitIn32 ZextWrapper_30_32_inst0$self_O (
    .in(ZextWrapper_30_32_inst0$self_O_in),
    .out(ZextWrapper_30_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_31_32_inst0$bit_const_0_None (
    .out(ZextWrapper_31_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_31_32_inst0$self_O_out;
assign ZextWrapper_31_32_inst0$self_O_out = {ZextWrapper_31_32_inst0$bit_const_0_None_out,config_reg_3_O};
mantle_wire__typeBitIn32 ZextWrapper_31_32_inst0$self_O (
    .in(ZextWrapper_31_32_inst0$self_O_in),
    .out(ZextWrapper_31_32_inst0$self_O_out)
);
coreir_and #(
    .width(1)
) and1_inst0 (
    .in0(coreir_eq_1_inst0_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst0_out)
);
coreir_and #(
    .width(1)
) and1_inst1 (
    .in0(coreir_eq_1_inst1_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst1_out)
);
coreir_and #(
    .width(1)
) and1_inst10 (
    .in0(coreir_eq_1_inst10_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst10_out)
);
coreir_and #(
    .width(1)
) and1_inst11 (
    .in0(coreir_eq_1_inst11_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst11_out)
);
coreir_and #(
    .width(1)
) and1_inst12 (
    .in0(coreir_eq_1_inst12_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst12_out)
);
coreir_and #(
    .width(1)
) and1_inst13 (
    .in0(coreir_eq_1_inst13_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst13_out)
);
coreir_and #(
    .width(1)
) and1_inst14 (
    .in0(coreir_eq_1_inst14_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst14_out)
);
coreir_and #(
    .width(1)
) and1_inst15 (
    .in0(coreir_eq_1_inst15_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst15_out)
);
coreir_and #(
    .width(1)
) and1_inst16 (
    .in0(coreir_eq_1_inst16_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst16_out)
);
coreir_and #(
    .width(1)
) and1_inst17 (
    .in0(coreir_eq_1_inst17_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst17_out)
);
coreir_and #(
    .width(1)
) and1_inst18 (
    .in0(coreir_eq_1_inst18_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst18_out)
);
coreir_and #(
    .width(1)
) and1_inst19 (
    .in0(coreir_eq_1_inst19_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst19_out)
);
coreir_and #(
    .width(1)
) and1_inst2 (
    .in0(coreir_eq_1_inst2_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst2_out)
);
coreir_and #(
    .width(1)
) and1_inst3 (
    .in0(coreir_eq_1_inst3_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst3_out)
);
coreir_and #(
    .width(1)
) and1_inst4 (
    .in0(coreir_eq_1_inst4_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst4_out)
);
coreir_and #(
    .width(1)
) and1_inst5 (
    .in0(coreir_eq_1_inst5_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst5_out)
);
coreir_and #(
    .width(1)
) and1_inst6 (
    .in0(coreir_eq_1_inst6_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst6_out)
);
coreir_and #(
    .width(1)
) and1_inst7 (
    .in0(coreir_eq_1_inst7_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst7_out)
);
coreir_and #(
    .width(1)
) and1_inst8 (
    .in0(coreir_eq_1_inst8_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst8_out)
);
coreir_and #(
    .width(1)
) and1_inst9 (
    .in0(coreir_eq_1_inst9_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst9_out)
);
wire [7:0] config_reg_0_config_addr;
assign config_reg_0_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_32_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_reg_0_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_1_config_addr;
assign config_reg_1_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_32_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_reg_1_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_2_config_addr;
assign config_reg_2_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_32_8_32_2 config_reg_2 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_2_O),
    .config_addr(config_reg_2_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_3_config_addr;
assign config_reg_3_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_31_8_32_3 config_reg_3 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_3_O),
    .config_addr(config_reg_3_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_4_config_addr;
assign config_reg_4_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_30_8_32_4 config_reg_4 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_4_O),
    .config_addr(config_reg_4_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_5_config_addr;
assign config_reg_5_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_23_8_32_5 config_reg_5 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_5_O),
    .config_addr(config_reg_5_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_const #(
    .value(1'h0),
    .width(1)
) const_0_1 (
    .out(const_0_1_out)
);
coreir_const #(
    .value(32'h00000000),
    .width(32)
) const_0_32 (
    .out(const_0_32_out)
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst0 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_NORTH_B1_sel_value_O),
    .out(coreir_eq_1_inst0_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst1 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_SOUTH_B1_sel_value_O),
    .out(coreir_eq_1_inst1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst10 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_EAST_B1_sel_value_O),
    .out(coreir_eq_1_inst10_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst11 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_WEST_B1_sel_value_O),
    .out(coreir_eq_1_inst11_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst12 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_NORTH_B1_sel_value_O),
    .out(coreir_eq_1_inst12_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst13 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_SOUTH_B1_sel_value_O),
    .out(coreir_eq_1_inst13_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst14 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_EAST_B1_sel_value_O),
    .out(coreir_eq_1_inst14_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst15 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_WEST_B1_sel_value_O),
    .out(coreir_eq_1_inst15_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst16 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_NORTH_B1_sel_value_O),
    .out(coreir_eq_1_inst16_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst17 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_SOUTH_B1_sel_value_O),
    .out(coreir_eq_1_inst17_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst18 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_EAST_B1_sel_value_O),
    .out(coreir_eq_1_inst18_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst19 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_WEST_B1_sel_value_O),
    .out(coreir_eq_1_inst19_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst2 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_EAST_B1_sel_value_O),
    .out(coreir_eq_1_inst2_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst3 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_WEST_B1_sel_value_O),
    .out(coreir_eq_1_inst3_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst4 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_NORTH_B1_sel_value_O),
    .out(coreir_eq_1_inst4_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst5 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_SOUTH_B1_sel_value_O),
    .out(coreir_eq_1_inst5_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst6 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_EAST_B1_sel_value_O),
    .out(coreir_eq_1_inst6_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst7 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_WEST_B1_sel_value_O),
    .out(coreir_eq_1_inst7_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst8 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_NORTH_B1_sel_value_O),
    .out(coreir_eq_1_inst8_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst9 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_SOUTH_B1_sel_value_O),
    .out(coreir_eq_1_inst9_out)
);
wire [31:0] mux_aoi_6_32_inst0_I [5:0];
assign mux_aoi_6_32_inst0_I[5] = ZextWrapper_23_32_inst0$self_O_in;
assign mux_aoi_6_32_inst0_I[4] = ZextWrapper_30_32_inst0$self_O_in;
assign mux_aoi_6_32_inst0_I[3] = ZextWrapper_31_32_inst0$self_O_in;
assign mux_aoi_6_32_inst0_I[2] = config_reg_2_O;
assign mux_aoi_6_32_inst0_I[1] = config_reg_1_O;
assign mux_aoi_6_32_inst0_I[0] = config_reg_0_O;
mux_aoi_6_32 mux_aoi_6_32_inst0 (
    .I(mux_aoi_6_32_inst0_I),
    .O(mux_aoi_6_32_inst0_O),
    .S(self_config_config_addr_out[2:0]),
    .out_sel(mux_aoi_6_32_inst0_out_sel)
);
mantle_wire__typeBit8 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
assign MEM_output_width_1_num_0_ready_out = CB_MEM_output_width_1_num_0_fan_in_O[0];
assign MEM_output_width_1_num_1_ready_out = CB_MEM_output_width_1_num_1_fan_in_O[0];
assign MEM_output_width_1_num_2_ready_out = CB_MEM_output_width_1_num_2_fan_in_O[0];
assign SB_T0_EAST_SB_IN_B1_enable = SB_T0_EAST_SB_IN_B1_enable_value_O[0];
assign SB_T0_EAST_SB_IN_B1_ready_out = WIRE_SB_T0_EAST_SB_IN_B1_ready_out;
assign SB_T0_EAST_SB_OUT_B1 = RMUX_T0_EAST_B1_O;
assign SB_T0_EAST_SB_OUT_B1_enable = SB_T0_EAST_SB_OUT_B1_enable_value_O[0];
assign SB_T0_EAST_SB_OUT_B1_valid_out = RMUX_T0_EAST_B1_valid_out;
assign SB_T0_NORTH_SB_IN_B1_enable = SB_T0_NORTH_SB_IN_B1_enable_value_O[0];
assign SB_T0_NORTH_SB_IN_B1_ready_out = WIRE_SB_T0_NORTH_SB_IN_B1_ready_out;
assign SB_T0_NORTH_SB_OUT_B1 = RMUX_T0_NORTH_B1_O;
assign SB_T0_NORTH_SB_OUT_B1_enable = SB_T0_NORTH_SB_OUT_B1_enable_value_O[0];
assign SB_T0_NORTH_SB_OUT_B1_valid_out = RMUX_T0_NORTH_B1_valid_out;
assign SB_T0_SOUTH_SB_IN_B1_enable = SB_T0_SOUTH_SB_IN_B1_enable_value_O[0];
assign SB_T0_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T0_SOUTH_SB_IN_B1_ready_out;
assign SB_T0_SOUTH_SB_OUT_B1 = RMUX_T0_SOUTH_B1_O;
assign SB_T0_SOUTH_SB_OUT_B1_enable = SB_T0_SOUTH_SB_OUT_B1_enable_value_O[0];
assign SB_T0_SOUTH_SB_OUT_B1_valid_out = RMUX_T0_SOUTH_B1_valid_out;
assign SB_T0_WEST_SB_IN_B1_enable = SB_T0_WEST_SB_IN_B1_enable_value_O[0];
assign SB_T0_WEST_SB_IN_B1_ready_out = WIRE_SB_T0_WEST_SB_IN_B1_ready_out;
assign SB_T0_WEST_SB_OUT_B1 = RMUX_T0_WEST_B1_O;
assign SB_T0_WEST_SB_OUT_B1_enable = SB_T0_WEST_SB_OUT_B1_enable_value_O[0];
assign SB_T0_WEST_SB_OUT_B1_valid_out = RMUX_T0_WEST_B1_valid_out;
assign SB_T1_EAST_SB_IN_B1_enable = SB_T1_EAST_SB_IN_B1_enable_value_O[0];
assign SB_T1_EAST_SB_IN_B1_ready_out = WIRE_SB_T1_EAST_SB_IN_B1_ready_out;
assign SB_T1_EAST_SB_OUT_B1 = RMUX_T1_EAST_B1_O;
assign SB_T1_EAST_SB_OUT_B1_enable = SB_T1_EAST_SB_OUT_B1_enable_value_O[0];
assign SB_T1_EAST_SB_OUT_B1_valid_out = RMUX_T1_EAST_B1_valid_out;
assign SB_T1_NORTH_SB_IN_B1_enable = SB_T1_NORTH_SB_IN_B1_enable_value_O[0];
assign SB_T1_NORTH_SB_IN_B1_ready_out = WIRE_SB_T1_NORTH_SB_IN_B1_ready_out;
assign SB_T1_NORTH_SB_OUT_B1 = RMUX_T1_NORTH_B1_O;
assign SB_T1_NORTH_SB_OUT_B1_enable = SB_T1_NORTH_SB_OUT_B1_enable_value_O[0];
assign SB_T1_NORTH_SB_OUT_B1_valid_out = RMUX_T1_NORTH_B1_valid_out;
assign SB_T1_SOUTH_SB_IN_B1_enable = SB_T1_SOUTH_SB_IN_B1_enable_value_O[0];
assign SB_T1_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T1_SOUTH_SB_IN_B1_ready_out;
assign SB_T1_SOUTH_SB_OUT_B1 = RMUX_T1_SOUTH_B1_O;
assign SB_T1_SOUTH_SB_OUT_B1_enable = SB_T1_SOUTH_SB_OUT_B1_enable_value_O[0];
assign SB_T1_SOUTH_SB_OUT_B1_valid_out = RMUX_T1_SOUTH_B1_valid_out;
assign SB_T1_WEST_SB_IN_B1_enable = SB_T1_WEST_SB_IN_B1_enable_value_O[0];
assign SB_T1_WEST_SB_IN_B1_ready_out = WIRE_SB_T1_WEST_SB_IN_B1_ready_out;
assign SB_T1_WEST_SB_OUT_B1 = RMUX_T1_WEST_B1_O;
assign SB_T1_WEST_SB_OUT_B1_enable = SB_T1_WEST_SB_OUT_B1_enable_value_O[0];
assign SB_T1_WEST_SB_OUT_B1_valid_out = RMUX_T1_WEST_B1_valid_out;
assign SB_T2_EAST_SB_IN_B1_enable = SB_T2_EAST_SB_IN_B1_enable_value_O[0];
assign SB_T2_EAST_SB_IN_B1_ready_out = WIRE_SB_T2_EAST_SB_IN_B1_ready_out;
assign SB_T2_EAST_SB_OUT_B1 = RMUX_T2_EAST_B1_O;
assign SB_T2_EAST_SB_OUT_B1_enable = SB_T2_EAST_SB_OUT_B1_enable_value_O[0];
assign SB_T2_EAST_SB_OUT_B1_valid_out = RMUX_T2_EAST_B1_valid_out;
assign SB_T2_NORTH_SB_IN_B1_enable = SB_T2_NORTH_SB_IN_B1_enable_value_O[0];
assign SB_T2_NORTH_SB_IN_B1_ready_out = WIRE_SB_T2_NORTH_SB_IN_B1_ready_out;
assign SB_T2_NORTH_SB_OUT_B1 = RMUX_T2_NORTH_B1_O;
assign SB_T2_NORTH_SB_OUT_B1_enable = SB_T2_NORTH_SB_OUT_B1_enable_value_O[0];
assign SB_T2_NORTH_SB_OUT_B1_valid_out = RMUX_T2_NORTH_B1_valid_out;
assign SB_T2_SOUTH_SB_IN_B1_enable = SB_T2_SOUTH_SB_IN_B1_enable_value_O[0];
assign SB_T2_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T2_SOUTH_SB_IN_B1_ready_out;
assign SB_T2_SOUTH_SB_OUT_B1 = RMUX_T2_SOUTH_B1_O;
assign SB_T2_SOUTH_SB_OUT_B1_enable = SB_T2_SOUTH_SB_OUT_B1_enable_value_O[0];
assign SB_T2_SOUTH_SB_OUT_B1_valid_out = RMUX_T2_SOUTH_B1_valid_out;
assign SB_T2_WEST_SB_IN_B1_enable = SB_T2_WEST_SB_IN_B1_enable_value_O[0];
assign SB_T2_WEST_SB_IN_B1_ready_out = WIRE_SB_T2_WEST_SB_IN_B1_ready_out;
assign SB_T2_WEST_SB_OUT_B1 = RMUX_T2_WEST_B1_O;
assign SB_T2_WEST_SB_OUT_B1_enable = SB_T2_WEST_SB_OUT_B1_enable_value_O[0];
assign SB_T2_WEST_SB_OUT_B1_valid_out = RMUX_T2_WEST_B1_valid_out;
assign SB_T3_EAST_SB_IN_B1_enable = SB_T3_EAST_SB_IN_B1_enable_value_O[0];
assign SB_T3_EAST_SB_IN_B1_ready_out = WIRE_SB_T3_EAST_SB_IN_B1_ready_out;
assign SB_T3_EAST_SB_OUT_B1 = RMUX_T3_EAST_B1_O;
assign SB_T3_EAST_SB_OUT_B1_enable = SB_T3_EAST_SB_OUT_B1_enable_value_O[0];
assign SB_T3_EAST_SB_OUT_B1_valid_out = RMUX_T3_EAST_B1_valid_out;
assign SB_T3_NORTH_SB_IN_B1_enable = SB_T3_NORTH_SB_IN_B1_enable_value_O[0];
assign SB_T3_NORTH_SB_IN_B1_ready_out = WIRE_SB_T3_NORTH_SB_IN_B1_ready_out;
assign SB_T3_NORTH_SB_OUT_B1 = RMUX_T3_NORTH_B1_O;
assign SB_T3_NORTH_SB_OUT_B1_enable = SB_T3_NORTH_SB_OUT_B1_enable_value_O[0];
assign SB_T3_NORTH_SB_OUT_B1_valid_out = RMUX_T3_NORTH_B1_valid_out;
assign SB_T3_SOUTH_SB_IN_B1_enable = SB_T3_SOUTH_SB_IN_B1_enable_value_O[0];
assign SB_T3_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T3_SOUTH_SB_IN_B1_ready_out;
assign SB_T3_SOUTH_SB_OUT_B1 = RMUX_T3_SOUTH_B1_O;
assign SB_T3_SOUTH_SB_OUT_B1_enable = SB_T3_SOUTH_SB_OUT_B1_enable_value_O[0];
assign SB_T3_SOUTH_SB_OUT_B1_valid_out = RMUX_T3_SOUTH_B1_valid_out;
assign SB_T3_WEST_SB_IN_B1_enable = SB_T3_WEST_SB_IN_B1_enable_value_O[0];
assign SB_T3_WEST_SB_IN_B1_ready_out = WIRE_SB_T3_WEST_SB_IN_B1_ready_out;
assign SB_T3_WEST_SB_OUT_B1 = RMUX_T3_WEST_B1_O;
assign SB_T3_WEST_SB_OUT_B1_enable = SB_T3_WEST_SB_OUT_B1_enable_value_O[0];
assign SB_T3_WEST_SB_OUT_B1_valid_out = RMUX_T3_WEST_B1_valid_out;
assign SB_T4_EAST_SB_IN_B1_enable = SB_T4_EAST_SB_IN_B1_enable_value_O[0];
assign SB_T4_EAST_SB_IN_B1_ready_out = WIRE_SB_T4_EAST_SB_IN_B1_ready_out;
assign SB_T4_EAST_SB_OUT_B1 = RMUX_T4_EAST_B1_O;
assign SB_T4_EAST_SB_OUT_B1_enable = SB_T4_EAST_SB_OUT_B1_enable_value_O[0];
assign SB_T4_EAST_SB_OUT_B1_valid_out = RMUX_T4_EAST_B1_valid_out;
assign SB_T4_NORTH_SB_IN_B1_enable = SB_T4_NORTH_SB_IN_B1_enable_value_O[0];
assign SB_T4_NORTH_SB_IN_B1_ready_out = WIRE_SB_T4_NORTH_SB_IN_B1_ready_out;
assign SB_T4_NORTH_SB_OUT_B1 = RMUX_T4_NORTH_B1_O;
assign SB_T4_NORTH_SB_OUT_B1_enable = SB_T4_NORTH_SB_OUT_B1_enable_value_O[0];
assign SB_T4_NORTH_SB_OUT_B1_valid_out = RMUX_T4_NORTH_B1_valid_out;
assign SB_T4_SOUTH_SB_IN_B1_enable = SB_T4_SOUTH_SB_IN_B1_enable_value_O[0];
assign SB_T4_SOUTH_SB_IN_B1_ready_out = WIRE_SB_T4_SOUTH_SB_IN_B1_ready_out;
assign SB_T4_SOUTH_SB_OUT_B1 = RMUX_T4_SOUTH_B1_O;
assign SB_T4_SOUTH_SB_OUT_B1_enable = SB_T4_SOUTH_SB_OUT_B1_enable_value_O[0];
assign SB_T4_SOUTH_SB_OUT_B1_valid_out = RMUX_T4_SOUTH_B1_valid_out;
assign SB_T4_WEST_SB_IN_B1_enable = SB_T4_WEST_SB_IN_B1_enable_value_O[0];
assign SB_T4_WEST_SB_IN_B1_ready_out = WIRE_SB_T4_WEST_SB_IN_B1_ready_out;
assign SB_T4_WEST_SB_OUT_B1 = RMUX_T4_WEST_B1_O;
assign SB_T4_WEST_SB_OUT_B1_enable = SB_T4_WEST_SB_OUT_B1_enable_value_O[0];
assign SB_T4_WEST_SB_OUT_B1_valid_out = RMUX_T4_WEST_B1_valid_out;
assign read_config_data = mux_aoi_6_32_inst0_O;
endmodule

module SB_ID0_5TRACKS_B17_PE (
    input [0:0] PE_input_width_17_num_0_enable,
    input [31:0] PE_input_width_17_num_0_out_sel,
    input PE_input_width_17_num_0_ready,
    input [0:0] PE_input_width_17_num_1_enable,
    input [31:0] PE_input_width_17_num_1_out_sel,
    input PE_input_width_17_num_1_ready,
    input [0:0] PE_input_width_17_num_2_enable,
    input [31:0] PE_input_width_17_num_2_out_sel,
    input PE_input_width_17_num_2_ready,
    input [0:0] PE_input_width_17_num_3_enable,
    input [31:0] PE_input_width_17_num_3_out_sel,
    input PE_input_width_17_num_3_ready,
    input [16:0] PE_output_width_17_num_0,
    output PE_output_width_17_num_0_ready_out,
    input PE_output_width_17_num_0_valid,
    input [16:0] PE_output_width_17_num_1,
    output PE_output_width_17_num_1_ready_out,
    input PE_output_width_17_num_1_valid,
    input [16:0] PE_output_width_17_num_2,
    output PE_output_width_17_num_2_ready_out,
    input PE_output_width_17_num_2_valid,
    input [0:0] PondTop_input_width_17_num_0_enable,
    input [31:0] PondTop_input_width_17_num_0_out_sel,
    input PondTop_input_width_17_num_0_ready,
    input [0:0] PondTop_input_width_17_num_1_enable,
    input [31:0] PondTop_input_width_17_num_1_out_sel,
    input PondTop_input_width_17_num_1_ready,
    output PondTop_output_width_17_num_0_ready_out,
    input PondTop_output_width_17_num_0_valid,
    input [16:0] PondTop_output_width_17_num_1,
    output PondTop_output_width_17_num_1_ready_out,
    input PondTop_output_width_17_num_1_valid,
    input [16:0] SB_T0_EAST_SB_IN_B17,
    output SB_T0_EAST_SB_IN_B17_enable,
    output SB_T0_EAST_SB_IN_B17_ready_out,
    input SB_T0_EAST_SB_IN_B17_valid_in,
    output [16:0] SB_T0_EAST_SB_OUT_B17,
    output SB_T0_EAST_SB_OUT_B17_enable,
    input SB_T0_EAST_SB_OUT_B17_ready_in,
    output SB_T0_EAST_SB_OUT_B17_valid_out,
    input [16:0] SB_T0_NORTH_SB_IN_B17,
    output SB_T0_NORTH_SB_IN_B17_enable,
    output SB_T0_NORTH_SB_IN_B17_ready_out,
    input SB_T0_NORTH_SB_IN_B17_valid_in,
    output [16:0] SB_T0_NORTH_SB_OUT_B17,
    output SB_T0_NORTH_SB_OUT_B17_enable,
    input SB_T0_NORTH_SB_OUT_B17_ready_in,
    output SB_T0_NORTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T0_SOUTH_SB_IN_B17,
    output SB_T0_SOUTH_SB_IN_B17_enable,
    output SB_T0_SOUTH_SB_IN_B17_ready_out,
    input SB_T0_SOUTH_SB_IN_B17_valid_in,
    output [16:0] SB_T0_SOUTH_SB_OUT_B17,
    output SB_T0_SOUTH_SB_OUT_B17_enable,
    input SB_T0_SOUTH_SB_OUT_B17_ready_in,
    output SB_T0_SOUTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T0_WEST_SB_IN_B17,
    output SB_T0_WEST_SB_IN_B17_enable,
    output SB_T0_WEST_SB_IN_B17_ready_out,
    input SB_T0_WEST_SB_IN_B17_valid_in,
    output [16:0] SB_T0_WEST_SB_OUT_B17,
    output SB_T0_WEST_SB_OUT_B17_enable,
    input SB_T0_WEST_SB_OUT_B17_ready_in,
    output SB_T0_WEST_SB_OUT_B17_valid_out,
    input [16:0] SB_T1_EAST_SB_IN_B17,
    output SB_T1_EAST_SB_IN_B17_enable,
    output SB_T1_EAST_SB_IN_B17_ready_out,
    input SB_T1_EAST_SB_IN_B17_valid_in,
    output [16:0] SB_T1_EAST_SB_OUT_B17,
    output SB_T1_EAST_SB_OUT_B17_enable,
    input SB_T1_EAST_SB_OUT_B17_ready_in,
    output SB_T1_EAST_SB_OUT_B17_valid_out,
    input [16:0] SB_T1_NORTH_SB_IN_B17,
    output SB_T1_NORTH_SB_IN_B17_enable,
    output SB_T1_NORTH_SB_IN_B17_ready_out,
    input SB_T1_NORTH_SB_IN_B17_valid_in,
    output [16:0] SB_T1_NORTH_SB_OUT_B17,
    output SB_T1_NORTH_SB_OUT_B17_enable,
    input SB_T1_NORTH_SB_OUT_B17_ready_in,
    output SB_T1_NORTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T1_SOUTH_SB_IN_B17,
    output SB_T1_SOUTH_SB_IN_B17_enable,
    output SB_T1_SOUTH_SB_IN_B17_ready_out,
    input SB_T1_SOUTH_SB_IN_B17_valid_in,
    output [16:0] SB_T1_SOUTH_SB_OUT_B17,
    output SB_T1_SOUTH_SB_OUT_B17_enable,
    input SB_T1_SOUTH_SB_OUT_B17_ready_in,
    output SB_T1_SOUTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T1_WEST_SB_IN_B17,
    output SB_T1_WEST_SB_IN_B17_enable,
    output SB_T1_WEST_SB_IN_B17_ready_out,
    input SB_T1_WEST_SB_IN_B17_valid_in,
    output [16:0] SB_T1_WEST_SB_OUT_B17,
    output SB_T1_WEST_SB_OUT_B17_enable,
    input SB_T1_WEST_SB_OUT_B17_ready_in,
    output SB_T1_WEST_SB_OUT_B17_valid_out,
    input [16:0] SB_T2_EAST_SB_IN_B17,
    output SB_T2_EAST_SB_IN_B17_enable,
    output SB_T2_EAST_SB_IN_B17_ready_out,
    input SB_T2_EAST_SB_IN_B17_valid_in,
    output [16:0] SB_T2_EAST_SB_OUT_B17,
    output SB_T2_EAST_SB_OUT_B17_enable,
    input SB_T2_EAST_SB_OUT_B17_ready_in,
    output SB_T2_EAST_SB_OUT_B17_valid_out,
    input [16:0] SB_T2_NORTH_SB_IN_B17,
    output SB_T2_NORTH_SB_IN_B17_enable,
    output SB_T2_NORTH_SB_IN_B17_ready_out,
    input SB_T2_NORTH_SB_IN_B17_valid_in,
    output [16:0] SB_T2_NORTH_SB_OUT_B17,
    output SB_T2_NORTH_SB_OUT_B17_enable,
    input SB_T2_NORTH_SB_OUT_B17_ready_in,
    output SB_T2_NORTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T2_SOUTH_SB_IN_B17,
    output SB_T2_SOUTH_SB_IN_B17_enable,
    output SB_T2_SOUTH_SB_IN_B17_ready_out,
    input SB_T2_SOUTH_SB_IN_B17_valid_in,
    output [16:0] SB_T2_SOUTH_SB_OUT_B17,
    output SB_T2_SOUTH_SB_OUT_B17_enable,
    input SB_T2_SOUTH_SB_OUT_B17_ready_in,
    output SB_T2_SOUTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T2_WEST_SB_IN_B17,
    output SB_T2_WEST_SB_IN_B17_enable,
    output SB_T2_WEST_SB_IN_B17_ready_out,
    input SB_T2_WEST_SB_IN_B17_valid_in,
    output [16:0] SB_T2_WEST_SB_OUT_B17,
    output SB_T2_WEST_SB_OUT_B17_enable,
    input SB_T2_WEST_SB_OUT_B17_ready_in,
    output SB_T2_WEST_SB_OUT_B17_valid_out,
    input [16:0] SB_T3_EAST_SB_IN_B17,
    output SB_T3_EAST_SB_IN_B17_enable,
    output SB_T3_EAST_SB_IN_B17_ready_out,
    input SB_T3_EAST_SB_IN_B17_valid_in,
    output [16:0] SB_T3_EAST_SB_OUT_B17,
    output SB_T3_EAST_SB_OUT_B17_enable,
    input SB_T3_EAST_SB_OUT_B17_ready_in,
    output SB_T3_EAST_SB_OUT_B17_valid_out,
    input [16:0] SB_T3_NORTH_SB_IN_B17,
    output SB_T3_NORTH_SB_IN_B17_enable,
    output SB_T3_NORTH_SB_IN_B17_ready_out,
    input SB_T3_NORTH_SB_IN_B17_valid_in,
    output [16:0] SB_T3_NORTH_SB_OUT_B17,
    output SB_T3_NORTH_SB_OUT_B17_enable,
    input SB_T3_NORTH_SB_OUT_B17_ready_in,
    output SB_T3_NORTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T3_SOUTH_SB_IN_B17,
    output SB_T3_SOUTH_SB_IN_B17_enable,
    output SB_T3_SOUTH_SB_IN_B17_ready_out,
    input SB_T3_SOUTH_SB_IN_B17_valid_in,
    output [16:0] SB_T3_SOUTH_SB_OUT_B17,
    output SB_T3_SOUTH_SB_OUT_B17_enable,
    input SB_T3_SOUTH_SB_OUT_B17_ready_in,
    output SB_T3_SOUTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T3_WEST_SB_IN_B17,
    output SB_T3_WEST_SB_IN_B17_enable,
    output SB_T3_WEST_SB_IN_B17_ready_out,
    input SB_T3_WEST_SB_IN_B17_valid_in,
    output [16:0] SB_T3_WEST_SB_OUT_B17,
    output SB_T3_WEST_SB_OUT_B17_enable,
    input SB_T3_WEST_SB_OUT_B17_ready_in,
    output SB_T3_WEST_SB_OUT_B17_valid_out,
    input [16:0] SB_T4_EAST_SB_IN_B17,
    output SB_T4_EAST_SB_IN_B17_enable,
    output SB_T4_EAST_SB_IN_B17_ready_out,
    input SB_T4_EAST_SB_IN_B17_valid_in,
    output [16:0] SB_T4_EAST_SB_OUT_B17,
    output SB_T4_EAST_SB_OUT_B17_enable,
    input SB_T4_EAST_SB_OUT_B17_ready_in,
    output SB_T4_EAST_SB_OUT_B17_valid_out,
    input [16:0] SB_T4_NORTH_SB_IN_B17,
    output SB_T4_NORTH_SB_IN_B17_enable,
    output SB_T4_NORTH_SB_IN_B17_ready_out,
    input SB_T4_NORTH_SB_IN_B17_valid_in,
    output [16:0] SB_T4_NORTH_SB_OUT_B17,
    output SB_T4_NORTH_SB_OUT_B17_enable,
    input SB_T4_NORTH_SB_OUT_B17_ready_in,
    output SB_T4_NORTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T4_SOUTH_SB_IN_B17,
    output SB_T4_SOUTH_SB_IN_B17_enable,
    output SB_T4_SOUTH_SB_IN_B17_ready_out,
    input SB_T4_SOUTH_SB_IN_B17_valid_in,
    output [16:0] SB_T4_SOUTH_SB_OUT_B17,
    output SB_T4_SOUTH_SB_OUT_B17_enable,
    input SB_T4_SOUTH_SB_OUT_B17_ready_in,
    output SB_T4_SOUTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T4_WEST_SB_IN_B17,
    output SB_T4_WEST_SB_IN_B17_enable,
    output SB_T4_WEST_SB_IN_B17_ready_out,
    input SB_T4_WEST_SB_IN_B17_valid_in,
    output [16:0] SB_T4_WEST_SB_OUT_B17,
    output SB_T4_WEST_SB_OUT_B17_enable,
    input SB_T4_WEST_SB_OUT_B17_ready_in,
    output SB_T4_WEST_SB_OUT_B17_valid_out,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset,
    input [0:0] stall
);
wire [0:0] CB_PE_output_width_17_num_0_fan_in_O;
wire [0:0] CB_PE_output_width_17_num_1_fan_in_O;
wire [0:0] CB_PE_output_width_17_num_2_fan_in_O;
wire [0:0] CB_PondTop_output_width_17_num_0_fan_in_O;
wire [0:0] CB_PondTop_output_width_17_num_1_fan_in_O;
wire [0:0] Invert1_inst0_out;
wire [16:0] MUX_SB_T0_EAST_SB_OUT_B17_O;
wire MUX_SB_T0_EAST_SB_OUT_B17_ready_out;
wire MUX_SB_T0_EAST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T0_EAST_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T0_NORTH_SB_OUT_B17_O;
wire MUX_SB_T0_NORTH_SB_OUT_B17_ready_out;
wire MUX_SB_T0_NORTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T0_NORTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T0_SOUTH_SB_OUT_B17_O;
wire MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out;
wire MUX_SB_T0_SOUTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T0_WEST_SB_OUT_B17_O;
wire MUX_SB_T0_WEST_SB_OUT_B17_ready_out;
wire MUX_SB_T0_WEST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T0_WEST_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T1_EAST_SB_OUT_B17_O;
wire MUX_SB_T1_EAST_SB_OUT_B17_ready_out;
wire MUX_SB_T1_EAST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T1_EAST_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T1_NORTH_SB_OUT_B17_O;
wire MUX_SB_T1_NORTH_SB_OUT_B17_ready_out;
wire MUX_SB_T1_NORTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T1_NORTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T1_SOUTH_SB_OUT_B17_O;
wire MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out;
wire MUX_SB_T1_SOUTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T1_WEST_SB_OUT_B17_O;
wire MUX_SB_T1_WEST_SB_OUT_B17_ready_out;
wire MUX_SB_T1_WEST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T1_WEST_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T2_EAST_SB_OUT_B17_O;
wire MUX_SB_T2_EAST_SB_OUT_B17_ready_out;
wire MUX_SB_T2_EAST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T2_EAST_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T2_NORTH_SB_OUT_B17_O;
wire MUX_SB_T2_NORTH_SB_OUT_B17_ready_out;
wire MUX_SB_T2_NORTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T2_NORTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T2_SOUTH_SB_OUT_B17_O;
wire MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out;
wire MUX_SB_T2_SOUTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T2_WEST_SB_OUT_B17_O;
wire MUX_SB_T2_WEST_SB_OUT_B17_ready_out;
wire MUX_SB_T2_WEST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T2_WEST_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T3_EAST_SB_OUT_B17_O;
wire MUX_SB_T3_EAST_SB_OUT_B17_ready_out;
wire MUX_SB_T3_EAST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T3_EAST_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T3_NORTH_SB_OUT_B17_O;
wire MUX_SB_T3_NORTH_SB_OUT_B17_ready_out;
wire MUX_SB_T3_NORTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T3_NORTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T3_SOUTH_SB_OUT_B17_O;
wire MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out;
wire MUX_SB_T3_SOUTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T3_WEST_SB_OUT_B17_O;
wire MUX_SB_T3_WEST_SB_OUT_B17_ready_out;
wire MUX_SB_T3_WEST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T3_WEST_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T4_EAST_SB_OUT_B17_O;
wire MUX_SB_T4_EAST_SB_OUT_B17_ready_out;
wire MUX_SB_T4_EAST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T4_EAST_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T4_NORTH_SB_OUT_B17_O;
wire MUX_SB_T4_NORTH_SB_OUT_B17_ready_out;
wire MUX_SB_T4_NORTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T4_NORTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T4_SOUTH_SB_OUT_B17_O;
wire MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out;
wire MUX_SB_T4_SOUTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T4_WEST_SB_OUT_B17_O;
wire MUX_SB_T4_WEST_SB_OUT_B17_ready_out;
wire MUX_SB_T4_WEST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T4_WEST_SB_OUT_B17_out_sel;
wire [0:0] REG_T0_EAST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T0_EAST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T0_EAST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T0_EAST_B17_end_value_O;
wire [0:0] REG_T0_EAST_B17_fifo_value_O;
wire [0:0] REG_T0_EAST_B17_start_value_O;
wire [0:0] REG_T0_NORTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T0_NORTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T0_NORTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T0_NORTH_B17_end_value_O;
wire [0:0] REG_T0_NORTH_B17_fifo_value_O;
wire [0:0] REG_T0_NORTH_B17_start_value_O;
wire [0:0] REG_T0_SOUTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T0_SOUTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T0_SOUTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T0_SOUTH_B17_end_value_O;
wire [0:0] REG_T0_SOUTH_B17_fifo_value_O;
wire [0:0] REG_T0_SOUTH_B17_start_value_O;
wire [0:0] REG_T0_WEST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T0_WEST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T0_WEST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T0_WEST_B17_end_value_O;
wire [0:0] REG_T0_WEST_B17_fifo_value_O;
wire [0:0] REG_T0_WEST_B17_start_value_O;
wire [0:0] REG_T1_EAST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T1_EAST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T1_EAST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T1_EAST_B17_end_value_O;
wire [0:0] REG_T1_EAST_B17_fifo_value_O;
wire [0:0] REG_T1_EAST_B17_start_value_O;
wire [0:0] REG_T1_NORTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T1_NORTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T1_NORTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T1_NORTH_B17_end_value_O;
wire [0:0] REG_T1_NORTH_B17_fifo_value_O;
wire [0:0] REG_T1_NORTH_B17_start_value_O;
wire [0:0] REG_T1_SOUTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T1_SOUTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T1_SOUTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T1_SOUTH_B17_end_value_O;
wire [0:0] REG_T1_SOUTH_B17_fifo_value_O;
wire [0:0] REG_T1_SOUTH_B17_start_value_O;
wire [0:0] REG_T1_WEST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T1_WEST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T1_WEST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T1_WEST_B17_end_value_O;
wire [0:0] REG_T1_WEST_B17_fifo_value_O;
wire [0:0] REG_T1_WEST_B17_start_value_O;
wire [0:0] REG_T2_EAST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T2_EAST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T2_EAST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T2_EAST_B17_end_value_O;
wire [0:0] REG_T2_EAST_B17_fifo_value_O;
wire [0:0] REG_T2_EAST_B17_start_value_O;
wire [0:0] REG_T2_NORTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T2_NORTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T2_NORTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T2_NORTH_B17_end_value_O;
wire [0:0] REG_T2_NORTH_B17_fifo_value_O;
wire [0:0] REG_T2_NORTH_B17_start_value_O;
wire [0:0] REG_T2_SOUTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T2_SOUTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T2_SOUTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T2_SOUTH_B17_end_value_O;
wire [0:0] REG_T2_SOUTH_B17_fifo_value_O;
wire [0:0] REG_T2_SOUTH_B17_start_value_O;
wire [0:0] REG_T2_WEST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T2_WEST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T2_WEST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T2_WEST_B17_end_value_O;
wire [0:0] REG_T2_WEST_B17_fifo_value_O;
wire [0:0] REG_T2_WEST_B17_start_value_O;
wire [0:0] REG_T3_EAST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T3_EAST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T3_EAST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T3_EAST_B17_end_value_O;
wire [0:0] REG_T3_EAST_B17_fifo_value_O;
wire [0:0] REG_T3_EAST_B17_start_value_O;
wire [0:0] REG_T3_NORTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T3_NORTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T3_NORTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T3_NORTH_B17_end_value_O;
wire [0:0] REG_T3_NORTH_B17_fifo_value_O;
wire [0:0] REG_T3_NORTH_B17_start_value_O;
wire [0:0] REG_T3_SOUTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T3_SOUTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T3_SOUTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T3_SOUTH_B17_end_value_O;
wire [0:0] REG_T3_SOUTH_B17_fifo_value_O;
wire [0:0] REG_T3_SOUTH_B17_start_value_O;
wire [0:0] REG_T3_WEST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T3_WEST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T3_WEST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T3_WEST_B17_end_value_O;
wire [0:0] REG_T3_WEST_B17_fifo_value_O;
wire [0:0] REG_T3_WEST_B17_start_value_O;
wire [0:0] REG_T4_EAST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T4_EAST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T4_EAST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T4_EAST_B17_end_value_O;
wire [0:0] REG_T4_EAST_B17_fifo_value_O;
wire [0:0] REG_T4_EAST_B17_start_value_O;
wire [0:0] REG_T4_NORTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T4_NORTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T4_NORTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T4_NORTH_B17_end_value_O;
wire [0:0] REG_T4_NORTH_B17_fifo_value_O;
wire [0:0] REG_T4_NORTH_B17_start_value_O;
wire [0:0] REG_T4_SOUTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T4_SOUTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T4_SOUTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T4_SOUTH_B17_end_value_O;
wire [0:0] REG_T4_SOUTH_B17_fifo_value_O;
wire [0:0] REG_T4_SOUTH_B17_start_value_O;
wire [0:0] REG_T4_WEST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T4_WEST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T4_WEST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T4_WEST_B17_end_value_O;
wire [0:0] REG_T4_WEST_B17_fifo_value_O;
wire [0:0] REG_T4_WEST_B17_start_value_O;
wire [16:0] RMUX_T0_EAST_B17_O;
wire RMUX_T0_EAST_B17_ready_out;
wire RMUX_T0_EAST_B17_valid_out;
wire [1:0] RMUX_T0_EAST_B17_out_sel;
wire [0:0] RMUX_T0_EAST_B17_sel_value_O;
wire [16:0] RMUX_T0_NORTH_B17_O;
wire RMUX_T0_NORTH_B17_ready_out;
wire RMUX_T0_NORTH_B17_valid_out;
wire [1:0] RMUX_T0_NORTH_B17_out_sel;
wire [0:0] RMUX_T0_NORTH_B17_sel_value_O;
wire [16:0] RMUX_T0_SOUTH_B17_O;
wire RMUX_T0_SOUTH_B17_ready_out;
wire RMUX_T0_SOUTH_B17_valid_out;
wire [1:0] RMUX_T0_SOUTH_B17_out_sel;
wire [0:0] RMUX_T0_SOUTH_B17_sel_value_O;
wire [16:0] RMUX_T0_WEST_B17_O;
wire RMUX_T0_WEST_B17_ready_out;
wire RMUX_T0_WEST_B17_valid_out;
wire [1:0] RMUX_T0_WEST_B17_out_sel;
wire [0:0] RMUX_T0_WEST_B17_sel_value_O;
wire [16:0] RMUX_T1_EAST_B17_O;
wire RMUX_T1_EAST_B17_ready_out;
wire RMUX_T1_EAST_B17_valid_out;
wire [1:0] RMUX_T1_EAST_B17_out_sel;
wire [0:0] RMUX_T1_EAST_B17_sel_value_O;
wire [16:0] RMUX_T1_NORTH_B17_O;
wire RMUX_T1_NORTH_B17_ready_out;
wire RMUX_T1_NORTH_B17_valid_out;
wire [1:0] RMUX_T1_NORTH_B17_out_sel;
wire [0:0] RMUX_T1_NORTH_B17_sel_value_O;
wire [16:0] RMUX_T1_SOUTH_B17_O;
wire RMUX_T1_SOUTH_B17_ready_out;
wire RMUX_T1_SOUTH_B17_valid_out;
wire [1:0] RMUX_T1_SOUTH_B17_out_sel;
wire [0:0] RMUX_T1_SOUTH_B17_sel_value_O;
wire [16:0] RMUX_T1_WEST_B17_O;
wire RMUX_T1_WEST_B17_ready_out;
wire RMUX_T1_WEST_B17_valid_out;
wire [1:0] RMUX_T1_WEST_B17_out_sel;
wire [0:0] RMUX_T1_WEST_B17_sel_value_O;
wire [16:0] RMUX_T2_EAST_B17_O;
wire RMUX_T2_EAST_B17_ready_out;
wire RMUX_T2_EAST_B17_valid_out;
wire [1:0] RMUX_T2_EAST_B17_out_sel;
wire [0:0] RMUX_T2_EAST_B17_sel_value_O;
wire [16:0] RMUX_T2_NORTH_B17_O;
wire RMUX_T2_NORTH_B17_ready_out;
wire RMUX_T2_NORTH_B17_valid_out;
wire [1:0] RMUX_T2_NORTH_B17_out_sel;
wire [0:0] RMUX_T2_NORTH_B17_sel_value_O;
wire [16:0] RMUX_T2_SOUTH_B17_O;
wire RMUX_T2_SOUTH_B17_ready_out;
wire RMUX_T2_SOUTH_B17_valid_out;
wire [1:0] RMUX_T2_SOUTH_B17_out_sel;
wire [0:0] RMUX_T2_SOUTH_B17_sel_value_O;
wire [16:0] RMUX_T2_WEST_B17_O;
wire RMUX_T2_WEST_B17_ready_out;
wire RMUX_T2_WEST_B17_valid_out;
wire [1:0] RMUX_T2_WEST_B17_out_sel;
wire [0:0] RMUX_T2_WEST_B17_sel_value_O;
wire [16:0] RMUX_T3_EAST_B17_O;
wire RMUX_T3_EAST_B17_ready_out;
wire RMUX_T3_EAST_B17_valid_out;
wire [1:0] RMUX_T3_EAST_B17_out_sel;
wire [0:0] RMUX_T3_EAST_B17_sel_value_O;
wire [16:0] RMUX_T3_NORTH_B17_O;
wire RMUX_T3_NORTH_B17_ready_out;
wire RMUX_T3_NORTH_B17_valid_out;
wire [1:0] RMUX_T3_NORTH_B17_out_sel;
wire [0:0] RMUX_T3_NORTH_B17_sel_value_O;
wire [16:0] RMUX_T3_SOUTH_B17_O;
wire RMUX_T3_SOUTH_B17_ready_out;
wire RMUX_T3_SOUTH_B17_valid_out;
wire [1:0] RMUX_T3_SOUTH_B17_out_sel;
wire [0:0] RMUX_T3_SOUTH_B17_sel_value_O;
wire [16:0] RMUX_T3_WEST_B17_O;
wire RMUX_T3_WEST_B17_ready_out;
wire RMUX_T3_WEST_B17_valid_out;
wire [1:0] RMUX_T3_WEST_B17_out_sel;
wire [0:0] RMUX_T3_WEST_B17_sel_value_O;
wire [16:0] RMUX_T4_EAST_B17_O;
wire RMUX_T4_EAST_B17_ready_out;
wire RMUX_T4_EAST_B17_valid_out;
wire [1:0] RMUX_T4_EAST_B17_out_sel;
wire [0:0] RMUX_T4_EAST_B17_sel_value_O;
wire [16:0] RMUX_T4_NORTH_B17_O;
wire RMUX_T4_NORTH_B17_ready_out;
wire RMUX_T4_NORTH_B17_valid_out;
wire [1:0] RMUX_T4_NORTH_B17_out_sel;
wire [0:0] RMUX_T4_NORTH_B17_sel_value_O;
wire [16:0] RMUX_T4_SOUTH_B17_O;
wire RMUX_T4_SOUTH_B17_ready_out;
wire RMUX_T4_SOUTH_B17_valid_out;
wire [1:0] RMUX_T4_SOUTH_B17_out_sel;
wire [0:0] RMUX_T4_SOUTH_B17_sel_value_O;
wire [16:0] RMUX_T4_WEST_B17_O;
wire RMUX_T4_WEST_B17_ready_out;
wire RMUX_T4_WEST_B17_valid_out;
wire [1:0] RMUX_T4_WEST_B17_out_sel;
wire [0:0] RMUX_T4_WEST_B17_sel_value_O;
wire [0:0] SB_T0_EAST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T0_EAST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T0_EAST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T0_EAST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T0_EAST_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T0_NORTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T0_NORTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T0_NORTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T0_NORTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T0_NORTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T0_SOUTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T0_SOUTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T0_SOUTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T0_SOUTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T0_SOUTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T0_WEST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T0_WEST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T0_WEST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T0_WEST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T0_WEST_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T1_EAST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T1_EAST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T1_EAST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T1_EAST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T1_EAST_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T1_NORTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T1_NORTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T1_NORTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T1_NORTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T1_NORTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T1_SOUTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T1_SOUTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T1_SOUTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T1_SOUTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T1_SOUTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T1_WEST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T1_WEST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T1_WEST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T1_WEST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T1_WEST_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T2_EAST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T2_EAST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T2_EAST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T2_EAST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T2_EAST_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T2_NORTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T2_NORTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T2_NORTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T2_NORTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T2_NORTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T2_SOUTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T2_SOUTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T2_SOUTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T2_SOUTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T2_SOUTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T2_WEST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T2_WEST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T2_WEST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T2_WEST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T2_WEST_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T3_EAST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T3_EAST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T3_EAST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T3_EAST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T3_EAST_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T3_NORTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T3_NORTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T3_NORTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T3_NORTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T3_NORTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T3_SOUTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T3_SOUTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T3_SOUTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T3_SOUTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T3_SOUTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T3_WEST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T3_WEST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T3_WEST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T3_WEST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T3_WEST_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T4_EAST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T4_EAST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T4_EAST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T4_EAST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T4_EAST_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T4_NORTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T4_NORTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T4_NORTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T4_NORTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T4_NORTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T4_SOUTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T4_SOUTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T4_SOUTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T4_SOUTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T4_SOUTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T4_WEST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T4_WEST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T4_WEST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T4_WEST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T4_WEST_SB_OUT_B17_sel_value_O;
wire [16:0] WIRE_SB_T0_EAST_SB_IN_B17_O;
wire WIRE_SB_T0_EAST_SB_IN_B17_ready_out;
wire WIRE_SB_T0_EAST_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T0_NORTH_SB_IN_B17_O;
wire WIRE_SB_T0_NORTH_SB_IN_B17_ready_out;
wire WIRE_SB_T0_NORTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T0_SOUTH_SB_IN_B17_O;
wire WIRE_SB_T0_SOUTH_SB_IN_B17_ready_out;
wire WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T0_WEST_SB_IN_B17_O;
wire WIRE_SB_T0_WEST_SB_IN_B17_ready_out;
wire WIRE_SB_T0_WEST_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T1_EAST_SB_IN_B17_O;
wire WIRE_SB_T1_EAST_SB_IN_B17_ready_out;
wire WIRE_SB_T1_EAST_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T1_NORTH_SB_IN_B17_O;
wire WIRE_SB_T1_NORTH_SB_IN_B17_ready_out;
wire WIRE_SB_T1_NORTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T1_SOUTH_SB_IN_B17_O;
wire WIRE_SB_T1_SOUTH_SB_IN_B17_ready_out;
wire WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T1_WEST_SB_IN_B17_O;
wire WIRE_SB_T1_WEST_SB_IN_B17_ready_out;
wire WIRE_SB_T1_WEST_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T2_EAST_SB_IN_B17_O;
wire WIRE_SB_T2_EAST_SB_IN_B17_ready_out;
wire WIRE_SB_T2_EAST_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T2_NORTH_SB_IN_B17_O;
wire WIRE_SB_T2_NORTH_SB_IN_B17_ready_out;
wire WIRE_SB_T2_NORTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T2_SOUTH_SB_IN_B17_O;
wire WIRE_SB_T2_SOUTH_SB_IN_B17_ready_out;
wire WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T2_WEST_SB_IN_B17_O;
wire WIRE_SB_T2_WEST_SB_IN_B17_ready_out;
wire WIRE_SB_T2_WEST_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T3_EAST_SB_IN_B17_O;
wire WIRE_SB_T3_EAST_SB_IN_B17_ready_out;
wire WIRE_SB_T3_EAST_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T3_NORTH_SB_IN_B17_O;
wire WIRE_SB_T3_NORTH_SB_IN_B17_ready_out;
wire WIRE_SB_T3_NORTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T3_SOUTH_SB_IN_B17_O;
wire WIRE_SB_T3_SOUTH_SB_IN_B17_ready_out;
wire WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T3_WEST_SB_IN_B17_O;
wire WIRE_SB_T3_WEST_SB_IN_B17_ready_out;
wire WIRE_SB_T3_WEST_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T4_EAST_SB_IN_B17_O;
wire WIRE_SB_T4_EAST_SB_IN_B17_ready_out;
wire WIRE_SB_T4_EAST_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T4_NORTH_SB_IN_B17_O;
wire WIRE_SB_T4_NORTH_SB_IN_B17_ready_out;
wire WIRE_SB_T4_NORTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T4_SOUTH_SB_IN_B17_O;
wire WIRE_SB_T4_SOUTH_SB_IN_B17_ready_out;
wire WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T4_WEST_SB_IN_B17_O;
wire WIRE_SB_T4_WEST_SB_IN_B17_ready_out;
wire WIRE_SB_T4_WEST_SB_IN_B17_valid_out;
wire ZextWrapper_23_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_23_32_inst0$self_O_in;
wire ZextWrapper_30_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_30_32_inst0$self_O_in;
wire ZextWrapper_31_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_31_32_inst0$self_O_in;
wire [0:0] and1_inst0_out;
wire [0:0] and1_inst1_out;
wire [0:0] and1_inst10_out;
wire [0:0] and1_inst11_out;
wire [0:0] and1_inst12_out;
wire [0:0] and1_inst13_out;
wire [0:0] and1_inst14_out;
wire [0:0] and1_inst15_out;
wire [0:0] and1_inst16_out;
wire [0:0] and1_inst17_out;
wire [0:0] and1_inst18_out;
wire [0:0] and1_inst19_out;
wire [0:0] and1_inst2_out;
wire [0:0] and1_inst3_out;
wire [0:0] and1_inst4_out;
wire [0:0] and1_inst5_out;
wire [0:0] and1_inst6_out;
wire [0:0] and1_inst7_out;
wire [0:0] and1_inst8_out;
wire [0:0] and1_inst9_out;
wire [31:0] config_reg_0_O;
wire [31:0] config_reg_1_O;
wire [31:0] config_reg_2_O;
wire [30:0] config_reg_3_O;
wire [29:0] config_reg_4_O;
wire [22:0] config_reg_5_O;
wire [0:0] const_1_1_out;
wire coreir_eq_1_inst0_out;
wire coreir_eq_1_inst1_out;
wire coreir_eq_1_inst10_out;
wire coreir_eq_1_inst11_out;
wire coreir_eq_1_inst12_out;
wire coreir_eq_1_inst13_out;
wire coreir_eq_1_inst14_out;
wire coreir_eq_1_inst15_out;
wire coreir_eq_1_inst16_out;
wire coreir_eq_1_inst17_out;
wire coreir_eq_1_inst18_out;
wire coreir_eq_1_inst19_out;
wire coreir_eq_1_inst2_out;
wire coreir_eq_1_inst3_out;
wire coreir_eq_1_inst4_out;
wire coreir_eq_1_inst5_out;
wire coreir_eq_1_inst6_out;
wire coreir_eq_1_inst7_out;
wire coreir_eq_1_inst8_out;
wire coreir_eq_1_inst9_out;
wire [31:0] mux_aoi_6_32_inst0_O;
wire [7:0] mux_aoi_6_32_inst0_out_sel;
wire [7:0] self_config_config_addr_out;
FanoutHash_330DF95D65589621 CB_PE_output_width_17_num_0_fan_in (
    .S13(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
    .E13(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
    .S6(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
    .E2(SB_T0_EAST_SB_OUT_B17_enable_value_O),
    .E12(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
    .E7(SB_T1_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
    .E18(SB_T4_EAST_SB_OUT_B17_enable_value_O),
    .I3(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
    .E19(SB_T4_WEST_SB_OUT_B17_enable_value_O),
    .I14(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
    .S14(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
    .I9(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
    .S12(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
    .E20(PondTop_input_width_17_num_0_enable),
    .S17(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
    .I21(PondTop_input_width_17_num_1_ready),
    .S21(PondTop_input_width_17_num_1_out_sel),
    .I13(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
    .S9(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
    .E10(SB_T2_EAST_SB_OUT_B17_enable_value_O),
    .E15(SB_T3_WEST_SB_OUT_B17_enable_value_O),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
    .E5(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
    .S10(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
    .E8(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
    .I11(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
    .I6(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
    .S15(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
    .I20(PondTop_input_width_17_num_0_ready),
    .S20(PondTop_input_width_17_num_0_out_sel),
    .E21(PondTop_input_width_17_num_1_enable),
    .I7(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
    .E14(SB_T3_EAST_SB_OUT_B17_enable_value_O),
    .I2(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
    .E11(SB_T2_WEST_SB_OUT_B17_enable_value_O),
    .S3(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
    .S8(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
    .I10(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
    .S16(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
    .E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
    .E16(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
    .E3(SB_T0_WEST_SB_OUT_B17_enable_value_O),
    .S18(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
    .S19(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
    .S2(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
    .S4(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
    .E9(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
    .I16(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
    .I12(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
    .S11(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
    .I17(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
    .I19(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
    .I18(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
    .S7(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
    .E4(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
    .E17(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
    .S5(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
    .I1(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
    .I5(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
    .E6(SB_T1_EAST_SB_OUT_B17_enable_value_O),
    .I4(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
    .I8(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
    .O(CB_PE_output_width_17_num_0_fan_in_O),
    .E1(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
    .I15(MUX_SB_T3_WEST_SB_OUT_B17_ready_out)
);
FanoutHash_82899D6851EDC11 CB_PE_output_width_17_num_1_fan_in (
    .S13(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
    .E13(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
    .S6(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
    .E2(SB_T0_EAST_SB_OUT_B17_enable_value_O),
    .E12(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
    .E7(SB_T1_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
    .E18(SB_T4_EAST_SB_OUT_B17_enable_value_O),
    .I3(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
    .E19(SB_T4_WEST_SB_OUT_B17_enable_value_O),
    .I14(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
    .S14(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
    .I9(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
    .S12(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
    .S17(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
    .I13(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
    .S9(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
    .E10(SB_T2_EAST_SB_OUT_B17_enable_value_O),
    .E15(SB_T3_WEST_SB_OUT_B17_enable_value_O),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
    .E5(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
    .S10(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
    .E8(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
    .I11(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
    .I6(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
    .S15(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
    .I7(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
    .E14(SB_T3_EAST_SB_OUT_B17_enable_value_O),
    .I2(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
    .E11(SB_T2_WEST_SB_OUT_B17_enable_value_O),
    .S3(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
    .S8(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
    .I10(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
    .S16(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
    .E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
    .E16(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
    .E3(SB_T0_WEST_SB_OUT_B17_enable_value_O),
    .S18(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
    .S19(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
    .S2(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
    .S4(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
    .E9(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
    .I16(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
    .I12(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
    .S11(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
    .I17(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
    .I19(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
    .I18(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
    .S7(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
    .E4(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
    .E17(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
    .S5(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
    .I1(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
    .I5(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
    .E6(SB_T1_EAST_SB_OUT_B17_enable_value_O),
    .I4(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
    .I8(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
    .O(CB_PE_output_width_17_num_1_fan_in_O),
    .E1(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
    .I15(MUX_SB_T3_WEST_SB_OUT_B17_ready_out)
);
FanoutHash_CE1AA874B742213 CB_PE_output_width_17_num_2_fan_in (
    .S13(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
    .E13(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
    .S6(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
    .E2(SB_T0_EAST_SB_OUT_B17_enable_value_O),
    .E12(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
    .E7(SB_T1_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
    .E18(SB_T4_EAST_SB_OUT_B17_enable_value_O),
    .I3(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
    .E19(SB_T4_WEST_SB_OUT_B17_enable_value_O),
    .I14(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
    .S14(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
    .I9(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
    .S12(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
    .S17(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
    .I13(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
    .S9(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
    .E10(SB_T2_EAST_SB_OUT_B17_enable_value_O),
    .E15(SB_T3_WEST_SB_OUT_B17_enable_value_O),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
    .E5(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
    .S10(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
    .E8(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
    .I11(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
    .I6(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
    .S15(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
    .I7(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
    .E14(SB_T3_EAST_SB_OUT_B17_enable_value_O),
    .I2(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
    .E11(SB_T2_WEST_SB_OUT_B17_enable_value_O),
    .S3(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
    .S8(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
    .I10(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
    .S16(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
    .E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
    .E16(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
    .E3(SB_T0_WEST_SB_OUT_B17_enable_value_O),
    .S18(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
    .S19(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
    .S2(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
    .S4(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
    .E9(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
    .I16(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
    .I12(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
    .S11(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
    .I17(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
    .I19(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
    .I18(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
    .S7(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
    .E4(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
    .E17(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
    .S5(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
    .I1(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
    .I5(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
    .E6(SB_T1_EAST_SB_OUT_B17_enable_value_O),
    .I4(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
    .I8(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
    .O(CB_PE_output_width_17_num_2_fan_in_O),
    .E1(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
    .I15(MUX_SB_T3_WEST_SB_OUT_B17_ready_out)
);
FanoutHash_14EBE1E8E49CA541 CB_PondTop_output_width_17_num_0_fan_in (
    .I2(PE_input_width_17_num_2_ready),
    .E2(PE_input_width_17_num_2_enable),
    .S1(PE_input_width_17_num_1_out_sel),
    .I1(PE_input_width_17_num_1_ready),
    .E0(PE_input_width_17_num_0_enable),
    .S2(PE_input_width_17_num_2_out_sel),
    .S0(PE_input_width_17_num_0_out_sel),
    .O(CB_PondTop_output_width_17_num_0_fan_in_O),
    .E1(PE_input_width_17_num_1_enable),
    .I0(PE_input_width_17_num_0_ready)
);
FanoutHash_1EBD0270673B29D7 CB_PondTop_output_width_17_num_1_fan_in (
    .S13(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
    .E13(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
    .S6(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
    .E2(SB_T0_EAST_SB_OUT_B17_enable_value_O),
    .E12(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
    .E7(SB_T1_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
    .E18(SB_T4_EAST_SB_OUT_B17_enable_value_O),
    .I3(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
    .E19(SB_T4_WEST_SB_OUT_B17_enable_value_O),
    .I14(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
    .S14(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
    .I9(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
    .S12(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
    .S17(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
    .I13(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
    .S9(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
    .E10(SB_T2_EAST_SB_OUT_B17_enable_value_O),
    .E15(SB_T3_WEST_SB_OUT_B17_enable_value_O),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
    .E5(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
    .S10(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
    .E8(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
    .I11(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
    .I6(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
    .S15(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
    .I7(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
    .E14(SB_T3_EAST_SB_OUT_B17_enable_value_O),
    .I2(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
    .E11(SB_T2_WEST_SB_OUT_B17_enable_value_O),
    .S3(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
    .S8(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
    .I10(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
    .S16(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
    .E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
    .E16(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
    .E3(SB_T0_WEST_SB_OUT_B17_enable_value_O),
    .S18(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
    .S19(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
    .S2(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
    .S4(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
    .E9(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
    .I16(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
    .I12(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
    .S11(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
    .I17(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
    .I19(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
    .I18(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
    .S7(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
    .E4(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
    .E17(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
    .S5(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
    .I1(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
    .I5(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
    .E6(SB_T1_EAST_SB_OUT_B17_enable_value_O),
    .I4(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
    .I8(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
    .O(CB_PondTop_output_width_17_num_1_fan_in_O),
    .E1(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
    .I15(MUX_SB_T3_WEST_SB_OUT_B17_ready_out)
);
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(stall),
    .out(Invert1_inst0_out)
);
wire [16:0] MUX_SB_T0_EAST_SB_OUT_B17_I [6:0];
assign MUX_SB_T0_EAST_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T0_EAST_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T0_EAST_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T0_EAST_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T0_EAST_SB_OUT_B17_I[2] = WIRE_SB_T4_NORTH_SB_IN_B17_O;
assign MUX_SB_T0_EAST_SB_OUT_B17_I[1] = WIRE_SB_T3_SOUTH_SB_IN_B17_O;
assign MUX_SB_T0_EAST_SB_OUT_B17_I[0] = WIRE_SB_T0_WEST_SB_IN_B17_O;
wire [6:0] MUX_SB_T0_EAST_SB_OUT_B17_valid_in;
assign MUX_SB_T0_EAST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T4_NORTH_SB_IN_B17_valid_out,WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T0_WEST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T0_EAST_SB_OUT_B17 (
    .I(MUX_SB_T0_EAST_SB_OUT_B17_I),
    .O(MUX_SB_T0_EAST_SB_OUT_B17_O),
    .ready_in(SB_T0_EAST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T0_EAST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T0_EAST_SB_OUT_B17_valid_out),
    .S(SB_T0_EAST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T0_EAST_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T0_NORTH_SB_OUT_B17_I [6:0];
assign MUX_SB_T0_NORTH_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T0_NORTH_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T0_NORTH_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T0_NORTH_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T0_NORTH_SB_OUT_B17_I[2] = WIRE_SB_T0_SOUTH_SB_IN_B17_O;
assign MUX_SB_T0_NORTH_SB_OUT_B17_I[1] = WIRE_SB_T1_EAST_SB_IN_B17_O;
assign MUX_SB_T0_NORTH_SB_OUT_B17_I[0] = WIRE_SB_T0_WEST_SB_IN_B17_O;
wire [6:0] MUX_SB_T0_NORTH_SB_OUT_B17_valid_in;
assign MUX_SB_T0_NORTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T1_EAST_SB_IN_B17_valid_out,WIRE_SB_T0_WEST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T0_NORTH_SB_OUT_B17 (
    .I(MUX_SB_T0_NORTH_SB_OUT_B17_I),
    .O(MUX_SB_T0_NORTH_SB_OUT_B17_O),
    .ready_in(SB_T0_NORTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T0_NORTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T0_NORTH_SB_OUT_B17_valid_out),
    .S(SB_T0_NORTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T0_SOUTH_SB_OUT_B17_I [6:0];
assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[2] = WIRE_SB_T1_WEST_SB_IN_B17_O;
assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[1] = WIRE_SB_T0_NORTH_SB_IN_B17_O;
assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[0] = WIRE_SB_T3_EAST_SB_IN_B17_O;
wire [6:0] MUX_SB_T0_SOUTH_SB_OUT_B17_valid_in;
assign MUX_SB_T0_SOUTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T1_WEST_SB_IN_B17_valid_out,WIRE_SB_T0_NORTH_SB_IN_B17_valid_out,WIRE_SB_T3_EAST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T0_SOUTH_SB_OUT_B17 (
    .I(MUX_SB_T0_SOUTH_SB_OUT_B17_I),
    .O(MUX_SB_T0_SOUTH_SB_OUT_B17_O),
    .ready_in(SB_T0_SOUTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T0_SOUTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T0_SOUTH_SB_OUT_B17_valid_out),
    .S(SB_T0_SOUTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T0_WEST_SB_OUT_B17_I [6:0];
assign MUX_SB_T0_WEST_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T0_WEST_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T0_WEST_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T0_WEST_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T0_WEST_SB_OUT_B17_I[2] = WIRE_SB_T0_EAST_SB_IN_B17_O;
assign MUX_SB_T0_WEST_SB_OUT_B17_I[1] = WIRE_SB_T4_SOUTH_SB_IN_B17_O;
assign MUX_SB_T0_WEST_SB_OUT_B17_I[0] = WIRE_SB_T0_NORTH_SB_IN_B17_O;
wire [6:0] MUX_SB_T0_WEST_SB_OUT_B17_valid_in;
assign MUX_SB_T0_WEST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T0_EAST_SB_IN_B17_valid_out,WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T0_NORTH_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T0_WEST_SB_OUT_B17 (
    .I(MUX_SB_T0_WEST_SB_OUT_B17_I),
    .O(MUX_SB_T0_WEST_SB_OUT_B17_O),
    .ready_in(SB_T0_WEST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T0_WEST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T0_WEST_SB_OUT_B17_valid_out),
    .S(SB_T0_WEST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T0_WEST_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T1_EAST_SB_OUT_B17_I [6:0];
assign MUX_SB_T1_EAST_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T1_EAST_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T1_EAST_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T1_EAST_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T1_EAST_SB_OUT_B17_I[2] = WIRE_SB_T2_SOUTH_SB_IN_B17_O;
assign MUX_SB_T1_EAST_SB_OUT_B17_I[1] = WIRE_SB_T1_WEST_SB_IN_B17_O;
assign MUX_SB_T1_EAST_SB_OUT_B17_I[0] = WIRE_SB_T0_NORTH_SB_IN_B17_O;
wire [6:0] MUX_SB_T1_EAST_SB_OUT_B17_valid_in;
assign MUX_SB_T1_EAST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T1_WEST_SB_IN_B17_valid_out,WIRE_SB_T0_NORTH_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T1_EAST_SB_OUT_B17 (
    .I(MUX_SB_T1_EAST_SB_OUT_B17_I),
    .O(MUX_SB_T1_EAST_SB_OUT_B17_O),
    .ready_in(SB_T1_EAST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T1_EAST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T1_EAST_SB_OUT_B17_valid_out),
    .S(SB_T1_EAST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T1_EAST_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T1_NORTH_SB_OUT_B17_I [6:0];
assign MUX_SB_T1_NORTH_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T1_NORTH_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T1_NORTH_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T1_NORTH_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T1_NORTH_SB_OUT_B17_I[2] = WIRE_SB_T4_WEST_SB_IN_B17_O;
assign MUX_SB_T1_NORTH_SB_OUT_B17_I[1] = WIRE_SB_T1_SOUTH_SB_IN_B17_O;
assign MUX_SB_T1_NORTH_SB_OUT_B17_I[0] = WIRE_SB_T2_EAST_SB_IN_B17_O;
wire [6:0] MUX_SB_T1_NORTH_SB_OUT_B17_valid_in;
assign MUX_SB_T1_NORTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T4_WEST_SB_IN_B17_valid_out,WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T2_EAST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T1_NORTH_SB_OUT_B17 (
    .I(MUX_SB_T1_NORTH_SB_OUT_B17_I),
    .O(MUX_SB_T1_NORTH_SB_OUT_B17_O),
    .ready_in(SB_T1_NORTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T1_NORTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T1_NORTH_SB_OUT_B17_valid_out),
    .S(SB_T1_NORTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T1_SOUTH_SB_OUT_B17_I [6:0];
assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[2] = WIRE_SB_T2_WEST_SB_IN_B17_O;
assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[1] = WIRE_SB_T1_NORTH_SB_IN_B17_O;
assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[0] = WIRE_SB_T2_EAST_SB_IN_B17_O;
wire [6:0] MUX_SB_T1_SOUTH_SB_OUT_B17_valid_in;
assign MUX_SB_T1_SOUTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T2_WEST_SB_IN_B17_valid_out,WIRE_SB_T1_NORTH_SB_IN_B17_valid_out,WIRE_SB_T2_EAST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T1_SOUTH_SB_OUT_B17 (
    .I(MUX_SB_T1_SOUTH_SB_OUT_B17_I),
    .O(MUX_SB_T1_SOUTH_SB_OUT_B17_O),
    .ready_in(SB_T1_SOUTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T1_SOUTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T1_SOUTH_SB_OUT_B17_valid_out),
    .S(SB_T1_SOUTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T1_WEST_SB_OUT_B17_I [6:0];
assign MUX_SB_T1_WEST_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T1_WEST_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T1_WEST_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T1_WEST_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T1_WEST_SB_OUT_B17_I[2] = WIRE_SB_T1_EAST_SB_IN_B17_O;
assign MUX_SB_T1_WEST_SB_OUT_B17_I[1] = WIRE_SB_T0_SOUTH_SB_IN_B17_O;
assign MUX_SB_T1_WEST_SB_OUT_B17_I[0] = WIRE_SB_T4_NORTH_SB_IN_B17_O;
wire [6:0] MUX_SB_T1_WEST_SB_OUT_B17_valid_in;
assign MUX_SB_T1_WEST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T1_EAST_SB_IN_B17_valid_out,WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T4_NORTH_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T1_WEST_SB_OUT_B17 (
    .I(MUX_SB_T1_WEST_SB_OUT_B17_I),
    .O(MUX_SB_T1_WEST_SB_OUT_B17_O),
    .ready_in(SB_T1_WEST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T1_WEST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T1_WEST_SB_OUT_B17_valid_out),
    .S(SB_T1_WEST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T1_WEST_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T2_EAST_SB_OUT_B17_I [6:0];
assign MUX_SB_T2_EAST_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T2_EAST_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T2_EAST_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T2_EAST_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T2_EAST_SB_OUT_B17_I[2] = WIRE_SB_T2_WEST_SB_IN_B17_O;
assign MUX_SB_T2_EAST_SB_OUT_B17_I[1] = WIRE_SB_T1_SOUTH_SB_IN_B17_O;
assign MUX_SB_T2_EAST_SB_OUT_B17_I[0] = WIRE_SB_T1_NORTH_SB_IN_B17_O;
wire [6:0] MUX_SB_T2_EAST_SB_OUT_B17_valid_in;
assign MUX_SB_T2_EAST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T2_WEST_SB_IN_B17_valid_out,WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T1_NORTH_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T2_EAST_SB_OUT_B17 (
    .I(MUX_SB_T2_EAST_SB_OUT_B17_I),
    .O(MUX_SB_T2_EAST_SB_OUT_B17_O),
    .ready_in(SB_T2_EAST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T2_EAST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T2_EAST_SB_OUT_B17_valid_out),
    .S(SB_T2_EAST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T2_EAST_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T2_NORTH_SB_OUT_B17_I [6:0];
assign MUX_SB_T2_NORTH_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T2_NORTH_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T2_NORTH_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T2_NORTH_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T2_NORTH_SB_OUT_B17_I[2] = WIRE_SB_T3_WEST_SB_IN_B17_O;
assign MUX_SB_T2_NORTH_SB_OUT_B17_I[1] = WIRE_SB_T2_SOUTH_SB_IN_B17_O;
assign MUX_SB_T2_NORTH_SB_OUT_B17_I[0] = WIRE_SB_T3_EAST_SB_IN_B17_O;
wire [6:0] MUX_SB_T2_NORTH_SB_OUT_B17_valid_in;
assign MUX_SB_T2_NORTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T3_WEST_SB_IN_B17_valid_out,WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T3_EAST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T2_NORTH_SB_OUT_B17 (
    .I(MUX_SB_T2_NORTH_SB_OUT_B17_I),
    .O(MUX_SB_T2_NORTH_SB_OUT_B17_O),
    .ready_in(SB_T2_NORTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T2_NORTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T2_NORTH_SB_OUT_B17_valid_out),
    .S(SB_T2_NORTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T2_SOUTH_SB_OUT_B17_I [6:0];
assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[2] = WIRE_SB_T3_WEST_SB_IN_B17_O;
assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[1] = WIRE_SB_T2_NORTH_SB_IN_B17_O;
assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[0] = WIRE_SB_T1_EAST_SB_IN_B17_O;
wire [6:0] MUX_SB_T2_SOUTH_SB_OUT_B17_valid_in;
assign MUX_SB_T2_SOUTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T3_WEST_SB_IN_B17_valid_out,WIRE_SB_T2_NORTH_SB_IN_B17_valid_out,WIRE_SB_T1_EAST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T2_SOUTH_SB_OUT_B17 (
    .I(MUX_SB_T2_SOUTH_SB_OUT_B17_I),
    .O(MUX_SB_T2_SOUTH_SB_OUT_B17_O),
    .ready_in(SB_T2_SOUTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T2_SOUTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T2_SOUTH_SB_OUT_B17_valid_out),
    .S(SB_T2_SOUTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T2_WEST_SB_OUT_B17_I [6:0];
assign MUX_SB_T2_WEST_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T2_WEST_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T2_WEST_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T2_WEST_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T2_WEST_SB_OUT_B17_I[2] = WIRE_SB_T2_EAST_SB_IN_B17_O;
assign MUX_SB_T2_WEST_SB_OUT_B17_I[1] = WIRE_SB_T1_SOUTH_SB_IN_B17_O;
assign MUX_SB_T2_WEST_SB_OUT_B17_I[0] = WIRE_SB_T3_NORTH_SB_IN_B17_O;
wire [6:0] MUX_SB_T2_WEST_SB_OUT_B17_valid_in;
assign MUX_SB_T2_WEST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T2_EAST_SB_IN_B17_valid_out,WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T3_NORTH_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T2_WEST_SB_OUT_B17 (
    .I(MUX_SB_T2_WEST_SB_OUT_B17_I),
    .O(MUX_SB_T2_WEST_SB_OUT_B17_O),
    .ready_in(SB_T2_WEST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T2_WEST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T2_WEST_SB_OUT_B17_valid_out),
    .S(SB_T2_WEST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T2_WEST_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T3_EAST_SB_OUT_B17_I [6:0];
assign MUX_SB_T3_EAST_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T3_EAST_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T3_EAST_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T3_EAST_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T3_EAST_SB_OUT_B17_I[2] = WIRE_SB_T3_WEST_SB_IN_B17_O;
assign MUX_SB_T3_EAST_SB_OUT_B17_I[1] = WIRE_SB_T2_NORTH_SB_IN_B17_O;
assign MUX_SB_T3_EAST_SB_OUT_B17_I[0] = WIRE_SB_T0_SOUTH_SB_IN_B17_O;
wire [6:0] MUX_SB_T3_EAST_SB_OUT_B17_valid_in;
assign MUX_SB_T3_EAST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T3_WEST_SB_IN_B17_valid_out,WIRE_SB_T2_NORTH_SB_IN_B17_valid_out,WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T3_EAST_SB_OUT_B17 (
    .I(MUX_SB_T3_EAST_SB_OUT_B17_I),
    .O(MUX_SB_T3_EAST_SB_OUT_B17_O),
    .ready_in(SB_T3_EAST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T3_EAST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T3_EAST_SB_OUT_B17_valid_out),
    .S(SB_T3_EAST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T3_EAST_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T3_NORTH_SB_OUT_B17_I [6:0];
assign MUX_SB_T3_NORTH_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T3_NORTH_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T3_NORTH_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T3_NORTH_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T3_NORTH_SB_OUT_B17_I[2] = WIRE_SB_T3_SOUTH_SB_IN_B17_O;
assign MUX_SB_T3_NORTH_SB_OUT_B17_I[1] = WIRE_SB_T4_EAST_SB_IN_B17_O;
assign MUX_SB_T3_NORTH_SB_OUT_B17_I[0] = WIRE_SB_T2_WEST_SB_IN_B17_O;
wire [6:0] MUX_SB_T3_NORTH_SB_OUT_B17_valid_in;
assign MUX_SB_T3_NORTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T4_EAST_SB_IN_B17_valid_out,WIRE_SB_T2_WEST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T3_NORTH_SB_OUT_B17 (
    .I(MUX_SB_T3_NORTH_SB_OUT_B17_I),
    .O(MUX_SB_T3_NORTH_SB_OUT_B17_O),
    .ready_in(SB_T3_NORTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T3_NORTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T3_NORTH_SB_OUT_B17_valid_out),
    .S(SB_T3_NORTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T3_SOUTH_SB_OUT_B17_I [6:0];
assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[2] = WIRE_SB_T4_WEST_SB_IN_B17_O;
assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[1] = WIRE_SB_T3_NORTH_SB_IN_B17_O;
assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[0] = WIRE_SB_T0_EAST_SB_IN_B17_O;
wire [6:0] MUX_SB_T3_SOUTH_SB_OUT_B17_valid_in;
assign MUX_SB_T3_SOUTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T4_WEST_SB_IN_B17_valid_out,WIRE_SB_T3_NORTH_SB_IN_B17_valid_out,WIRE_SB_T0_EAST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T3_SOUTH_SB_OUT_B17 (
    .I(MUX_SB_T3_SOUTH_SB_OUT_B17_I),
    .O(MUX_SB_T3_SOUTH_SB_OUT_B17_O),
    .ready_in(SB_T3_SOUTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T3_SOUTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T3_SOUTH_SB_OUT_B17_valid_out),
    .S(SB_T3_SOUTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T3_WEST_SB_OUT_B17_I [6:0];
assign MUX_SB_T3_WEST_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T3_WEST_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T3_WEST_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T3_WEST_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T3_WEST_SB_OUT_B17_I[2] = WIRE_SB_T3_EAST_SB_IN_B17_O;
assign MUX_SB_T3_WEST_SB_OUT_B17_I[1] = WIRE_SB_T2_SOUTH_SB_IN_B17_O;
assign MUX_SB_T3_WEST_SB_OUT_B17_I[0] = WIRE_SB_T2_NORTH_SB_IN_B17_O;
wire [6:0] MUX_SB_T3_WEST_SB_OUT_B17_valid_in;
assign MUX_SB_T3_WEST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T3_EAST_SB_IN_B17_valid_out,WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T2_NORTH_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T3_WEST_SB_OUT_B17 (
    .I(MUX_SB_T3_WEST_SB_OUT_B17_I),
    .O(MUX_SB_T3_WEST_SB_OUT_B17_O),
    .ready_in(SB_T3_WEST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T3_WEST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T3_WEST_SB_OUT_B17_valid_out),
    .S(SB_T3_WEST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T3_WEST_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T4_EAST_SB_OUT_B17_I [6:0];
assign MUX_SB_T4_EAST_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T4_EAST_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T4_EAST_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T4_EAST_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T4_EAST_SB_OUT_B17_I[2] = WIRE_SB_T4_WEST_SB_IN_B17_O;
assign MUX_SB_T4_EAST_SB_OUT_B17_I[1] = WIRE_SB_T4_SOUTH_SB_IN_B17_O;
assign MUX_SB_T4_EAST_SB_OUT_B17_I[0] = WIRE_SB_T3_NORTH_SB_IN_B17_O;
wire [6:0] MUX_SB_T4_EAST_SB_OUT_B17_valid_in;
assign MUX_SB_T4_EAST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T4_WEST_SB_IN_B17_valid_out,WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T3_NORTH_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T4_EAST_SB_OUT_B17 (
    .I(MUX_SB_T4_EAST_SB_OUT_B17_I),
    .O(MUX_SB_T4_EAST_SB_OUT_B17_O),
    .ready_in(SB_T4_EAST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T4_EAST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T4_EAST_SB_OUT_B17_valid_out),
    .S(SB_T4_EAST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T4_EAST_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T4_NORTH_SB_OUT_B17_I [6:0];
assign MUX_SB_T4_NORTH_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T4_NORTH_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T4_NORTH_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T4_NORTH_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T4_NORTH_SB_OUT_B17_I[2] = WIRE_SB_T4_SOUTH_SB_IN_B17_O;
assign MUX_SB_T4_NORTH_SB_OUT_B17_I[1] = WIRE_SB_T0_EAST_SB_IN_B17_O;
assign MUX_SB_T4_NORTH_SB_OUT_B17_I[0] = WIRE_SB_T1_WEST_SB_IN_B17_O;
wire [6:0] MUX_SB_T4_NORTH_SB_OUT_B17_valid_in;
assign MUX_SB_T4_NORTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T0_EAST_SB_IN_B17_valid_out,WIRE_SB_T1_WEST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T4_NORTH_SB_OUT_B17 (
    .I(MUX_SB_T4_NORTH_SB_OUT_B17_I),
    .O(MUX_SB_T4_NORTH_SB_OUT_B17_O),
    .ready_in(SB_T4_NORTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T4_NORTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T4_NORTH_SB_OUT_B17_valid_out),
    .S(SB_T4_NORTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T4_SOUTH_SB_OUT_B17_I [6:0];
assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[2] = WIRE_SB_T4_NORTH_SB_IN_B17_O;
assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[1] = WIRE_SB_T4_EAST_SB_IN_B17_O;
assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[0] = WIRE_SB_T0_WEST_SB_IN_B17_O;
wire [6:0] MUX_SB_T4_SOUTH_SB_OUT_B17_valid_in;
assign MUX_SB_T4_SOUTH_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T4_NORTH_SB_IN_B17_valid_out,WIRE_SB_T4_EAST_SB_IN_B17_valid_out,WIRE_SB_T0_WEST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T4_SOUTH_SB_OUT_B17 (
    .I(MUX_SB_T4_SOUTH_SB_OUT_B17_I),
    .O(MUX_SB_T4_SOUTH_SB_OUT_B17_O),
    .ready_in(SB_T4_SOUTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T4_SOUTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T4_SOUTH_SB_OUT_B17_valid_out),
    .S(SB_T4_SOUTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T4_WEST_SB_OUT_B17_I [6:0];
assign MUX_SB_T4_WEST_SB_OUT_B17_I[6] = PondTop_output_width_17_num_1;
assign MUX_SB_T4_WEST_SB_OUT_B17_I[5] = PE_output_width_17_num_2;
assign MUX_SB_T4_WEST_SB_OUT_B17_I[4] = PE_output_width_17_num_1;
assign MUX_SB_T4_WEST_SB_OUT_B17_I[3] = PE_output_width_17_num_0;
assign MUX_SB_T4_WEST_SB_OUT_B17_I[2] = WIRE_SB_T4_EAST_SB_IN_B17_O;
assign MUX_SB_T4_WEST_SB_OUT_B17_I[1] = WIRE_SB_T3_SOUTH_SB_IN_B17_O;
assign MUX_SB_T4_WEST_SB_OUT_B17_I[0] = WIRE_SB_T1_NORTH_SB_IN_B17_O;
wire [6:0] MUX_SB_T4_WEST_SB_OUT_B17_valid_in;
assign MUX_SB_T4_WEST_SB_OUT_B17_valid_in = {PondTop_output_width_17_num_1_valid,PE_output_width_17_num_2_valid,PE_output_width_17_num_1_valid,PE_output_width_17_num_0_valid,WIRE_SB_T4_EAST_SB_IN_B17_valid_out,WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T1_NORTH_SB_IN_B17_valid_out};
mux_aoi_ready_valid_7_17 MUX_SB_T4_WEST_SB_OUT_B17 (
    .I(MUX_SB_T4_WEST_SB_OUT_B17_I),
    .O(MUX_SB_T4_WEST_SB_OUT_B17_O),
    .ready_in(SB_T4_WEST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T4_WEST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T4_WEST_SB_OUT_B17_valid_out),
    .S(SB_T4_WEST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T4_WEST_SB_OUT_B17_out_sel)
);
SplitFifo_17 REG_T0_EAST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T0_EAST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T0_EAST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T0_EAST_B17_fifo_value_O[0]),
    .end_fifo(REG_T0_EAST_B17_end_value_O[0]),
    .data_in(MUX_SB_T0_EAST_SB_OUT_B17_O),
    .ready1(RMUX_T0_EAST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T0_EAST_SB_OUT_B17_valid_out),
    .data_out(REG_T0_EAST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T0_EAST_B17_start_value_O[0]),
    .clk_en(and1_inst2_out[0])
);
SliceWrapper_32_0_1 REG_T0_EAST_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T0_EAST_B17_end_value_O)
);
SliceWrapper_32_1_2 REG_T0_EAST_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T0_EAST_B17_fifo_value_O)
);
SliceWrapper_32_2_3 REG_T0_EAST_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T0_EAST_B17_start_value_O)
);
SplitFifo_17 REG_T0_NORTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T0_NORTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T0_NORTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T0_NORTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T0_NORTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T0_NORTH_SB_OUT_B17_O),
    .ready1(RMUX_T0_NORTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T0_NORTH_SB_OUT_B17_valid_out),
    .data_out(REG_T0_NORTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T0_NORTH_B17_start_value_O[0]),
    .clk_en(and1_inst0_out[0])
);
SliceWrapper_32_3_4 REG_T0_NORTH_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T0_NORTH_B17_end_value_O)
);
SliceWrapper_32_4_5 REG_T0_NORTH_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T0_NORTH_B17_fifo_value_O)
);
SliceWrapper_32_5_6 REG_T0_NORTH_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T0_NORTH_B17_start_value_O)
);
SplitFifo_17 REG_T0_SOUTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T0_SOUTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T0_SOUTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T0_SOUTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T0_SOUTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T0_SOUTH_SB_OUT_B17_O),
    .ready1(RMUX_T0_SOUTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T0_SOUTH_SB_OUT_B17_valid_out),
    .data_out(REG_T0_SOUTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T0_SOUTH_B17_start_value_O[0]),
    .clk_en(and1_inst1_out[0])
);
SliceWrapper_32_6_7 REG_T0_SOUTH_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T0_SOUTH_B17_end_value_O)
);
SliceWrapper_32_7_8 REG_T0_SOUTH_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T0_SOUTH_B17_fifo_value_O)
);
SliceWrapper_32_8_9 REG_T0_SOUTH_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T0_SOUTH_B17_start_value_O)
);
SplitFifo_17 REG_T0_WEST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T0_WEST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T0_WEST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T0_WEST_B17_fifo_value_O[0]),
    .end_fifo(REG_T0_WEST_B17_end_value_O[0]),
    .data_in(MUX_SB_T0_WEST_SB_OUT_B17_O),
    .ready1(RMUX_T0_WEST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T0_WEST_SB_OUT_B17_valid_out),
    .data_out(REG_T0_WEST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T0_WEST_B17_start_value_O[0]),
    .clk_en(and1_inst3_out[0])
);
SliceWrapper_32_9_10 REG_T0_WEST_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T0_WEST_B17_end_value_O)
);
SliceWrapper_32_10_11 REG_T0_WEST_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T0_WEST_B17_fifo_value_O)
);
SliceWrapper_32_11_12 REG_T0_WEST_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T0_WEST_B17_start_value_O)
);
SplitFifo_17 REG_T1_EAST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T1_EAST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T1_EAST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T1_EAST_B17_fifo_value_O[0]),
    .end_fifo(REG_T1_EAST_B17_end_value_O[0]),
    .data_in(MUX_SB_T1_EAST_SB_OUT_B17_O),
    .ready1(RMUX_T1_EAST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T1_EAST_SB_OUT_B17_valid_out),
    .data_out(REG_T1_EAST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T1_EAST_B17_start_value_O[0]),
    .clk_en(and1_inst6_out[0])
);
SliceWrapper_32_12_13 REG_T1_EAST_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T1_EAST_B17_end_value_O)
);
SliceWrapper_32_13_14 REG_T1_EAST_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T1_EAST_B17_fifo_value_O)
);
SliceWrapper_32_14_15 REG_T1_EAST_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T1_EAST_B17_start_value_O)
);
SplitFifo_17 REG_T1_NORTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T1_NORTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T1_NORTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T1_NORTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T1_NORTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T1_NORTH_SB_OUT_B17_O),
    .ready1(RMUX_T1_NORTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T1_NORTH_SB_OUT_B17_valid_out),
    .data_out(REG_T1_NORTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T1_NORTH_B17_start_value_O[0]),
    .clk_en(and1_inst4_out[0])
);
SliceWrapper_32_15_16 REG_T1_NORTH_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T1_NORTH_B17_end_value_O)
);
SliceWrapper_32_16_17 REG_T1_NORTH_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T1_NORTH_B17_fifo_value_O)
);
SliceWrapper_32_17_18 REG_T1_NORTH_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T1_NORTH_B17_start_value_O)
);
SplitFifo_17 REG_T1_SOUTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T1_SOUTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T1_SOUTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T1_SOUTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T1_SOUTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T1_SOUTH_SB_OUT_B17_O),
    .ready1(RMUX_T1_SOUTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T1_SOUTH_SB_OUT_B17_valid_out),
    .data_out(REG_T1_SOUTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T1_SOUTH_B17_start_value_O[0]),
    .clk_en(and1_inst5_out[0])
);
SliceWrapper_32_18_19 REG_T1_SOUTH_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T1_SOUTH_B17_end_value_O)
);
SliceWrapper_32_19_20 REG_T1_SOUTH_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T1_SOUTH_B17_fifo_value_O)
);
SliceWrapper_32_20_21 REG_T1_SOUTH_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T1_SOUTH_B17_start_value_O)
);
SplitFifo_17 REG_T1_WEST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T1_WEST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T1_WEST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T1_WEST_B17_fifo_value_O[0]),
    .end_fifo(REG_T1_WEST_B17_end_value_O[0]),
    .data_in(MUX_SB_T1_WEST_SB_OUT_B17_O),
    .ready1(RMUX_T1_WEST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T1_WEST_SB_OUT_B17_valid_out),
    .data_out(REG_T1_WEST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T1_WEST_B17_start_value_O[0]),
    .clk_en(and1_inst7_out[0])
);
SliceWrapper_32_21_22 REG_T1_WEST_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T1_WEST_B17_end_value_O)
);
SliceWrapper_32_22_23 REG_T1_WEST_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T1_WEST_B17_fifo_value_O)
);
SliceWrapper_32_23_24 REG_T1_WEST_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T1_WEST_B17_start_value_O)
);
SplitFifo_17 REG_T2_EAST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T2_EAST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T2_EAST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T2_EAST_B17_fifo_value_O[0]),
    .end_fifo(REG_T2_EAST_B17_end_value_O[0]),
    .data_in(MUX_SB_T2_EAST_SB_OUT_B17_O),
    .ready1(RMUX_T2_EAST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T2_EAST_SB_OUT_B17_valid_out),
    .data_out(REG_T2_EAST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T2_EAST_B17_start_value_O[0]),
    .clk_en(and1_inst10_out[0])
);
SliceWrapper_32_24_25 REG_T2_EAST_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T2_EAST_B17_end_value_O)
);
SliceWrapper_32_25_26 REG_T2_EAST_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T2_EAST_B17_fifo_value_O)
);
SliceWrapper_32_26_27 REG_T2_EAST_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T2_EAST_B17_start_value_O)
);
SplitFifo_17 REG_T2_NORTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T2_NORTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T2_NORTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T2_NORTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T2_NORTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T2_NORTH_SB_OUT_B17_O),
    .ready1(RMUX_T2_NORTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T2_NORTH_SB_OUT_B17_valid_out),
    .data_out(REG_T2_NORTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T2_NORTH_B17_start_value_O[0]),
    .clk_en(and1_inst8_out[0])
);
SliceWrapper_32_27_28 REG_T2_NORTH_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T2_NORTH_B17_end_value_O)
);
SliceWrapper_32_28_29 REG_T2_NORTH_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T2_NORTH_B17_fifo_value_O)
);
SliceWrapper_32_29_30 REG_T2_NORTH_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T2_NORTH_B17_start_value_O)
);
SplitFifo_17 REG_T2_SOUTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T2_SOUTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T2_SOUTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T2_SOUTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T2_SOUTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T2_SOUTH_SB_OUT_B17_O),
    .ready1(RMUX_T2_SOUTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T2_SOUTH_SB_OUT_B17_valid_out),
    .data_out(REG_T2_SOUTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T2_SOUTH_B17_start_value_O[0]),
    .clk_en(and1_inst9_out[0])
);
SliceWrapper_32_30_31 REG_T2_SOUTH_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T2_SOUTH_B17_end_value_O)
);
SliceWrapper_32_31_32 REG_T2_SOUTH_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T2_SOUTH_B17_fifo_value_O)
);
SliceWrapper_32_0_1 REG_T2_SOUTH_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T2_SOUTH_B17_start_value_O)
);
SplitFifo_17 REG_T2_WEST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T2_WEST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T2_WEST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T2_WEST_B17_fifo_value_O[0]),
    .end_fifo(REG_T2_WEST_B17_end_value_O[0]),
    .data_in(MUX_SB_T2_WEST_SB_OUT_B17_O),
    .ready1(RMUX_T2_WEST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T2_WEST_SB_OUT_B17_valid_out),
    .data_out(REG_T2_WEST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T2_WEST_B17_start_value_O[0]),
    .clk_en(and1_inst11_out[0])
);
SliceWrapper_32_1_2 REG_T2_WEST_B17_end_value (
    .I(config_reg_1_O),
    .O(REG_T2_WEST_B17_end_value_O)
);
SliceWrapper_32_2_3 REG_T2_WEST_B17_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T2_WEST_B17_fifo_value_O)
);
SliceWrapper_32_3_4 REG_T2_WEST_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T2_WEST_B17_start_value_O)
);
SplitFifo_17 REG_T3_EAST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T3_EAST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T3_EAST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T3_EAST_B17_fifo_value_O[0]),
    .end_fifo(REG_T3_EAST_B17_end_value_O[0]),
    .data_in(MUX_SB_T3_EAST_SB_OUT_B17_O),
    .ready1(RMUX_T3_EAST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T3_EAST_SB_OUT_B17_valid_out),
    .data_out(REG_T3_EAST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T3_EAST_B17_start_value_O[0]),
    .clk_en(and1_inst14_out[0])
);
SliceWrapper_32_4_5 REG_T3_EAST_B17_end_value (
    .I(config_reg_1_O),
    .O(REG_T3_EAST_B17_end_value_O)
);
SliceWrapper_32_5_6 REG_T3_EAST_B17_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T3_EAST_B17_fifo_value_O)
);
SliceWrapper_32_6_7 REG_T3_EAST_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T3_EAST_B17_start_value_O)
);
SplitFifo_17 REG_T3_NORTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T3_NORTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T3_NORTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T3_NORTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T3_NORTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T3_NORTH_SB_OUT_B17_O),
    .ready1(RMUX_T3_NORTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T3_NORTH_SB_OUT_B17_valid_out),
    .data_out(REG_T3_NORTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T3_NORTH_B17_start_value_O[0]),
    .clk_en(and1_inst12_out[0])
);
SliceWrapper_32_7_8 REG_T3_NORTH_B17_end_value (
    .I(config_reg_1_O),
    .O(REG_T3_NORTH_B17_end_value_O)
);
SliceWrapper_32_8_9 REG_T3_NORTH_B17_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T3_NORTH_B17_fifo_value_O)
);
SliceWrapper_32_9_10 REG_T3_NORTH_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T3_NORTH_B17_start_value_O)
);
SplitFifo_17 REG_T3_SOUTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T3_SOUTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T3_SOUTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T3_SOUTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T3_SOUTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T3_SOUTH_SB_OUT_B17_O),
    .ready1(RMUX_T3_SOUTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T3_SOUTH_SB_OUT_B17_valid_out),
    .data_out(REG_T3_SOUTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T3_SOUTH_B17_start_value_O[0]),
    .clk_en(and1_inst13_out[0])
);
SliceWrapper_32_10_11 REG_T3_SOUTH_B17_end_value (
    .I(config_reg_1_O),
    .O(REG_T3_SOUTH_B17_end_value_O)
);
SliceWrapper_32_11_12 REG_T3_SOUTH_B17_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T3_SOUTH_B17_fifo_value_O)
);
SliceWrapper_32_12_13 REG_T3_SOUTH_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T3_SOUTH_B17_start_value_O)
);
SplitFifo_17 REG_T3_WEST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T3_WEST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T3_WEST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T3_WEST_B17_fifo_value_O[0]),
    .end_fifo(REG_T3_WEST_B17_end_value_O[0]),
    .data_in(MUX_SB_T3_WEST_SB_OUT_B17_O),
    .ready1(RMUX_T3_WEST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T3_WEST_SB_OUT_B17_valid_out),
    .data_out(REG_T3_WEST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T3_WEST_B17_start_value_O[0]),
    .clk_en(and1_inst15_out[0])
);
SliceWrapper_32_13_14 REG_T3_WEST_B17_end_value (
    .I(config_reg_1_O),
    .O(REG_T3_WEST_B17_end_value_O)
);
SliceWrapper_32_14_15 REG_T3_WEST_B17_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T3_WEST_B17_fifo_value_O)
);
SliceWrapper_32_15_16 REG_T3_WEST_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T3_WEST_B17_start_value_O)
);
SplitFifo_17 REG_T4_EAST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T4_EAST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T4_EAST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T4_EAST_B17_fifo_value_O[0]),
    .end_fifo(REG_T4_EAST_B17_end_value_O[0]),
    .data_in(MUX_SB_T4_EAST_SB_OUT_B17_O),
    .ready1(RMUX_T4_EAST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T4_EAST_SB_OUT_B17_valid_out),
    .data_out(REG_T4_EAST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T4_EAST_B17_start_value_O[0]),
    .clk_en(and1_inst18_out[0])
);
SliceWrapper_32_16_17 REG_T4_EAST_B17_end_value (
    .I(config_reg_1_O),
    .O(REG_T4_EAST_B17_end_value_O)
);
SliceWrapper_32_17_18 REG_T4_EAST_B17_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T4_EAST_B17_fifo_value_O)
);
SliceWrapper_32_18_19 REG_T4_EAST_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T4_EAST_B17_start_value_O)
);
SplitFifo_17 REG_T4_NORTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T4_NORTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T4_NORTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T4_NORTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T4_NORTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T4_NORTH_SB_OUT_B17_O),
    .ready1(RMUX_T4_NORTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T4_NORTH_SB_OUT_B17_valid_out),
    .data_out(REG_T4_NORTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T4_NORTH_B17_start_value_O[0]),
    .clk_en(and1_inst16_out[0])
);
SliceWrapper_32_19_20 REG_T4_NORTH_B17_end_value (
    .I(config_reg_1_O),
    .O(REG_T4_NORTH_B17_end_value_O)
);
SliceWrapper_32_20_21 REG_T4_NORTH_B17_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T4_NORTH_B17_fifo_value_O)
);
SliceWrapper_32_21_22 REG_T4_NORTH_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T4_NORTH_B17_start_value_O)
);
SplitFifo_17 REG_T4_SOUTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T4_SOUTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T4_SOUTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T4_SOUTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T4_SOUTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T4_SOUTH_SB_OUT_B17_O),
    .ready1(RMUX_T4_SOUTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T4_SOUTH_SB_OUT_B17_valid_out),
    .data_out(REG_T4_SOUTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T4_SOUTH_B17_start_value_O[0]),
    .clk_en(and1_inst17_out[0])
);
SliceWrapper_32_22_23 REG_T4_SOUTH_B17_end_value (
    .I(config_reg_1_O),
    .O(REG_T4_SOUTH_B17_end_value_O)
);
SliceWrapper_32_23_24 REG_T4_SOUTH_B17_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T4_SOUTH_B17_fifo_value_O)
);
SliceWrapper_32_24_25 REG_T4_SOUTH_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T4_SOUTH_B17_start_value_O)
);
SplitFifo_17 REG_T4_WEST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T4_WEST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T4_WEST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T4_WEST_B17_fifo_value_O[0]),
    .end_fifo(REG_T4_WEST_B17_end_value_O[0]),
    .data_in(MUX_SB_T4_WEST_SB_OUT_B17_O),
    .ready1(RMUX_T4_WEST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T4_WEST_SB_OUT_B17_valid_out),
    .data_out(REG_T4_WEST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T4_WEST_B17_start_value_O[0]),
    .clk_en(and1_inst19_out[0])
);
SliceWrapper_32_25_26 REG_T4_WEST_B17_end_value (
    .I(config_reg_1_O),
    .O(REG_T4_WEST_B17_end_value_O)
);
SliceWrapper_32_26_27 REG_T4_WEST_B17_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T4_WEST_B17_fifo_value_O)
);
SliceWrapper_32_27_28 REG_T4_WEST_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T4_WEST_B17_start_value_O)
);
wire [16:0] RMUX_T0_EAST_B17_I [1:0];
assign RMUX_T0_EAST_B17_I[1] = REG_T0_EAST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T0_EAST_B17_I[0] = MUX_SB_T0_EAST_SB_OUT_B17_O;
wire [1:0] RMUX_T0_EAST_B17_valid_in;
assign RMUX_T0_EAST_B17_valid_in = {REG_T0_EAST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T0_EAST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T0_EAST_B17 (
    .I(RMUX_T0_EAST_B17_I),
    .O(RMUX_T0_EAST_B17_O),
    .ready_in(SB_T0_EAST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T0_EAST_B17_ready_out),
    .valid_in(RMUX_T0_EAST_B17_valid_in),
    .valid_out(RMUX_T0_EAST_B17_valid_out),
    .S(RMUX_T0_EAST_B17_sel_value_O),
    .out_sel(RMUX_T0_EAST_B17_out_sel)
);
SliceWrapper_32_28_29 RMUX_T0_EAST_B17_sel_value (
    .I(config_reg_1_O),
    .O(RMUX_T0_EAST_B17_sel_value_O)
);
wire [16:0] RMUX_T0_NORTH_B17_I [1:0];
assign RMUX_T0_NORTH_B17_I[1] = REG_T0_NORTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T0_NORTH_B17_I[0] = MUX_SB_T0_NORTH_SB_OUT_B17_O;
wire [1:0] RMUX_T0_NORTH_B17_valid_in;
assign RMUX_T0_NORTH_B17_valid_in = {REG_T0_NORTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T0_NORTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T0_NORTH_B17 (
    .I(RMUX_T0_NORTH_B17_I),
    .O(RMUX_T0_NORTH_B17_O),
    .ready_in(SB_T0_NORTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T0_NORTH_B17_ready_out),
    .valid_in(RMUX_T0_NORTH_B17_valid_in),
    .valid_out(RMUX_T0_NORTH_B17_valid_out),
    .S(RMUX_T0_NORTH_B17_sel_value_O),
    .out_sel(RMUX_T0_NORTH_B17_out_sel)
);
SliceWrapper_32_29_30 RMUX_T0_NORTH_B17_sel_value (
    .I(config_reg_1_O),
    .O(RMUX_T0_NORTH_B17_sel_value_O)
);
wire [16:0] RMUX_T0_SOUTH_B17_I [1:0];
assign RMUX_T0_SOUTH_B17_I[1] = REG_T0_SOUTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T0_SOUTH_B17_I[0] = MUX_SB_T0_SOUTH_SB_OUT_B17_O;
wire [1:0] RMUX_T0_SOUTH_B17_valid_in;
assign RMUX_T0_SOUTH_B17_valid_in = {REG_T0_SOUTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T0_SOUTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T0_SOUTH_B17 (
    .I(RMUX_T0_SOUTH_B17_I),
    .O(RMUX_T0_SOUTH_B17_O),
    .ready_in(SB_T0_SOUTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T0_SOUTH_B17_ready_out),
    .valid_in(RMUX_T0_SOUTH_B17_valid_in),
    .valid_out(RMUX_T0_SOUTH_B17_valid_out),
    .S(RMUX_T0_SOUTH_B17_sel_value_O),
    .out_sel(RMUX_T0_SOUTH_B17_out_sel)
);
SliceWrapper_32_30_31 RMUX_T0_SOUTH_B17_sel_value (
    .I(config_reg_1_O),
    .O(RMUX_T0_SOUTH_B17_sel_value_O)
);
wire [16:0] RMUX_T0_WEST_B17_I [1:0];
assign RMUX_T0_WEST_B17_I[1] = REG_T0_WEST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T0_WEST_B17_I[0] = MUX_SB_T0_WEST_SB_OUT_B17_O;
wire [1:0] RMUX_T0_WEST_B17_valid_in;
assign RMUX_T0_WEST_B17_valid_in = {REG_T0_WEST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T0_WEST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T0_WEST_B17 (
    .I(RMUX_T0_WEST_B17_I),
    .O(RMUX_T0_WEST_B17_O),
    .ready_in(SB_T0_WEST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T0_WEST_B17_ready_out),
    .valid_in(RMUX_T0_WEST_B17_valid_in),
    .valid_out(RMUX_T0_WEST_B17_valid_out),
    .S(RMUX_T0_WEST_B17_sel_value_O),
    .out_sel(RMUX_T0_WEST_B17_out_sel)
);
SliceWrapper_32_31_32 RMUX_T0_WEST_B17_sel_value (
    .I(config_reg_1_O),
    .O(RMUX_T0_WEST_B17_sel_value_O)
);
wire [16:0] RMUX_T1_EAST_B17_I [1:0];
assign RMUX_T1_EAST_B17_I[1] = REG_T1_EAST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T1_EAST_B17_I[0] = MUX_SB_T1_EAST_SB_OUT_B17_O;
wire [1:0] RMUX_T1_EAST_B17_valid_in;
assign RMUX_T1_EAST_B17_valid_in = {REG_T1_EAST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T1_EAST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T1_EAST_B17 (
    .I(RMUX_T1_EAST_B17_I),
    .O(RMUX_T1_EAST_B17_O),
    .ready_in(SB_T1_EAST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T1_EAST_B17_ready_out),
    .valid_in(RMUX_T1_EAST_B17_valid_in),
    .valid_out(RMUX_T1_EAST_B17_valid_out),
    .S(RMUX_T1_EAST_B17_sel_value_O),
    .out_sel(RMUX_T1_EAST_B17_out_sel)
);
SliceWrapper_32_0_1 RMUX_T1_EAST_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T1_EAST_B17_sel_value_O)
);
wire [16:0] RMUX_T1_NORTH_B17_I [1:0];
assign RMUX_T1_NORTH_B17_I[1] = REG_T1_NORTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T1_NORTH_B17_I[0] = MUX_SB_T1_NORTH_SB_OUT_B17_O;
wire [1:0] RMUX_T1_NORTH_B17_valid_in;
assign RMUX_T1_NORTH_B17_valid_in = {REG_T1_NORTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T1_NORTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T1_NORTH_B17 (
    .I(RMUX_T1_NORTH_B17_I),
    .O(RMUX_T1_NORTH_B17_O),
    .ready_in(SB_T1_NORTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T1_NORTH_B17_ready_out),
    .valid_in(RMUX_T1_NORTH_B17_valid_in),
    .valid_out(RMUX_T1_NORTH_B17_valid_out),
    .S(RMUX_T1_NORTH_B17_sel_value_O),
    .out_sel(RMUX_T1_NORTH_B17_out_sel)
);
SliceWrapper_32_1_2 RMUX_T1_NORTH_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T1_NORTH_B17_sel_value_O)
);
wire [16:0] RMUX_T1_SOUTH_B17_I [1:0];
assign RMUX_T1_SOUTH_B17_I[1] = REG_T1_SOUTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T1_SOUTH_B17_I[0] = MUX_SB_T1_SOUTH_SB_OUT_B17_O;
wire [1:0] RMUX_T1_SOUTH_B17_valid_in;
assign RMUX_T1_SOUTH_B17_valid_in = {REG_T1_SOUTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T1_SOUTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T1_SOUTH_B17 (
    .I(RMUX_T1_SOUTH_B17_I),
    .O(RMUX_T1_SOUTH_B17_O),
    .ready_in(SB_T1_SOUTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T1_SOUTH_B17_ready_out),
    .valid_in(RMUX_T1_SOUTH_B17_valid_in),
    .valid_out(RMUX_T1_SOUTH_B17_valid_out),
    .S(RMUX_T1_SOUTH_B17_sel_value_O),
    .out_sel(RMUX_T1_SOUTH_B17_out_sel)
);
SliceWrapper_32_2_3 RMUX_T1_SOUTH_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T1_SOUTH_B17_sel_value_O)
);
wire [16:0] RMUX_T1_WEST_B17_I [1:0];
assign RMUX_T1_WEST_B17_I[1] = REG_T1_WEST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T1_WEST_B17_I[0] = MUX_SB_T1_WEST_SB_OUT_B17_O;
wire [1:0] RMUX_T1_WEST_B17_valid_in;
assign RMUX_T1_WEST_B17_valid_in = {REG_T1_WEST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T1_WEST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T1_WEST_B17 (
    .I(RMUX_T1_WEST_B17_I),
    .O(RMUX_T1_WEST_B17_O),
    .ready_in(SB_T1_WEST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T1_WEST_B17_ready_out),
    .valid_in(RMUX_T1_WEST_B17_valid_in),
    .valid_out(RMUX_T1_WEST_B17_valid_out),
    .S(RMUX_T1_WEST_B17_sel_value_O),
    .out_sel(RMUX_T1_WEST_B17_out_sel)
);
SliceWrapper_32_3_4 RMUX_T1_WEST_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T1_WEST_B17_sel_value_O)
);
wire [16:0] RMUX_T2_EAST_B17_I [1:0];
assign RMUX_T2_EAST_B17_I[1] = REG_T2_EAST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T2_EAST_B17_I[0] = MUX_SB_T2_EAST_SB_OUT_B17_O;
wire [1:0] RMUX_T2_EAST_B17_valid_in;
assign RMUX_T2_EAST_B17_valid_in = {REG_T2_EAST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T2_EAST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T2_EAST_B17 (
    .I(RMUX_T2_EAST_B17_I),
    .O(RMUX_T2_EAST_B17_O),
    .ready_in(SB_T2_EAST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T2_EAST_B17_ready_out),
    .valid_in(RMUX_T2_EAST_B17_valid_in),
    .valid_out(RMUX_T2_EAST_B17_valid_out),
    .S(RMUX_T2_EAST_B17_sel_value_O),
    .out_sel(RMUX_T2_EAST_B17_out_sel)
);
SliceWrapper_32_4_5 RMUX_T2_EAST_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T2_EAST_B17_sel_value_O)
);
wire [16:0] RMUX_T2_NORTH_B17_I [1:0];
assign RMUX_T2_NORTH_B17_I[1] = REG_T2_NORTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T2_NORTH_B17_I[0] = MUX_SB_T2_NORTH_SB_OUT_B17_O;
wire [1:0] RMUX_T2_NORTH_B17_valid_in;
assign RMUX_T2_NORTH_B17_valid_in = {REG_T2_NORTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T2_NORTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T2_NORTH_B17 (
    .I(RMUX_T2_NORTH_B17_I),
    .O(RMUX_T2_NORTH_B17_O),
    .ready_in(SB_T2_NORTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T2_NORTH_B17_ready_out),
    .valid_in(RMUX_T2_NORTH_B17_valid_in),
    .valid_out(RMUX_T2_NORTH_B17_valid_out),
    .S(RMUX_T2_NORTH_B17_sel_value_O),
    .out_sel(RMUX_T2_NORTH_B17_out_sel)
);
SliceWrapper_32_5_6 RMUX_T2_NORTH_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T2_NORTH_B17_sel_value_O)
);
wire [16:0] RMUX_T2_SOUTH_B17_I [1:0];
assign RMUX_T2_SOUTH_B17_I[1] = REG_T2_SOUTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T2_SOUTH_B17_I[0] = MUX_SB_T2_SOUTH_SB_OUT_B17_O;
wire [1:0] RMUX_T2_SOUTH_B17_valid_in;
assign RMUX_T2_SOUTH_B17_valid_in = {REG_T2_SOUTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T2_SOUTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T2_SOUTH_B17 (
    .I(RMUX_T2_SOUTH_B17_I),
    .O(RMUX_T2_SOUTH_B17_O),
    .ready_in(SB_T2_SOUTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T2_SOUTH_B17_ready_out),
    .valid_in(RMUX_T2_SOUTH_B17_valid_in),
    .valid_out(RMUX_T2_SOUTH_B17_valid_out),
    .S(RMUX_T2_SOUTH_B17_sel_value_O),
    .out_sel(RMUX_T2_SOUTH_B17_out_sel)
);
SliceWrapper_32_6_7 RMUX_T2_SOUTH_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T2_SOUTH_B17_sel_value_O)
);
wire [16:0] RMUX_T2_WEST_B17_I [1:0];
assign RMUX_T2_WEST_B17_I[1] = REG_T2_WEST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T2_WEST_B17_I[0] = MUX_SB_T2_WEST_SB_OUT_B17_O;
wire [1:0] RMUX_T2_WEST_B17_valid_in;
assign RMUX_T2_WEST_B17_valid_in = {REG_T2_WEST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T2_WEST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T2_WEST_B17 (
    .I(RMUX_T2_WEST_B17_I),
    .O(RMUX_T2_WEST_B17_O),
    .ready_in(SB_T2_WEST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T2_WEST_B17_ready_out),
    .valid_in(RMUX_T2_WEST_B17_valid_in),
    .valid_out(RMUX_T2_WEST_B17_valid_out),
    .S(RMUX_T2_WEST_B17_sel_value_O),
    .out_sel(RMUX_T2_WEST_B17_out_sel)
);
SliceWrapper_32_7_8 RMUX_T2_WEST_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T2_WEST_B17_sel_value_O)
);
wire [16:0] RMUX_T3_EAST_B17_I [1:0];
assign RMUX_T3_EAST_B17_I[1] = REG_T3_EAST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T3_EAST_B17_I[0] = MUX_SB_T3_EAST_SB_OUT_B17_O;
wire [1:0] RMUX_T3_EAST_B17_valid_in;
assign RMUX_T3_EAST_B17_valid_in = {REG_T3_EAST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T3_EAST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T3_EAST_B17 (
    .I(RMUX_T3_EAST_B17_I),
    .O(RMUX_T3_EAST_B17_O),
    .ready_in(SB_T3_EAST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T3_EAST_B17_ready_out),
    .valid_in(RMUX_T3_EAST_B17_valid_in),
    .valid_out(RMUX_T3_EAST_B17_valid_out),
    .S(RMUX_T3_EAST_B17_sel_value_O),
    .out_sel(RMUX_T3_EAST_B17_out_sel)
);
SliceWrapper_32_8_9 RMUX_T3_EAST_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T3_EAST_B17_sel_value_O)
);
wire [16:0] RMUX_T3_NORTH_B17_I [1:0];
assign RMUX_T3_NORTH_B17_I[1] = REG_T3_NORTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T3_NORTH_B17_I[0] = MUX_SB_T3_NORTH_SB_OUT_B17_O;
wire [1:0] RMUX_T3_NORTH_B17_valid_in;
assign RMUX_T3_NORTH_B17_valid_in = {REG_T3_NORTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T3_NORTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T3_NORTH_B17 (
    .I(RMUX_T3_NORTH_B17_I),
    .O(RMUX_T3_NORTH_B17_O),
    .ready_in(SB_T3_NORTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T3_NORTH_B17_ready_out),
    .valid_in(RMUX_T3_NORTH_B17_valid_in),
    .valid_out(RMUX_T3_NORTH_B17_valid_out),
    .S(RMUX_T3_NORTH_B17_sel_value_O),
    .out_sel(RMUX_T3_NORTH_B17_out_sel)
);
SliceWrapper_32_9_10 RMUX_T3_NORTH_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T3_NORTH_B17_sel_value_O)
);
wire [16:0] RMUX_T3_SOUTH_B17_I [1:0];
assign RMUX_T3_SOUTH_B17_I[1] = REG_T3_SOUTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T3_SOUTH_B17_I[0] = MUX_SB_T3_SOUTH_SB_OUT_B17_O;
wire [1:0] RMUX_T3_SOUTH_B17_valid_in;
assign RMUX_T3_SOUTH_B17_valid_in = {REG_T3_SOUTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T3_SOUTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T3_SOUTH_B17 (
    .I(RMUX_T3_SOUTH_B17_I),
    .O(RMUX_T3_SOUTH_B17_O),
    .ready_in(SB_T3_SOUTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T3_SOUTH_B17_ready_out),
    .valid_in(RMUX_T3_SOUTH_B17_valid_in),
    .valid_out(RMUX_T3_SOUTH_B17_valid_out),
    .S(RMUX_T3_SOUTH_B17_sel_value_O),
    .out_sel(RMUX_T3_SOUTH_B17_out_sel)
);
SliceWrapper_32_10_11 RMUX_T3_SOUTH_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T3_SOUTH_B17_sel_value_O)
);
wire [16:0] RMUX_T3_WEST_B17_I [1:0];
assign RMUX_T3_WEST_B17_I[1] = REG_T3_WEST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T3_WEST_B17_I[0] = MUX_SB_T3_WEST_SB_OUT_B17_O;
wire [1:0] RMUX_T3_WEST_B17_valid_in;
assign RMUX_T3_WEST_B17_valid_in = {REG_T3_WEST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T3_WEST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T3_WEST_B17 (
    .I(RMUX_T3_WEST_B17_I),
    .O(RMUX_T3_WEST_B17_O),
    .ready_in(SB_T3_WEST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T3_WEST_B17_ready_out),
    .valid_in(RMUX_T3_WEST_B17_valid_in),
    .valid_out(RMUX_T3_WEST_B17_valid_out),
    .S(RMUX_T3_WEST_B17_sel_value_O),
    .out_sel(RMUX_T3_WEST_B17_out_sel)
);
SliceWrapper_32_11_12 RMUX_T3_WEST_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T3_WEST_B17_sel_value_O)
);
wire [16:0] RMUX_T4_EAST_B17_I [1:0];
assign RMUX_T4_EAST_B17_I[1] = REG_T4_EAST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T4_EAST_B17_I[0] = MUX_SB_T4_EAST_SB_OUT_B17_O;
wire [1:0] RMUX_T4_EAST_B17_valid_in;
assign RMUX_T4_EAST_B17_valid_in = {REG_T4_EAST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T4_EAST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T4_EAST_B17 (
    .I(RMUX_T4_EAST_B17_I),
    .O(RMUX_T4_EAST_B17_O),
    .ready_in(SB_T4_EAST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T4_EAST_B17_ready_out),
    .valid_in(RMUX_T4_EAST_B17_valid_in),
    .valid_out(RMUX_T4_EAST_B17_valid_out),
    .S(RMUX_T4_EAST_B17_sel_value_O),
    .out_sel(RMUX_T4_EAST_B17_out_sel)
);
SliceWrapper_32_12_13 RMUX_T4_EAST_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T4_EAST_B17_sel_value_O)
);
wire [16:0] RMUX_T4_NORTH_B17_I [1:0];
assign RMUX_T4_NORTH_B17_I[1] = REG_T4_NORTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T4_NORTH_B17_I[0] = MUX_SB_T4_NORTH_SB_OUT_B17_O;
wire [1:0] RMUX_T4_NORTH_B17_valid_in;
assign RMUX_T4_NORTH_B17_valid_in = {REG_T4_NORTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T4_NORTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T4_NORTH_B17 (
    .I(RMUX_T4_NORTH_B17_I),
    .O(RMUX_T4_NORTH_B17_O),
    .ready_in(SB_T4_NORTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T4_NORTH_B17_ready_out),
    .valid_in(RMUX_T4_NORTH_B17_valid_in),
    .valid_out(RMUX_T4_NORTH_B17_valid_out),
    .S(RMUX_T4_NORTH_B17_sel_value_O),
    .out_sel(RMUX_T4_NORTH_B17_out_sel)
);
SliceWrapper_32_13_14 RMUX_T4_NORTH_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T4_NORTH_B17_sel_value_O)
);
wire [16:0] RMUX_T4_SOUTH_B17_I [1:0];
assign RMUX_T4_SOUTH_B17_I[1] = REG_T4_SOUTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T4_SOUTH_B17_I[0] = MUX_SB_T4_SOUTH_SB_OUT_B17_O;
wire [1:0] RMUX_T4_SOUTH_B17_valid_in;
assign RMUX_T4_SOUTH_B17_valid_in = {REG_T4_SOUTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T4_SOUTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T4_SOUTH_B17 (
    .I(RMUX_T4_SOUTH_B17_I),
    .O(RMUX_T4_SOUTH_B17_O),
    .ready_in(SB_T4_SOUTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T4_SOUTH_B17_ready_out),
    .valid_in(RMUX_T4_SOUTH_B17_valid_in),
    .valid_out(RMUX_T4_SOUTH_B17_valid_out),
    .S(RMUX_T4_SOUTH_B17_sel_value_O),
    .out_sel(RMUX_T4_SOUTH_B17_out_sel)
);
SliceWrapper_32_14_15 RMUX_T4_SOUTH_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T4_SOUTH_B17_sel_value_O)
);
wire [16:0] RMUX_T4_WEST_B17_I [1:0];
assign RMUX_T4_WEST_B17_I[1] = REG_T4_WEST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T4_WEST_B17_I[0] = MUX_SB_T4_WEST_SB_OUT_B17_O;
wire [1:0] RMUX_T4_WEST_B17_valid_in;
assign RMUX_T4_WEST_B17_valid_in = {REG_T4_WEST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T4_WEST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T4_WEST_B17 (
    .I(RMUX_T4_WEST_B17_I),
    .O(RMUX_T4_WEST_B17_O),
    .ready_in(SB_T4_WEST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T4_WEST_B17_ready_out),
    .valid_in(RMUX_T4_WEST_B17_valid_in),
    .valid_out(RMUX_T4_WEST_B17_valid_out),
    .S(RMUX_T4_WEST_B17_sel_value_O),
    .out_sel(RMUX_T4_WEST_B17_out_sel)
);
SliceWrapper_32_15_16 RMUX_T4_WEST_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T4_WEST_B17_sel_value_O)
);
SliceWrapper_32_16_17 SB_T0_EAST_SB_IN_B17_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_EAST_SB_IN_B17_enable_value_O)
);
FanoutHash_55B00FA90A0098BB SB_T0_EAST_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T0_WEST_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T0_EAST_SB_IN_B17_fan_in_O),
    .E1(SB_T3_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T0_EAST_SB_OUT_B17_FANOUT_I;
assign SB_T0_EAST_SB_OUT_B17_FANOUT_I = {REG_T0_EAST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T0_EAST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T0_EAST_SB_OUT_B17_FANOUT (
    .S(RMUX_T0_EAST_B17_out_sel),
    .O(SB_T0_EAST_SB_OUT_B17_FANOUT_O),
    .I(SB_T0_EAST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_32_17_18 SB_T0_EAST_SB_OUT_B17_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_EAST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_32_18_21 SB_T0_EAST_SB_OUT_B17_sel_value (
    .I(config_reg_2_O),
    .O(SB_T0_EAST_SB_OUT_B17_sel_value_O)
);
SliceWrapper_32_21_22 SB_T0_NORTH_SB_IN_B17_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_NORTH_SB_IN_B17_enable_value_O)
);
FanoutHash_3A6A5822E84DCC71 SB_T0_NORTH_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T0_WEST_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T0_NORTH_SB_IN_B17_fan_in_O),
    .E1(SB_T1_EAST_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T0_NORTH_SB_OUT_B17_FANOUT_I;
assign SB_T0_NORTH_SB_OUT_B17_FANOUT_I = {REG_T0_NORTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T0_NORTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T0_NORTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T0_NORTH_B17_out_sel),
    .O(SB_T0_NORTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T0_NORTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_32_22_23 SB_T0_NORTH_SB_OUT_B17_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_NORTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_32_23_26 SB_T0_NORTH_SB_OUT_B17_sel_value (
    .I(config_reg_2_O),
    .O(SB_T0_NORTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_32_26_27 SB_T0_SOUTH_SB_IN_B17_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_SOUTH_SB_IN_B17_enable_value_O)
);
FanoutHash_3E05574A9CE9CA8A SB_T0_SOUTH_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T1_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T3_EAST_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T0_SOUTH_SB_IN_B17_fan_in_O),
    .E1(SB_T0_NORTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T0_SOUTH_SB_OUT_B17_FANOUT_I;
assign SB_T0_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T0_SOUTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T0_SOUTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T0_SOUTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T0_SOUTH_B17_out_sel),
    .O(SB_T0_SOUTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T0_SOUTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_32_27_28 SB_T0_SOUTH_SB_OUT_B17_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_SOUTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_32_28_31 SB_T0_SOUTH_SB_OUT_B17_sel_value (
    .I(config_reg_2_O),
    .O(SB_T0_SOUTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_32_31_32 SB_T0_WEST_SB_IN_B17_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_WEST_SB_IN_B17_enable_value_O)
);
FanoutHash_87642A353688B49 SB_T0_WEST_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T0_EAST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T0_WEST_SB_IN_B17_fan_in_O),
    .E1(SB_T4_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T0_WEST_SB_OUT_B17_FANOUT_I;
assign SB_T0_WEST_SB_OUT_B17_FANOUT_I = {REG_T0_WEST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T0_WEST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T0_WEST_SB_OUT_B17_FANOUT (
    .S(RMUX_T0_WEST_B17_out_sel),
    .O(SB_T0_WEST_SB_OUT_B17_FANOUT_O),
    .I(SB_T0_WEST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_31_0_1 SB_T0_WEST_SB_OUT_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T0_WEST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_31_1_4 SB_T0_WEST_SB_OUT_B17_sel_value (
    .I(config_reg_3_O),
    .O(SB_T0_WEST_SB_OUT_B17_sel_value_O)
);
SliceWrapper_31_4_5 SB_T1_EAST_SB_IN_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_EAST_SB_IN_B17_enable_value_O)
);
FanoutHash_245560850976C879 SB_T1_EAST_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T1_EAST_SB_IN_B17_fan_in_O),
    .E1(SB_T1_WEST_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T1_EAST_SB_OUT_B17_FANOUT_I;
assign SB_T1_EAST_SB_OUT_B17_FANOUT_I = {REG_T1_EAST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T1_EAST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T1_EAST_SB_OUT_B17_FANOUT (
    .S(RMUX_T1_EAST_B17_out_sel),
    .O(SB_T1_EAST_SB_OUT_B17_FANOUT_O),
    .I(SB_T1_EAST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_31_5_6 SB_T1_EAST_SB_OUT_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_EAST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_31_6_9 SB_T1_EAST_SB_OUT_B17_sel_value (
    .I(config_reg_3_O),
    .O(SB_T1_EAST_SB_OUT_B17_sel_value_O)
);
SliceWrapper_31_9_10 SB_T1_NORTH_SB_IN_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_NORTH_SB_IN_B17_enable_value_O)
);
FanoutHash_37E9FE88073C5BAC SB_T1_NORTH_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T4_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T2_EAST_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T1_NORTH_SB_IN_B17_fan_in_O),
    .E1(SB_T1_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T1_NORTH_SB_OUT_B17_FANOUT_I;
assign SB_T1_NORTH_SB_OUT_B17_FANOUT_I = {REG_T1_NORTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T1_NORTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T1_NORTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T1_NORTH_B17_out_sel),
    .O(SB_T1_NORTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T1_NORTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_31_10_11 SB_T1_NORTH_SB_OUT_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_NORTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_31_11_14 SB_T1_NORTH_SB_OUT_B17_sel_value (
    .I(config_reg_3_O),
    .O(SB_T1_NORTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_31_14_15 SB_T1_SOUTH_SB_IN_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_SOUTH_SB_IN_B17_enable_value_O)
);
FanoutHash_2F92967E9F56D548 SB_T1_SOUTH_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T2_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T2_EAST_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T1_SOUTH_SB_IN_B17_fan_in_O),
    .E1(SB_T1_NORTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T1_SOUTH_SB_OUT_B17_FANOUT_I;
assign SB_T1_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T1_SOUTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T1_SOUTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T1_SOUTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T1_SOUTH_B17_out_sel),
    .O(SB_T1_SOUTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T1_SOUTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_31_15_16 SB_T1_SOUTH_SB_OUT_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_SOUTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_31_16_19 SB_T1_SOUTH_SB_OUT_B17_sel_value (
    .I(config_reg_3_O),
    .O(SB_T1_SOUTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_31_19_20 SB_T1_WEST_SB_IN_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_WEST_SB_IN_B17_enable_value_O)
);
FanoutHash_653384C8EF52B5E3 SB_T1_WEST_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T1_EAST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T1_WEST_SB_IN_B17_fan_in_O),
    .E1(SB_T0_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T1_WEST_SB_OUT_B17_FANOUT_I;
assign SB_T1_WEST_SB_OUT_B17_FANOUT_I = {REG_T1_WEST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T1_WEST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T1_WEST_SB_OUT_B17_FANOUT (
    .S(RMUX_T1_WEST_B17_out_sel),
    .O(SB_T1_WEST_SB_OUT_B17_FANOUT_O),
    .I(SB_T1_WEST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_31_20_21 SB_T1_WEST_SB_OUT_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_WEST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_31_21_24 SB_T1_WEST_SB_OUT_B17_sel_value (
    .I(config_reg_3_O),
    .O(SB_T1_WEST_SB_OUT_B17_sel_value_O)
);
SliceWrapper_31_24_25 SB_T2_EAST_SB_IN_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T2_EAST_SB_IN_B17_enable_value_O)
);
FanoutHash_5CD8077D054B887B SB_T2_EAST_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T2_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T2_EAST_SB_IN_B17_fan_in_O),
    .E1(SB_T1_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T2_EAST_SB_OUT_B17_FANOUT_I;
assign SB_T2_EAST_SB_OUT_B17_FANOUT_I = {REG_T2_EAST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T2_EAST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T2_EAST_SB_OUT_B17_FANOUT (
    .S(RMUX_T2_EAST_B17_out_sel),
    .O(SB_T2_EAST_SB_OUT_B17_FANOUT_O),
    .I(SB_T2_EAST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_31_25_26 SB_T2_EAST_SB_OUT_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T2_EAST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_31_26_29 SB_T2_EAST_SB_OUT_B17_sel_value (
    .I(config_reg_3_O),
    .O(SB_T2_EAST_SB_OUT_B17_sel_value_O)
);
SliceWrapper_31_29_30 SB_T2_NORTH_SB_IN_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T2_NORTH_SB_IN_B17_enable_value_O)
);
FanoutHash_74A3E41836ECED62 SB_T2_NORTH_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T3_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T3_EAST_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T2_NORTH_SB_IN_B17_fan_in_O),
    .E1(SB_T2_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T2_NORTH_SB_OUT_B17_FANOUT_I;
assign SB_T2_NORTH_SB_OUT_B17_FANOUT_I = {REG_T2_NORTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T2_NORTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T2_NORTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T2_NORTH_B17_out_sel),
    .O(SB_T2_NORTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T2_NORTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_31_30_31 SB_T2_NORTH_SB_OUT_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T2_NORTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_30_0_3 SB_T2_NORTH_SB_OUT_B17_sel_value (
    .I(config_reg_4_O),
    .O(SB_T2_NORTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_30_3_4 SB_T2_SOUTH_SB_IN_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T2_SOUTH_SB_IN_B17_enable_value_O)
);
FanoutHash_2CE3041FDDDDEC1A SB_T2_SOUTH_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T3_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T1_EAST_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T2_SOUTH_SB_IN_B17_fan_in_O),
    .E1(SB_T2_NORTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T2_SOUTH_SB_OUT_B17_FANOUT_I;
assign SB_T2_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T2_SOUTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T2_SOUTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T2_SOUTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T2_SOUTH_B17_out_sel),
    .O(SB_T2_SOUTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T2_SOUTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_30_4_5 SB_T2_SOUTH_SB_OUT_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T2_SOUTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_30_5_8 SB_T2_SOUTH_SB_OUT_B17_sel_value (
    .I(config_reg_4_O),
    .O(SB_T2_SOUTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_30_8_9 SB_T2_WEST_SB_IN_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T2_WEST_SB_IN_B17_enable_value_O)
);
FanoutHash_4A74B16B611BA7E4 SB_T2_WEST_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T2_EAST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T2_WEST_SB_IN_B17_fan_in_O),
    .E1(SB_T1_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T2_WEST_SB_OUT_B17_FANOUT_I;
assign SB_T2_WEST_SB_OUT_B17_FANOUT_I = {REG_T2_WEST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T2_WEST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T2_WEST_SB_OUT_B17_FANOUT (
    .S(RMUX_T2_WEST_B17_out_sel),
    .O(SB_T2_WEST_SB_OUT_B17_FANOUT_O),
    .I(SB_T2_WEST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_30_9_10 SB_T2_WEST_SB_OUT_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T2_WEST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_30_10_13 SB_T2_WEST_SB_OUT_B17_sel_value (
    .I(config_reg_4_O),
    .O(SB_T2_WEST_SB_OUT_B17_sel_value_O)
);
SliceWrapper_30_13_14 SB_T3_EAST_SB_IN_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_EAST_SB_IN_B17_enable_value_O)
);
FanoutHash_276F8381CE025648 SB_T3_EAST_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T3_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T3_EAST_SB_IN_B17_fan_in_O),
    .E1(SB_T2_NORTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T3_EAST_SB_OUT_B17_FANOUT_I;
assign SB_T3_EAST_SB_OUT_B17_FANOUT_I = {REG_T3_EAST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T3_EAST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T3_EAST_SB_OUT_B17_FANOUT (
    .S(RMUX_T3_EAST_B17_out_sel),
    .O(SB_T3_EAST_SB_OUT_B17_FANOUT_O),
    .I(SB_T3_EAST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_30_14_15 SB_T3_EAST_SB_OUT_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_EAST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_30_15_18 SB_T3_EAST_SB_OUT_B17_sel_value (
    .I(config_reg_4_O),
    .O(SB_T3_EAST_SB_OUT_B17_sel_value_O)
);
SliceWrapper_30_18_19 SB_T3_NORTH_SB_IN_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_NORTH_SB_IN_B17_enable_value_O)
);
FanoutHash_7E22D83B42537D1D SB_T3_NORTH_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T2_WEST_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T3_NORTH_SB_IN_B17_fan_in_O),
    .E1(SB_T4_EAST_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T3_NORTH_SB_OUT_B17_FANOUT_I;
assign SB_T3_NORTH_SB_OUT_B17_FANOUT_I = {REG_T3_NORTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T3_NORTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T3_NORTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T3_NORTH_B17_out_sel),
    .O(SB_T3_NORTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T3_NORTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_30_19_20 SB_T3_NORTH_SB_OUT_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_NORTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_30_20_23 SB_T3_NORTH_SB_OUT_B17_sel_value (
    .I(config_reg_4_O),
    .O(SB_T3_NORTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_30_23_24 SB_T3_SOUTH_SB_IN_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_SOUTH_SB_IN_B17_enable_value_O)
);
FanoutHash_59B7E37DAE2221E3 SB_T3_SOUTH_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T4_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T0_EAST_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T3_SOUTH_SB_IN_B17_fan_in_O),
    .E1(SB_T3_NORTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T3_SOUTH_SB_OUT_B17_FANOUT_I;
assign SB_T3_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T3_SOUTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T3_SOUTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T3_SOUTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T3_SOUTH_B17_out_sel),
    .O(SB_T3_SOUTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T3_SOUTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_30_24_25 SB_T3_SOUTH_SB_OUT_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_SOUTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_30_25_28 SB_T3_SOUTH_SB_OUT_B17_sel_value (
    .I(config_reg_4_O),
    .O(SB_T3_SOUTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_30_28_29 SB_T3_WEST_SB_IN_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_WEST_SB_IN_B17_enable_value_O)
);
FanoutHash_41D739158D58E184 SB_T3_WEST_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T3_EAST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T3_WEST_SB_IN_B17_fan_in_O),
    .E1(SB_T2_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T3_WEST_SB_OUT_B17_FANOUT_I;
assign SB_T3_WEST_SB_OUT_B17_FANOUT_I = {REG_T3_WEST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T3_WEST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T3_WEST_SB_OUT_B17_FANOUT (
    .S(RMUX_T3_WEST_B17_out_sel),
    .O(SB_T3_WEST_SB_OUT_B17_FANOUT_O),
    .I(SB_T3_WEST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_30_29_30 SB_T3_WEST_SB_OUT_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_WEST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_23_0_3 SB_T3_WEST_SB_OUT_B17_sel_value (
    .I(config_reg_5_O),
    .O(SB_T3_WEST_SB_OUT_B17_sel_value_O)
);
SliceWrapper_23_3_4 SB_T4_EAST_SB_IN_B17_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_EAST_SB_IN_B17_enable_value_O)
);
FanoutHash_55169EB19E10AA09 SB_T4_EAST_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T4_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T4_EAST_SB_IN_B17_fan_in_O),
    .E1(SB_T4_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T4_EAST_SB_OUT_B17_FANOUT_I;
assign SB_T4_EAST_SB_OUT_B17_FANOUT_I = {REG_T4_EAST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T4_EAST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T4_EAST_SB_OUT_B17_FANOUT (
    .S(RMUX_T4_EAST_B17_out_sel),
    .O(SB_T4_EAST_SB_OUT_B17_FANOUT_O),
    .I(SB_T4_EAST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_23_4_5 SB_T4_EAST_SB_OUT_B17_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_EAST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_23_5_8 SB_T4_EAST_SB_OUT_B17_sel_value (
    .I(config_reg_5_O),
    .O(SB_T4_EAST_SB_OUT_B17_sel_value_O)
);
SliceWrapper_23_8_9 SB_T4_NORTH_SB_IN_B17_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_NORTH_SB_IN_B17_enable_value_O)
);
FanoutHash_244497FCED8BEB80 SB_T4_NORTH_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T1_WEST_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T4_NORTH_SB_IN_B17_fan_in_O),
    .E1(SB_T0_EAST_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T4_NORTH_SB_OUT_B17_FANOUT_I;
assign SB_T4_NORTH_SB_OUT_B17_FANOUT_I = {REG_T4_NORTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T4_NORTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T4_NORTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T4_NORTH_B17_out_sel),
    .O(SB_T4_NORTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T4_NORTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_23_9_10 SB_T4_NORTH_SB_OUT_B17_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_NORTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_23_10_13 SB_T4_NORTH_SB_OUT_B17_sel_value (
    .I(config_reg_5_O),
    .O(SB_T4_NORTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_23_13_14 SB_T4_SOUTH_SB_IN_B17_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_SOUTH_SB_IN_B17_enable_value_O)
);
FanoutHash_AE7392256DF8B0F SB_T4_SOUTH_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T0_WEST_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T4_SOUTH_SB_IN_B17_fan_in_O),
    .E1(SB_T4_EAST_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T4_SOUTH_SB_OUT_B17_FANOUT_I;
assign SB_T4_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T4_SOUTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T4_SOUTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T4_SOUTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T4_SOUTH_B17_out_sel),
    .O(SB_T4_SOUTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T4_SOUTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_23_14_15 SB_T4_SOUTH_SB_OUT_B17_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_SOUTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_23_15_18 SB_T4_SOUTH_SB_OUT_B17_sel_value (
    .I(config_reg_5_O),
    .O(SB_T4_SOUTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_23_18_19 SB_T4_WEST_SB_IN_B17_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_WEST_SB_IN_B17_enable_value_O)
);
FanoutHash_6E1094CE0D0F6DFA SB_T4_WEST_SB_IN_B17_fan_in (
    .S6(PE_input_width_17_num_3_out_sel),
    .E2(SB_T4_EAST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
    .E7(PondTop_input_width_17_num_0_enable),
    .I3(PE_input_width_17_num_0_ready),
    .S0(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
    .E5(PE_input_width_17_num_2_enable),
    .E8(PondTop_input_width_17_num_1_enable),
    .I6(PE_input_width_17_num_3_ready),
    .I7(PondTop_input_width_17_num_0_ready),
    .I2(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
    .S3(PE_input_width_17_num_0_out_sel),
    .S8(PondTop_input_width_17_num_1_out_sel),
    .S2(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
    .E3(PE_input_width_17_num_0_enable),
    .E0(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
    .S4(PE_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
    .S7(PondTop_input_width_17_num_0_out_sel),
    .E4(PE_input_width_17_num_1_enable),
    .S5(PE_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
    .I5(PE_input_width_17_num_2_ready),
    .E6(PE_input_width_17_num_3_enable),
    .I4(PE_input_width_17_num_1_ready),
    .I8(PondTop_input_width_17_num_1_ready),
    .O(SB_T4_WEST_SB_IN_B17_fan_in_O),
    .E1(SB_T3_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T4_WEST_SB_OUT_B17_FANOUT_I;
assign SB_T4_WEST_SB_OUT_B17_FANOUT_I = {REG_T4_WEST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T4_WEST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T4_WEST_SB_OUT_B17_FANOUT (
    .S(RMUX_T4_WEST_B17_out_sel),
    .O(SB_T4_WEST_SB_OUT_B17_FANOUT_O),
    .I(SB_T4_WEST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_23_19_20 SB_T4_WEST_SB_OUT_B17_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_WEST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_23_20_23 SB_T4_WEST_SB_OUT_B17_sel_value (
    .I(config_reg_5_O),
    .O(SB_T4_WEST_SB_OUT_B17_sel_value_O)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T0_EAST_SB_IN_B17 (
    .I(SB_T0_EAST_SB_IN_B17),
    .O(WIRE_SB_T0_EAST_SB_IN_B17_O),
    .ready_in(SB_T0_EAST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T0_EAST_SB_IN_B17_ready_out),
    .valid_in(SB_T0_EAST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T0_EAST_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T0_NORTH_SB_IN_B17 (
    .I(SB_T0_NORTH_SB_IN_B17),
    .O(WIRE_SB_T0_NORTH_SB_IN_B17_O),
    .ready_in(SB_T0_NORTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T0_NORTH_SB_IN_B17_ready_out),
    .valid_in(SB_T0_NORTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T0_NORTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T0_SOUTH_SB_IN_B17 (
    .I(SB_T0_SOUTH_SB_IN_B17),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B17_O),
    .ready_in(SB_T0_SOUTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T0_SOUTH_SB_IN_B17_ready_out),
    .valid_in(SB_T0_SOUTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T0_WEST_SB_IN_B17 (
    .I(SB_T0_WEST_SB_IN_B17),
    .O(WIRE_SB_T0_WEST_SB_IN_B17_O),
    .ready_in(SB_T0_WEST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T0_WEST_SB_IN_B17_ready_out),
    .valid_in(SB_T0_WEST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T0_WEST_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T1_EAST_SB_IN_B17 (
    .I(SB_T1_EAST_SB_IN_B17),
    .O(WIRE_SB_T1_EAST_SB_IN_B17_O),
    .ready_in(SB_T1_EAST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T1_EAST_SB_IN_B17_ready_out),
    .valid_in(SB_T1_EAST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T1_EAST_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T1_NORTH_SB_IN_B17 (
    .I(SB_T1_NORTH_SB_IN_B17),
    .O(WIRE_SB_T1_NORTH_SB_IN_B17_O),
    .ready_in(SB_T1_NORTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T1_NORTH_SB_IN_B17_ready_out),
    .valid_in(SB_T1_NORTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T1_NORTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T1_SOUTH_SB_IN_B17 (
    .I(SB_T1_SOUTH_SB_IN_B17),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B17_O),
    .ready_in(SB_T1_SOUTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T1_SOUTH_SB_IN_B17_ready_out),
    .valid_in(SB_T1_SOUTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T1_WEST_SB_IN_B17 (
    .I(SB_T1_WEST_SB_IN_B17),
    .O(WIRE_SB_T1_WEST_SB_IN_B17_O),
    .ready_in(SB_T1_WEST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T1_WEST_SB_IN_B17_ready_out),
    .valid_in(SB_T1_WEST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T1_WEST_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T2_EAST_SB_IN_B17 (
    .I(SB_T2_EAST_SB_IN_B17),
    .O(WIRE_SB_T2_EAST_SB_IN_B17_O),
    .ready_in(SB_T2_EAST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T2_EAST_SB_IN_B17_ready_out),
    .valid_in(SB_T2_EAST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T2_EAST_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T2_NORTH_SB_IN_B17 (
    .I(SB_T2_NORTH_SB_IN_B17),
    .O(WIRE_SB_T2_NORTH_SB_IN_B17_O),
    .ready_in(SB_T2_NORTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T2_NORTH_SB_IN_B17_ready_out),
    .valid_in(SB_T2_NORTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T2_NORTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T2_SOUTH_SB_IN_B17 (
    .I(SB_T2_SOUTH_SB_IN_B17),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B17_O),
    .ready_in(SB_T2_SOUTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T2_SOUTH_SB_IN_B17_ready_out),
    .valid_in(SB_T2_SOUTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T2_WEST_SB_IN_B17 (
    .I(SB_T2_WEST_SB_IN_B17),
    .O(WIRE_SB_T2_WEST_SB_IN_B17_O),
    .ready_in(SB_T2_WEST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T2_WEST_SB_IN_B17_ready_out),
    .valid_in(SB_T2_WEST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T2_WEST_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T3_EAST_SB_IN_B17 (
    .I(SB_T3_EAST_SB_IN_B17),
    .O(WIRE_SB_T3_EAST_SB_IN_B17_O),
    .ready_in(SB_T3_EAST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T3_EAST_SB_IN_B17_ready_out),
    .valid_in(SB_T3_EAST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T3_EAST_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T3_NORTH_SB_IN_B17 (
    .I(SB_T3_NORTH_SB_IN_B17),
    .O(WIRE_SB_T3_NORTH_SB_IN_B17_O),
    .ready_in(SB_T3_NORTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T3_NORTH_SB_IN_B17_ready_out),
    .valid_in(SB_T3_NORTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T3_NORTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T3_SOUTH_SB_IN_B17 (
    .I(SB_T3_SOUTH_SB_IN_B17),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B17_O),
    .ready_in(SB_T3_SOUTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T3_SOUTH_SB_IN_B17_ready_out),
    .valid_in(SB_T3_SOUTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T3_WEST_SB_IN_B17 (
    .I(SB_T3_WEST_SB_IN_B17),
    .O(WIRE_SB_T3_WEST_SB_IN_B17_O),
    .ready_in(SB_T3_WEST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T3_WEST_SB_IN_B17_ready_out),
    .valid_in(SB_T3_WEST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T3_WEST_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T4_EAST_SB_IN_B17 (
    .I(SB_T4_EAST_SB_IN_B17),
    .O(WIRE_SB_T4_EAST_SB_IN_B17_O),
    .ready_in(SB_T4_EAST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T4_EAST_SB_IN_B17_ready_out),
    .valid_in(SB_T4_EAST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T4_EAST_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T4_NORTH_SB_IN_B17 (
    .I(SB_T4_NORTH_SB_IN_B17),
    .O(WIRE_SB_T4_NORTH_SB_IN_B17_O),
    .ready_in(SB_T4_NORTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T4_NORTH_SB_IN_B17_ready_out),
    .valid_in(SB_T4_NORTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T4_NORTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T4_SOUTH_SB_IN_B17 (
    .I(SB_T4_SOUTH_SB_IN_B17),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B17_O),
    .ready_in(SB_T4_SOUTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T4_SOUTH_SB_IN_B17_ready_out),
    .valid_in(SB_T4_SOUTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T4_WEST_SB_IN_B17 (
    .I(SB_T4_WEST_SB_IN_B17),
    .O(WIRE_SB_T4_WEST_SB_IN_B17_O),
    .ready_in(SB_T4_WEST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T4_WEST_SB_IN_B17_ready_out),
    .valid_in(SB_T4_WEST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T4_WEST_SB_IN_B17_valid_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_23_32_inst0$bit_const_0_None (
    .out(ZextWrapper_23_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_23_32_inst0$self_O_out;
assign ZextWrapper_23_32_inst0$self_O_out = {ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,config_reg_5_O};
mantle_wire__typeBitIn32 ZextWrapper_23_32_inst0$self_O (
    .in(ZextWrapper_23_32_inst0$self_O_in),
    .out(ZextWrapper_23_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_30_32_inst0$bit_const_0_None (
    .out(ZextWrapper_30_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_30_32_inst0$self_O_out;
assign ZextWrapper_30_32_inst0$self_O_out = {ZextWrapper_30_32_inst0$bit_const_0_None_out,ZextWrapper_30_32_inst0$bit_const_0_None_out,config_reg_4_O};
mantle_wire__typeBitIn32 ZextWrapper_30_32_inst0$self_O (
    .in(ZextWrapper_30_32_inst0$self_O_in),
    .out(ZextWrapper_30_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_31_32_inst0$bit_const_0_None (
    .out(ZextWrapper_31_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_31_32_inst0$self_O_out;
assign ZextWrapper_31_32_inst0$self_O_out = {ZextWrapper_31_32_inst0$bit_const_0_None_out,config_reg_3_O};
mantle_wire__typeBitIn32 ZextWrapper_31_32_inst0$self_O (
    .in(ZextWrapper_31_32_inst0$self_O_in),
    .out(ZextWrapper_31_32_inst0$self_O_out)
);
coreir_and #(
    .width(1)
) and1_inst0 (
    .in0(coreir_eq_1_inst0_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst0_out)
);
coreir_and #(
    .width(1)
) and1_inst1 (
    .in0(coreir_eq_1_inst1_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst1_out)
);
coreir_and #(
    .width(1)
) and1_inst10 (
    .in0(coreir_eq_1_inst10_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst10_out)
);
coreir_and #(
    .width(1)
) and1_inst11 (
    .in0(coreir_eq_1_inst11_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst11_out)
);
coreir_and #(
    .width(1)
) and1_inst12 (
    .in0(coreir_eq_1_inst12_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst12_out)
);
coreir_and #(
    .width(1)
) and1_inst13 (
    .in0(coreir_eq_1_inst13_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst13_out)
);
coreir_and #(
    .width(1)
) and1_inst14 (
    .in0(coreir_eq_1_inst14_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst14_out)
);
coreir_and #(
    .width(1)
) and1_inst15 (
    .in0(coreir_eq_1_inst15_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst15_out)
);
coreir_and #(
    .width(1)
) and1_inst16 (
    .in0(coreir_eq_1_inst16_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst16_out)
);
coreir_and #(
    .width(1)
) and1_inst17 (
    .in0(coreir_eq_1_inst17_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst17_out)
);
coreir_and #(
    .width(1)
) and1_inst18 (
    .in0(coreir_eq_1_inst18_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst18_out)
);
coreir_and #(
    .width(1)
) and1_inst19 (
    .in0(coreir_eq_1_inst19_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst19_out)
);
coreir_and #(
    .width(1)
) and1_inst2 (
    .in0(coreir_eq_1_inst2_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst2_out)
);
coreir_and #(
    .width(1)
) and1_inst3 (
    .in0(coreir_eq_1_inst3_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst3_out)
);
coreir_and #(
    .width(1)
) and1_inst4 (
    .in0(coreir_eq_1_inst4_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst4_out)
);
coreir_and #(
    .width(1)
) and1_inst5 (
    .in0(coreir_eq_1_inst5_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst5_out)
);
coreir_and #(
    .width(1)
) and1_inst6 (
    .in0(coreir_eq_1_inst6_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst6_out)
);
coreir_and #(
    .width(1)
) and1_inst7 (
    .in0(coreir_eq_1_inst7_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst7_out)
);
coreir_and #(
    .width(1)
) and1_inst8 (
    .in0(coreir_eq_1_inst8_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst8_out)
);
coreir_and #(
    .width(1)
) and1_inst9 (
    .in0(coreir_eq_1_inst9_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst9_out)
);
wire [7:0] config_reg_0_config_addr;
assign config_reg_0_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_32_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_reg_0_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_1_config_addr;
assign config_reg_1_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_32_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_reg_1_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_2_config_addr;
assign config_reg_2_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_32_8_32_2 config_reg_2 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_2_O),
    .config_addr(config_reg_2_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_3_config_addr;
assign config_reg_3_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_31_8_32_3 config_reg_3 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_3_O),
    .config_addr(config_reg_3_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_4_config_addr;
assign config_reg_4_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_30_8_32_4 config_reg_4 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_4_O),
    .config_addr(config_reg_4_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_5_config_addr;
assign config_reg_5_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_23_8_32_5 config_reg_5 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_5_O),
    .config_addr(config_reg_5_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst0 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_NORTH_B17_sel_value_O),
    .out(coreir_eq_1_inst0_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst1 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_SOUTH_B17_sel_value_O),
    .out(coreir_eq_1_inst1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst10 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_EAST_B17_sel_value_O),
    .out(coreir_eq_1_inst10_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst11 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_WEST_B17_sel_value_O),
    .out(coreir_eq_1_inst11_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst12 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_NORTH_B17_sel_value_O),
    .out(coreir_eq_1_inst12_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst13 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_SOUTH_B17_sel_value_O),
    .out(coreir_eq_1_inst13_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst14 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_EAST_B17_sel_value_O),
    .out(coreir_eq_1_inst14_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst15 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_WEST_B17_sel_value_O),
    .out(coreir_eq_1_inst15_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst16 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_NORTH_B17_sel_value_O),
    .out(coreir_eq_1_inst16_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst17 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_SOUTH_B17_sel_value_O),
    .out(coreir_eq_1_inst17_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst18 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_EAST_B17_sel_value_O),
    .out(coreir_eq_1_inst18_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst19 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_WEST_B17_sel_value_O),
    .out(coreir_eq_1_inst19_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst2 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_EAST_B17_sel_value_O),
    .out(coreir_eq_1_inst2_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst3 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_WEST_B17_sel_value_O),
    .out(coreir_eq_1_inst3_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst4 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_NORTH_B17_sel_value_O),
    .out(coreir_eq_1_inst4_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst5 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_SOUTH_B17_sel_value_O),
    .out(coreir_eq_1_inst5_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst6 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_EAST_B17_sel_value_O),
    .out(coreir_eq_1_inst6_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst7 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_WEST_B17_sel_value_O),
    .out(coreir_eq_1_inst7_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst8 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_NORTH_B17_sel_value_O),
    .out(coreir_eq_1_inst8_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst9 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_SOUTH_B17_sel_value_O),
    .out(coreir_eq_1_inst9_out)
);
wire [31:0] mux_aoi_6_32_inst0_I [5:0];
assign mux_aoi_6_32_inst0_I[5] = ZextWrapper_23_32_inst0$self_O_in;
assign mux_aoi_6_32_inst0_I[4] = ZextWrapper_30_32_inst0$self_O_in;
assign mux_aoi_6_32_inst0_I[3] = ZextWrapper_31_32_inst0$self_O_in;
assign mux_aoi_6_32_inst0_I[2] = config_reg_2_O;
assign mux_aoi_6_32_inst0_I[1] = config_reg_1_O;
assign mux_aoi_6_32_inst0_I[0] = config_reg_0_O;
mux_aoi_6_32 mux_aoi_6_32_inst0 (
    .I(mux_aoi_6_32_inst0_I),
    .O(mux_aoi_6_32_inst0_O),
    .S(self_config_config_addr_out[2:0]),
    .out_sel(mux_aoi_6_32_inst0_out_sel)
);
mantle_wire__typeBit8 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
assign PE_output_width_17_num_0_ready_out = CB_PE_output_width_17_num_0_fan_in_O[0];
assign PE_output_width_17_num_1_ready_out = CB_PE_output_width_17_num_1_fan_in_O[0];
assign PE_output_width_17_num_2_ready_out = CB_PE_output_width_17_num_2_fan_in_O[0];
assign PondTop_output_width_17_num_0_ready_out = CB_PondTop_output_width_17_num_0_fan_in_O[0];
assign PondTop_output_width_17_num_1_ready_out = CB_PondTop_output_width_17_num_1_fan_in_O[0];
assign SB_T0_EAST_SB_IN_B17_enable = SB_T0_EAST_SB_IN_B17_enable_value_O[0];
assign SB_T0_EAST_SB_IN_B17_ready_out = WIRE_SB_T0_EAST_SB_IN_B17_ready_out;
assign SB_T0_EAST_SB_OUT_B17 = RMUX_T0_EAST_B17_O;
assign SB_T0_EAST_SB_OUT_B17_enable = SB_T0_EAST_SB_OUT_B17_enable_value_O[0];
assign SB_T0_EAST_SB_OUT_B17_valid_out = RMUX_T0_EAST_B17_valid_out;
assign SB_T0_NORTH_SB_IN_B17_enable = SB_T0_NORTH_SB_IN_B17_enable_value_O[0];
assign SB_T0_NORTH_SB_IN_B17_ready_out = WIRE_SB_T0_NORTH_SB_IN_B17_ready_out;
assign SB_T0_NORTH_SB_OUT_B17 = RMUX_T0_NORTH_B17_O;
assign SB_T0_NORTH_SB_OUT_B17_enable = SB_T0_NORTH_SB_OUT_B17_enable_value_O[0];
assign SB_T0_NORTH_SB_OUT_B17_valid_out = RMUX_T0_NORTH_B17_valid_out;
assign SB_T0_SOUTH_SB_IN_B17_enable = SB_T0_SOUTH_SB_IN_B17_enable_value_O[0];
assign SB_T0_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T0_SOUTH_SB_IN_B17_ready_out;
assign SB_T0_SOUTH_SB_OUT_B17 = RMUX_T0_SOUTH_B17_O;
assign SB_T0_SOUTH_SB_OUT_B17_enable = SB_T0_SOUTH_SB_OUT_B17_enable_value_O[0];
assign SB_T0_SOUTH_SB_OUT_B17_valid_out = RMUX_T0_SOUTH_B17_valid_out;
assign SB_T0_WEST_SB_IN_B17_enable = SB_T0_WEST_SB_IN_B17_enable_value_O[0];
assign SB_T0_WEST_SB_IN_B17_ready_out = WIRE_SB_T0_WEST_SB_IN_B17_ready_out;
assign SB_T0_WEST_SB_OUT_B17 = RMUX_T0_WEST_B17_O;
assign SB_T0_WEST_SB_OUT_B17_enable = SB_T0_WEST_SB_OUT_B17_enable_value_O[0];
assign SB_T0_WEST_SB_OUT_B17_valid_out = RMUX_T0_WEST_B17_valid_out;
assign SB_T1_EAST_SB_IN_B17_enable = SB_T1_EAST_SB_IN_B17_enable_value_O[0];
assign SB_T1_EAST_SB_IN_B17_ready_out = WIRE_SB_T1_EAST_SB_IN_B17_ready_out;
assign SB_T1_EAST_SB_OUT_B17 = RMUX_T1_EAST_B17_O;
assign SB_T1_EAST_SB_OUT_B17_enable = SB_T1_EAST_SB_OUT_B17_enable_value_O[0];
assign SB_T1_EAST_SB_OUT_B17_valid_out = RMUX_T1_EAST_B17_valid_out;
assign SB_T1_NORTH_SB_IN_B17_enable = SB_T1_NORTH_SB_IN_B17_enable_value_O[0];
assign SB_T1_NORTH_SB_IN_B17_ready_out = WIRE_SB_T1_NORTH_SB_IN_B17_ready_out;
assign SB_T1_NORTH_SB_OUT_B17 = RMUX_T1_NORTH_B17_O;
assign SB_T1_NORTH_SB_OUT_B17_enable = SB_T1_NORTH_SB_OUT_B17_enable_value_O[0];
assign SB_T1_NORTH_SB_OUT_B17_valid_out = RMUX_T1_NORTH_B17_valid_out;
assign SB_T1_SOUTH_SB_IN_B17_enable = SB_T1_SOUTH_SB_IN_B17_enable_value_O[0];
assign SB_T1_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T1_SOUTH_SB_IN_B17_ready_out;
assign SB_T1_SOUTH_SB_OUT_B17 = RMUX_T1_SOUTH_B17_O;
assign SB_T1_SOUTH_SB_OUT_B17_enable = SB_T1_SOUTH_SB_OUT_B17_enable_value_O[0];
assign SB_T1_SOUTH_SB_OUT_B17_valid_out = RMUX_T1_SOUTH_B17_valid_out;
assign SB_T1_WEST_SB_IN_B17_enable = SB_T1_WEST_SB_IN_B17_enable_value_O[0];
assign SB_T1_WEST_SB_IN_B17_ready_out = WIRE_SB_T1_WEST_SB_IN_B17_ready_out;
assign SB_T1_WEST_SB_OUT_B17 = RMUX_T1_WEST_B17_O;
assign SB_T1_WEST_SB_OUT_B17_enable = SB_T1_WEST_SB_OUT_B17_enable_value_O[0];
assign SB_T1_WEST_SB_OUT_B17_valid_out = RMUX_T1_WEST_B17_valid_out;
assign SB_T2_EAST_SB_IN_B17_enable = SB_T2_EAST_SB_IN_B17_enable_value_O[0];
assign SB_T2_EAST_SB_IN_B17_ready_out = WIRE_SB_T2_EAST_SB_IN_B17_ready_out;
assign SB_T2_EAST_SB_OUT_B17 = RMUX_T2_EAST_B17_O;
assign SB_T2_EAST_SB_OUT_B17_enable = SB_T2_EAST_SB_OUT_B17_enable_value_O[0];
assign SB_T2_EAST_SB_OUT_B17_valid_out = RMUX_T2_EAST_B17_valid_out;
assign SB_T2_NORTH_SB_IN_B17_enable = SB_T2_NORTH_SB_IN_B17_enable_value_O[0];
assign SB_T2_NORTH_SB_IN_B17_ready_out = WIRE_SB_T2_NORTH_SB_IN_B17_ready_out;
assign SB_T2_NORTH_SB_OUT_B17 = RMUX_T2_NORTH_B17_O;
assign SB_T2_NORTH_SB_OUT_B17_enable = SB_T2_NORTH_SB_OUT_B17_enable_value_O[0];
assign SB_T2_NORTH_SB_OUT_B17_valid_out = RMUX_T2_NORTH_B17_valid_out;
assign SB_T2_SOUTH_SB_IN_B17_enable = SB_T2_SOUTH_SB_IN_B17_enable_value_O[0];
assign SB_T2_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T2_SOUTH_SB_IN_B17_ready_out;
assign SB_T2_SOUTH_SB_OUT_B17 = RMUX_T2_SOUTH_B17_O;
assign SB_T2_SOUTH_SB_OUT_B17_enable = SB_T2_SOUTH_SB_OUT_B17_enable_value_O[0];
assign SB_T2_SOUTH_SB_OUT_B17_valid_out = RMUX_T2_SOUTH_B17_valid_out;
assign SB_T2_WEST_SB_IN_B17_enable = SB_T2_WEST_SB_IN_B17_enable_value_O[0];
assign SB_T2_WEST_SB_IN_B17_ready_out = WIRE_SB_T2_WEST_SB_IN_B17_ready_out;
assign SB_T2_WEST_SB_OUT_B17 = RMUX_T2_WEST_B17_O;
assign SB_T2_WEST_SB_OUT_B17_enable = SB_T2_WEST_SB_OUT_B17_enable_value_O[0];
assign SB_T2_WEST_SB_OUT_B17_valid_out = RMUX_T2_WEST_B17_valid_out;
assign SB_T3_EAST_SB_IN_B17_enable = SB_T3_EAST_SB_IN_B17_enable_value_O[0];
assign SB_T3_EAST_SB_IN_B17_ready_out = WIRE_SB_T3_EAST_SB_IN_B17_ready_out;
assign SB_T3_EAST_SB_OUT_B17 = RMUX_T3_EAST_B17_O;
assign SB_T3_EAST_SB_OUT_B17_enable = SB_T3_EAST_SB_OUT_B17_enable_value_O[0];
assign SB_T3_EAST_SB_OUT_B17_valid_out = RMUX_T3_EAST_B17_valid_out;
assign SB_T3_NORTH_SB_IN_B17_enable = SB_T3_NORTH_SB_IN_B17_enable_value_O[0];
assign SB_T3_NORTH_SB_IN_B17_ready_out = WIRE_SB_T3_NORTH_SB_IN_B17_ready_out;
assign SB_T3_NORTH_SB_OUT_B17 = RMUX_T3_NORTH_B17_O;
assign SB_T3_NORTH_SB_OUT_B17_enable = SB_T3_NORTH_SB_OUT_B17_enable_value_O[0];
assign SB_T3_NORTH_SB_OUT_B17_valid_out = RMUX_T3_NORTH_B17_valid_out;
assign SB_T3_SOUTH_SB_IN_B17_enable = SB_T3_SOUTH_SB_IN_B17_enable_value_O[0];
assign SB_T3_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T3_SOUTH_SB_IN_B17_ready_out;
assign SB_T3_SOUTH_SB_OUT_B17 = RMUX_T3_SOUTH_B17_O;
assign SB_T3_SOUTH_SB_OUT_B17_enable = SB_T3_SOUTH_SB_OUT_B17_enable_value_O[0];
assign SB_T3_SOUTH_SB_OUT_B17_valid_out = RMUX_T3_SOUTH_B17_valid_out;
assign SB_T3_WEST_SB_IN_B17_enable = SB_T3_WEST_SB_IN_B17_enable_value_O[0];
assign SB_T3_WEST_SB_IN_B17_ready_out = WIRE_SB_T3_WEST_SB_IN_B17_ready_out;
assign SB_T3_WEST_SB_OUT_B17 = RMUX_T3_WEST_B17_O;
assign SB_T3_WEST_SB_OUT_B17_enable = SB_T3_WEST_SB_OUT_B17_enable_value_O[0];
assign SB_T3_WEST_SB_OUT_B17_valid_out = RMUX_T3_WEST_B17_valid_out;
assign SB_T4_EAST_SB_IN_B17_enable = SB_T4_EAST_SB_IN_B17_enable_value_O[0];
assign SB_T4_EAST_SB_IN_B17_ready_out = WIRE_SB_T4_EAST_SB_IN_B17_ready_out;
assign SB_T4_EAST_SB_OUT_B17 = RMUX_T4_EAST_B17_O;
assign SB_T4_EAST_SB_OUT_B17_enable = SB_T4_EAST_SB_OUT_B17_enable_value_O[0];
assign SB_T4_EAST_SB_OUT_B17_valid_out = RMUX_T4_EAST_B17_valid_out;
assign SB_T4_NORTH_SB_IN_B17_enable = SB_T4_NORTH_SB_IN_B17_enable_value_O[0];
assign SB_T4_NORTH_SB_IN_B17_ready_out = WIRE_SB_T4_NORTH_SB_IN_B17_ready_out;
assign SB_T4_NORTH_SB_OUT_B17 = RMUX_T4_NORTH_B17_O;
assign SB_T4_NORTH_SB_OUT_B17_enable = SB_T4_NORTH_SB_OUT_B17_enable_value_O[0];
assign SB_T4_NORTH_SB_OUT_B17_valid_out = RMUX_T4_NORTH_B17_valid_out;
assign SB_T4_SOUTH_SB_IN_B17_enable = SB_T4_SOUTH_SB_IN_B17_enable_value_O[0];
assign SB_T4_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T4_SOUTH_SB_IN_B17_ready_out;
assign SB_T4_SOUTH_SB_OUT_B17 = RMUX_T4_SOUTH_B17_O;
assign SB_T4_SOUTH_SB_OUT_B17_enable = SB_T4_SOUTH_SB_OUT_B17_enable_value_O[0];
assign SB_T4_SOUTH_SB_OUT_B17_valid_out = RMUX_T4_SOUTH_B17_valid_out;
assign SB_T4_WEST_SB_IN_B17_enable = SB_T4_WEST_SB_IN_B17_enable_value_O[0];
assign SB_T4_WEST_SB_IN_B17_ready_out = WIRE_SB_T4_WEST_SB_IN_B17_ready_out;
assign SB_T4_WEST_SB_OUT_B17 = RMUX_T4_WEST_B17_O;
assign SB_T4_WEST_SB_OUT_B17_enable = SB_T4_WEST_SB_OUT_B17_enable_value_O[0];
assign SB_T4_WEST_SB_OUT_B17_valid_out = RMUX_T4_WEST_B17_valid_out;
assign read_config_data = mux_aoi_6_32_inst0_O;
endmodule

module SB_ID0_5TRACKS_B17_MemCore (
    input [0:0] MEM_input_width_17_num_0_enable,
    input [31:0] MEM_input_width_17_num_0_out_sel,
    input MEM_input_width_17_num_0_ready,
    input [0:0] MEM_input_width_17_num_1_enable,
    input [31:0] MEM_input_width_17_num_1_out_sel,
    input MEM_input_width_17_num_1_ready,
    input [0:0] MEM_input_width_17_num_2_enable,
    input [31:0] MEM_input_width_17_num_2_out_sel,
    input MEM_input_width_17_num_2_ready,
    input [0:0] MEM_input_width_17_num_3_enable,
    input [31:0] MEM_input_width_17_num_3_out_sel,
    input MEM_input_width_17_num_3_ready,
    input [16:0] MEM_output_width_17_num_0,
    output MEM_output_width_17_num_0_ready_out,
    input MEM_output_width_17_num_0_valid,
    input [16:0] MEM_output_width_17_num_1,
    output MEM_output_width_17_num_1_ready_out,
    input MEM_output_width_17_num_1_valid,
    input [16:0] MEM_output_width_17_num_2,
    output MEM_output_width_17_num_2_ready_out,
    input MEM_output_width_17_num_2_valid,
    input [16:0] SB_T0_EAST_SB_IN_B17,
    output SB_T0_EAST_SB_IN_B17_enable,
    output SB_T0_EAST_SB_IN_B17_ready_out,
    input SB_T0_EAST_SB_IN_B17_valid_in,
    output [16:0] SB_T0_EAST_SB_OUT_B17,
    output SB_T0_EAST_SB_OUT_B17_enable,
    input SB_T0_EAST_SB_OUT_B17_ready_in,
    output SB_T0_EAST_SB_OUT_B17_valid_out,
    input [16:0] SB_T0_NORTH_SB_IN_B17,
    output SB_T0_NORTH_SB_IN_B17_enable,
    output SB_T0_NORTH_SB_IN_B17_ready_out,
    input SB_T0_NORTH_SB_IN_B17_valid_in,
    output [16:0] SB_T0_NORTH_SB_OUT_B17,
    output SB_T0_NORTH_SB_OUT_B17_enable,
    input SB_T0_NORTH_SB_OUT_B17_ready_in,
    output SB_T0_NORTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T0_SOUTH_SB_IN_B17,
    output SB_T0_SOUTH_SB_IN_B17_enable,
    output SB_T0_SOUTH_SB_IN_B17_ready_out,
    input SB_T0_SOUTH_SB_IN_B17_valid_in,
    output [16:0] SB_T0_SOUTH_SB_OUT_B17,
    output SB_T0_SOUTH_SB_OUT_B17_enable,
    input SB_T0_SOUTH_SB_OUT_B17_ready_in,
    output SB_T0_SOUTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T0_WEST_SB_IN_B17,
    output SB_T0_WEST_SB_IN_B17_enable,
    output SB_T0_WEST_SB_IN_B17_ready_out,
    input SB_T0_WEST_SB_IN_B17_valid_in,
    output [16:0] SB_T0_WEST_SB_OUT_B17,
    output SB_T0_WEST_SB_OUT_B17_enable,
    input SB_T0_WEST_SB_OUT_B17_ready_in,
    output SB_T0_WEST_SB_OUT_B17_valid_out,
    input [16:0] SB_T1_EAST_SB_IN_B17,
    output SB_T1_EAST_SB_IN_B17_enable,
    output SB_T1_EAST_SB_IN_B17_ready_out,
    input SB_T1_EAST_SB_IN_B17_valid_in,
    output [16:0] SB_T1_EAST_SB_OUT_B17,
    output SB_T1_EAST_SB_OUT_B17_enable,
    input SB_T1_EAST_SB_OUT_B17_ready_in,
    output SB_T1_EAST_SB_OUT_B17_valid_out,
    input [16:0] SB_T1_NORTH_SB_IN_B17,
    output SB_T1_NORTH_SB_IN_B17_enable,
    output SB_T1_NORTH_SB_IN_B17_ready_out,
    input SB_T1_NORTH_SB_IN_B17_valid_in,
    output [16:0] SB_T1_NORTH_SB_OUT_B17,
    output SB_T1_NORTH_SB_OUT_B17_enable,
    input SB_T1_NORTH_SB_OUT_B17_ready_in,
    output SB_T1_NORTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T1_SOUTH_SB_IN_B17,
    output SB_T1_SOUTH_SB_IN_B17_enable,
    output SB_T1_SOUTH_SB_IN_B17_ready_out,
    input SB_T1_SOUTH_SB_IN_B17_valid_in,
    output [16:0] SB_T1_SOUTH_SB_OUT_B17,
    output SB_T1_SOUTH_SB_OUT_B17_enable,
    input SB_T1_SOUTH_SB_OUT_B17_ready_in,
    output SB_T1_SOUTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T1_WEST_SB_IN_B17,
    output SB_T1_WEST_SB_IN_B17_enable,
    output SB_T1_WEST_SB_IN_B17_ready_out,
    input SB_T1_WEST_SB_IN_B17_valid_in,
    output [16:0] SB_T1_WEST_SB_OUT_B17,
    output SB_T1_WEST_SB_OUT_B17_enable,
    input SB_T1_WEST_SB_OUT_B17_ready_in,
    output SB_T1_WEST_SB_OUT_B17_valid_out,
    input [16:0] SB_T2_EAST_SB_IN_B17,
    output SB_T2_EAST_SB_IN_B17_enable,
    output SB_T2_EAST_SB_IN_B17_ready_out,
    input SB_T2_EAST_SB_IN_B17_valid_in,
    output [16:0] SB_T2_EAST_SB_OUT_B17,
    output SB_T2_EAST_SB_OUT_B17_enable,
    input SB_T2_EAST_SB_OUT_B17_ready_in,
    output SB_T2_EAST_SB_OUT_B17_valid_out,
    input [16:0] SB_T2_NORTH_SB_IN_B17,
    output SB_T2_NORTH_SB_IN_B17_enable,
    output SB_T2_NORTH_SB_IN_B17_ready_out,
    input SB_T2_NORTH_SB_IN_B17_valid_in,
    output [16:0] SB_T2_NORTH_SB_OUT_B17,
    output SB_T2_NORTH_SB_OUT_B17_enable,
    input SB_T2_NORTH_SB_OUT_B17_ready_in,
    output SB_T2_NORTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T2_SOUTH_SB_IN_B17,
    output SB_T2_SOUTH_SB_IN_B17_enable,
    output SB_T2_SOUTH_SB_IN_B17_ready_out,
    input SB_T2_SOUTH_SB_IN_B17_valid_in,
    output [16:0] SB_T2_SOUTH_SB_OUT_B17,
    output SB_T2_SOUTH_SB_OUT_B17_enable,
    input SB_T2_SOUTH_SB_OUT_B17_ready_in,
    output SB_T2_SOUTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T2_WEST_SB_IN_B17,
    output SB_T2_WEST_SB_IN_B17_enable,
    output SB_T2_WEST_SB_IN_B17_ready_out,
    input SB_T2_WEST_SB_IN_B17_valid_in,
    output [16:0] SB_T2_WEST_SB_OUT_B17,
    output SB_T2_WEST_SB_OUT_B17_enable,
    input SB_T2_WEST_SB_OUT_B17_ready_in,
    output SB_T2_WEST_SB_OUT_B17_valid_out,
    input [16:0] SB_T3_EAST_SB_IN_B17,
    output SB_T3_EAST_SB_IN_B17_enable,
    output SB_T3_EAST_SB_IN_B17_ready_out,
    input SB_T3_EAST_SB_IN_B17_valid_in,
    output [16:0] SB_T3_EAST_SB_OUT_B17,
    output SB_T3_EAST_SB_OUT_B17_enable,
    input SB_T3_EAST_SB_OUT_B17_ready_in,
    output SB_T3_EAST_SB_OUT_B17_valid_out,
    input [16:0] SB_T3_NORTH_SB_IN_B17,
    output SB_T3_NORTH_SB_IN_B17_enable,
    output SB_T3_NORTH_SB_IN_B17_ready_out,
    input SB_T3_NORTH_SB_IN_B17_valid_in,
    output [16:0] SB_T3_NORTH_SB_OUT_B17,
    output SB_T3_NORTH_SB_OUT_B17_enable,
    input SB_T3_NORTH_SB_OUT_B17_ready_in,
    output SB_T3_NORTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T3_SOUTH_SB_IN_B17,
    output SB_T3_SOUTH_SB_IN_B17_enable,
    output SB_T3_SOUTH_SB_IN_B17_ready_out,
    input SB_T3_SOUTH_SB_IN_B17_valid_in,
    output [16:0] SB_T3_SOUTH_SB_OUT_B17,
    output SB_T3_SOUTH_SB_OUT_B17_enable,
    input SB_T3_SOUTH_SB_OUT_B17_ready_in,
    output SB_T3_SOUTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T3_WEST_SB_IN_B17,
    output SB_T3_WEST_SB_IN_B17_enable,
    output SB_T3_WEST_SB_IN_B17_ready_out,
    input SB_T3_WEST_SB_IN_B17_valid_in,
    output [16:0] SB_T3_WEST_SB_OUT_B17,
    output SB_T3_WEST_SB_OUT_B17_enable,
    input SB_T3_WEST_SB_OUT_B17_ready_in,
    output SB_T3_WEST_SB_OUT_B17_valid_out,
    input [16:0] SB_T4_EAST_SB_IN_B17,
    output SB_T4_EAST_SB_IN_B17_enable,
    output SB_T4_EAST_SB_IN_B17_ready_out,
    input SB_T4_EAST_SB_IN_B17_valid_in,
    output [16:0] SB_T4_EAST_SB_OUT_B17,
    output SB_T4_EAST_SB_OUT_B17_enable,
    input SB_T4_EAST_SB_OUT_B17_ready_in,
    output SB_T4_EAST_SB_OUT_B17_valid_out,
    input [16:0] SB_T4_NORTH_SB_IN_B17,
    output SB_T4_NORTH_SB_IN_B17_enable,
    output SB_T4_NORTH_SB_IN_B17_ready_out,
    input SB_T4_NORTH_SB_IN_B17_valid_in,
    output [16:0] SB_T4_NORTH_SB_OUT_B17,
    output SB_T4_NORTH_SB_OUT_B17_enable,
    input SB_T4_NORTH_SB_OUT_B17_ready_in,
    output SB_T4_NORTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T4_SOUTH_SB_IN_B17,
    output SB_T4_SOUTH_SB_IN_B17_enable,
    output SB_T4_SOUTH_SB_IN_B17_ready_out,
    input SB_T4_SOUTH_SB_IN_B17_valid_in,
    output [16:0] SB_T4_SOUTH_SB_OUT_B17,
    output SB_T4_SOUTH_SB_OUT_B17_enable,
    input SB_T4_SOUTH_SB_OUT_B17_ready_in,
    output SB_T4_SOUTH_SB_OUT_B17_valid_out,
    input [16:0] SB_T4_WEST_SB_IN_B17,
    output SB_T4_WEST_SB_IN_B17_enable,
    output SB_T4_WEST_SB_IN_B17_ready_out,
    input SB_T4_WEST_SB_IN_B17_valid_in,
    output [16:0] SB_T4_WEST_SB_OUT_B17,
    output SB_T4_WEST_SB_OUT_B17_enable,
    input SB_T4_WEST_SB_OUT_B17_ready_in,
    output SB_T4_WEST_SB_OUT_B17_valid_out,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset,
    input [0:0] stall
);
wire [0:0] CB_MEM_output_width_17_num_0_fan_in_O;
wire [0:0] CB_MEM_output_width_17_num_1_fan_in_O;
wire [0:0] CB_MEM_output_width_17_num_2_fan_in_O;
wire [0:0] Invert1_inst0_out;
wire [16:0] MUX_SB_T0_EAST_SB_OUT_B17_O;
wire MUX_SB_T0_EAST_SB_OUT_B17_ready_out;
wire MUX_SB_T0_EAST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T0_EAST_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T0_NORTH_SB_OUT_B17_O;
wire MUX_SB_T0_NORTH_SB_OUT_B17_ready_out;
wire MUX_SB_T0_NORTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T0_NORTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T0_SOUTH_SB_OUT_B17_O;
wire MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out;
wire MUX_SB_T0_SOUTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T0_WEST_SB_OUT_B17_O;
wire MUX_SB_T0_WEST_SB_OUT_B17_ready_out;
wire MUX_SB_T0_WEST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T0_WEST_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T1_EAST_SB_OUT_B17_O;
wire MUX_SB_T1_EAST_SB_OUT_B17_ready_out;
wire MUX_SB_T1_EAST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T1_EAST_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T1_NORTH_SB_OUT_B17_O;
wire MUX_SB_T1_NORTH_SB_OUT_B17_ready_out;
wire MUX_SB_T1_NORTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T1_NORTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T1_SOUTH_SB_OUT_B17_O;
wire MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out;
wire MUX_SB_T1_SOUTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T1_WEST_SB_OUT_B17_O;
wire MUX_SB_T1_WEST_SB_OUT_B17_ready_out;
wire MUX_SB_T1_WEST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T1_WEST_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T2_EAST_SB_OUT_B17_O;
wire MUX_SB_T2_EAST_SB_OUT_B17_ready_out;
wire MUX_SB_T2_EAST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T2_EAST_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T2_NORTH_SB_OUT_B17_O;
wire MUX_SB_T2_NORTH_SB_OUT_B17_ready_out;
wire MUX_SB_T2_NORTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T2_NORTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T2_SOUTH_SB_OUT_B17_O;
wire MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out;
wire MUX_SB_T2_SOUTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T2_WEST_SB_OUT_B17_O;
wire MUX_SB_T2_WEST_SB_OUT_B17_ready_out;
wire MUX_SB_T2_WEST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T2_WEST_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T3_EAST_SB_OUT_B17_O;
wire MUX_SB_T3_EAST_SB_OUT_B17_ready_out;
wire MUX_SB_T3_EAST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T3_EAST_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T3_NORTH_SB_OUT_B17_O;
wire MUX_SB_T3_NORTH_SB_OUT_B17_ready_out;
wire MUX_SB_T3_NORTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T3_NORTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T3_SOUTH_SB_OUT_B17_O;
wire MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out;
wire MUX_SB_T3_SOUTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T3_WEST_SB_OUT_B17_O;
wire MUX_SB_T3_WEST_SB_OUT_B17_ready_out;
wire MUX_SB_T3_WEST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T3_WEST_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T4_EAST_SB_OUT_B17_O;
wire MUX_SB_T4_EAST_SB_OUT_B17_ready_out;
wire MUX_SB_T4_EAST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T4_EAST_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T4_NORTH_SB_OUT_B17_O;
wire MUX_SB_T4_NORTH_SB_OUT_B17_ready_out;
wire MUX_SB_T4_NORTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T4_NORTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T4_SOUTH_SB_OUT_B17_O;
wire MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out;
wire MUX_SB_T4_SOUTH_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel;
wire [16:0] MUX_SB_T4_WEST_SB_OUT_B17_O;
wire MUX_SB_T4_WEST_SB_OUT_B17_ready_out;
wire MUX_SB_T4_WEST_SB_OUT_B17_valid_out;
wire [7:0] MUX_SB_T4_WEST_SB_OUT_B17_out_sel;
wire [0:0] REG_T0_EAST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T0_EAST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T0_EAST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T0_EAST_B17_end_value_O;
wire [0:0] REG_T0_EAST_B17_fifo_value_O;
wire [0:0] REG_T0_EAST_B17_start_value_O;
wire [0:0] REG_T0_NORTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T0_NORTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T0_NORTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T0_NORTH_B17_end_value_O;
wire [0:0] REG_T0_NORTH_B17_fifo_value_O;
wire [0:0] REG_T0_NORTH_B17_start_value_O;
wire [0:0] REG_T0_SOUTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T0_SOUTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T0_SOUTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T0_SOUTH_B17_end_value_O;
wire [0:0] REG_T0_SOUTH_B17_fifo_value_O;
wire [0:0] REG_T0_SOUTH_B17_start_value_O;
wire [0:0] REG_T0_WEST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T0_WEST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T0_WEST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T0_WEST_B17_end_value_O;
wire [0:0] REG_T0_WEST_B17_fifo_value_O;
wire [0:0] REG_T0_WEST_B17_start_value_O;
wire [0:0] REG_T1_EAST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T1_EAST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T1_EAST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T1_EAST_B17_end_value_O;
wire [0:0] REG_T1_EAST_B17_fifo_value_O;
wire [0:0] REG_T1_EAST_B17_start_value_O;
wire [0:0] REG_T1_NORTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T1_NORTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T1_NORTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T1_NORTH_B17_end_value_O;
wire [0:0] REG_T1_NORTH_B17_fifo_value_O;
wire [0:0] REG_T1_NORTH_B17_start_value_O;
wire [0:0] REG_T1_SOUTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T1_SOUTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T1_SOUTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T1_SOUTH_B17_end_value_O;
wire [0:0] REG_T1_SOUTH_B17_fifo_value_O;
wire [0:0] REG_T1_SOUTH_B17_start_value_O;
wire [0:0] REG_T1_WEST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T1_WEST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T1_WEST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T1_WEST_B17_end_value_O;
wire [0:0] REG_T1_WEST_B17_fifo_value_O;
wire [0:0] REG_T1_WEST_B17_start_value_O;
wire [0:0] REG_T2_EAST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T2_EAST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T2_EAST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T2_EAST_B17_end_value_O;
wire [0:0] REG_T2_EAST_B17_fifo_value_O;
wire [0:0] REG_T2_EAST_B17_start_value_O;
wire [0:0] REG_T2_NORTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T2_NORTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T2_NORTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T2_NORTH_B17_end_value_O;
wire [0:0] REG_T2_NORTH_B17_fifo_value_O;
wire [0:0] REG_T2_NORTH_B17_start_value_O;
wire [0:0] REG_T2_SOUTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T2_SOUTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T2_SOUTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T2_SOUTH_B17_end_value_O;
wire [0:0] REG_T2_SOUTH_B17_fifo_value_O;
wire [0:0] REG_T2_SOUTH_B17_start_value_O;
wire [0:0] REG_T2_WEST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T2_WEST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T2_WEST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T2_WEST_B17_end_value_O;
wire [0:0] REG_T2_WEST_B17_fifo_value_O;
wire [0:0] REG_T2_WEST_B17_start_value_O;
wire [0:0] REG_T3_EAST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T3_EAST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T3_EAST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T3_EAST_B17_end_value_O;
wire [0:0] REG_T3_EAST_B17_fifo_value_O;
wire [0:0] REG_T3_EAST_B17_start_value_O;
wire [0:0] REG_T3_NORTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T3_NORTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T3_NORTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T3_NORTH_B17_end_value_O;
wire [0:0] REG_T3_NORTH_B17_fifo_value_O;
wire [0:0] REG_T3_NORTH_B17_start_value_O;
wire [0:0] REG_T3_SOUTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T3_SOUTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T3_SOUTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T3_SOUTH_B17_end_value_O;
wire [0:0] REG_T3_SOUTH_B17_fifo_value_O;
wire [0:0] REG_T3_SOUTH_B17_start_value_O;
wire [0:0] REG_T3_WEST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T3_WEST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T3_WEST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T3_WEST_B17_end_value_O;
wire [0:0] REG_T3_WEST_B17_fifo_value_O;
wire [0:0] REG_T3_WEST_B17_start_value_O;
wire [0:0] REG_T4_EAST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T4_EAST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T4_EAST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T4_EAST_B17_end_value_O;
wire [0:0] REG_T4_EAST_B17_fifo_value_O;
wire [0:0] REG_T4_EAST_B17_start_value_O;
wire [0:0] REG_T4_NORTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T4_NORTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T4_NORTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T4_NORTH_B17_end_value_O;
wire [0:0] REG_T4_NORTH_B17_fifo_value_O;
wire [0:0] REG_T4_NORTH_B17_start_value_O;
wire [0:0] REG_T4_SOUTH_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T4_SOUTH_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T4_SOUTH_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T4_SOUTH_B17_end_value_O;
wire [0:0] REG_T4_SOUTH_B17_fifo_value_O;
wire [0:0] REG_T4_SOUTH_B17_start_value_O;
wire [0:0] REG_T4_WEST_B17$SplitFifo_17_inst0_ready0;
wire [0:0] REG_T4_WEST_B17$SplitFifo_17_inst0_valid1;
wire [16:0] REG_T4_WEST_B17$SplitFifo_17_inst0_data_out;
wire [0:0] REG_T4_WEST_B17_end_value_O;
wire [0:0] REG_T4_WEST_B17_fifo_value_O;
wire [0:0] REG_T4_WEST_B17_start_value_O;
wire [16:0] RMUX_T0_EAST_B17_O;
wire RMUX_T0_EAST_B17_ready_out;
wire RMUX_T0_EAST_B17_valid_out;
wire [1:0] RMUX_T0_EAST_B17_out_sel;
wire [0:0] RMUX_T0_EAST_B17_sel_value_O;
wire [16:0] RMUX_T0_NORTH_B17_O;
wire RMUX_T0_NORTH_B17_ready_out;
wire RMUX_T0_NORTH_B17_valid_out;
wire [1:0] RMUX_T0_NORTH_B17_out_sel;
wire [0:0] RMUX_T0_NORTH_B17_sel_value_O;
wire [16:0] RMUX_T0_SOUTH_B17_O;
wire RMUX_T0_SOUTH_B17_ready_out;
wire RMUX_T0_SOUTH_B17_valid_out;
wire [1:0] RMUX_T0_SOUTH_B17_out_sel;
wire [0:0] RMUX_T0_SOUTH_B17_sel_value_O;
wire [16:0] RMUX_T0_WEST_B17_O;
wire RMUX_T0_WEST_B17_ready_out;
wire RMUX_T0_WEST_B17_valid_out;
wire [1:0] RMUX_T0_WEST_B17_out_sel;
wire [0:0] RMUX_T0_WEST_B17_sel_value_O;
wire [16:0] RMUX_T1_EAST_B17_O;
wire RMUX_T1_EAST_B17_ready_out;
wire RMUX_T1_EAST_B17_valid_out;
wire [1:0] RMUX_T1_EAST_B17_out_sel;
wire [0:0] RMUX_T1_EAST_B17_sel_value_O;
wire [16:0] RMUX_T1_NORTH_B17_O;
wire RMUX_T1_NORTH_B17_ready_out;
wire RMUX_T1_NORTH_B17_valid_out;
wire [1:0] RMUX_T1_NORTH_B17_out_sel;
wire [0:0] RMUX_T1_NORTH_B17_sel_value_O;
wire [16:0] RMUX_T1_SOUTH_B17_O;
wire RMUX_T1_SOUTH_B17_ready_out;
wire RMUX_T1_SOUTH_B17_valid_out;
wire [1:0] RMUX_T1_SOUTH_B17_out_sel;
wire [0:0] RMUX_T1_SOUTH_B17_sel_value_O;
wire [16:0] RMUX_T1_WEST_B17_O;
wire RMUX_T1_WEST_B17_ready_out;
wire RMUX_T1_WEST_B17_valid_out;
wire [1:0] RMUX_T1_WEST_B17_out_sel;
wire [0:0] RMUX_T1_WEST_B17_sel_value_O;
wire [16:0] RMUX_T2_EAST_B17_O;
wire RMUX_T2_EAST_B17_ready_out;
wire RMUX_T2_EAST_B17_valid_out;
wire [1:0] RMUX_T2_EAST_B17_out_sel;
wire [0:0] RMUX_T2_EAST_B17_sel_value_O;
wire [16:0] RMUX_T2_NORTH_B17_O;
wire RMUX_T2_NORTH_B17_ready_out;
wire RMUX_T2_NORTH_B17_valid_out;
wire [1:0] RMUX_T2_NORTH_B17_out_sel;
wire [0:0] RMUX_T2_NORTH_B17_sel_value_O;
wire [16:0] RMUX_T2_SOUTH_B17_O;
wire RMUX_T2_SOUTH_B17_ready_out;
wire RMUX_T2_SOUTH_B17_valid_out;
wire [1:0] RMUX_T2_SOUTH_B17_out_sel;
wire [0:0] RMUX_T2_SOUTH_B17_sel_value_O;
wire [16:0] RMUX_T2_WEST_B17_O;
wire RMUX_T2_WEST_B17_ready_out;
wire RMUX_T2_WEST_B17_valid_out;
wire [1:0] RMUX_T2_WEST_B17_out_sel;
wire [0:0] RMUX_T2_WEST_B17_sel_value_O;
wire [16:0] RMUX_T3_EAST_B17_O;
wire RMUX_T3_EAST_B17_ready_out;
wire RMUX_T3_EAST_B17_valid_out;
wire [1:0] RMUX_T3_EAST_B17_out_sel;
wire [0:0] RMUX_T3_EAST_B17_sel_value_O;
wire [16:0] RMUX_T3_NORTH_B17_O;
wire RMUX_T3_NORTH_B17_ready_out;
wire RMUX_T3_NORTH_B17_valid_out;
wire [1:0] RMUX_T3_NORTH_B17_out_sel;
wire [0:0] RMUX_T3_NORTH_B17_sel_value_O;
wire [16:0] RMUX_T3_SOUTH_B17_O;
wire RMUX_T3_SOUTH_B17_ready_out;
wire RMUX_T3_SOUTH_B17_valid_out;
wire [1:0] RMUX_T3_SOUTH_B17_out_sel;
wire [0:0] RMUX_T3_SOUTH_B17_sel_value_O;
wire [16:0] RMUX_T3_WEST_B17_O;
wire RMUX_T3_WEST_B17_ready_out;
wire RMUX_T3_WEST_B17_valid_out;
wire [1:0] RMUX_T3_WEST_B17_out_sel;
wire [0:0] RMUX_T3_WEST_B17_sel_value_O;
wire [16:0] RMUX_T4_EAST_B17_O;
wire RMUX_T4_EAST_B17_ready_out;
wire RMUX_T4_EAST_B17_valid_out;
wire [1:0] RMUX_T4_EAST_B17_out_sel;
wire [0:0] RMUX_T4_EAST_B17_sel_value_O;
wire [16:0] RMUX_T4_NORTH_B17_O;
wire RMUX_T4_NORTH_B17_ready_out;
wire RMUX_T4_NORTH_B17_valid_out;
wire [1:0] RMUX_T4_NORTH_B17_out_sel;
wire [0:0] RMUX_T4_NORTH_B17_sel_value_O;
wire [16:0] RMUX_T4_SOUTH_B17_O;
wire RMUX_T4_SOUTH_B17_ready_out;
wire RMUX_T4_SOUTH_B17_valid_out;
wire [1:0] RMUX_T4_SOUTH_B17_out_sel;
wire [0:0] RMUX_T4_SOUTH_B17_sel_value_O;
wire [16:0] RMUX_T4_WEST_B17_O;
wire RMUX_T4_WEST_B17_ready_out;
wire RMUX_T4_WEST_B17_valid_out;
wire [1:0] RMUX_T4_WEST_B17_out_sel;
wire [0:0] RMUX_T4_WEST_B17_sel_value_O;
wire [0:0] SB_T0_EAST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T0_EAST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T0_EAST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T0_EAST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T0_EAST_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T0_NORTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T0_NORTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T0_NORTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T0_NORTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T0_NORTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T0_SOUTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T0_SOUTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T0_SOUTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T0_SOUTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T0_SOUTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T0_WEST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T0_WEST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T0_WEST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T0_WEST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T0_WEST_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T1_EAST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T1_EAST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T1_EAST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T1_EAST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T1_EAST_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T1_NORTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T1_NORTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T1_NORTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T1_NORTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T1_NORTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T1_SOUTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T1_SOUTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T1_SOUTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T1_SOUTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T1_SOUTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T1_WEST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T1_WEST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T1_WEST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T1_WEST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T1_WEST_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T2_EAST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T2_EAST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T2_EAST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T2_EAST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T2_EAST_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T2_NORTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T2_NORTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T2_NORTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T2_NORTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T2_NORTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T2_SOUTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T2_SOUTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T2_SOUTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T2_SOUTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T2_SOUTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T2_WEST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T2_WEST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T2_WEST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T2_WEST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T2_WEST_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T3_EAST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T3_EAST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T3_EAST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T3_EAST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T3_EAST_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T3_NORTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T3_NORTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T3_NORTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T3_NORTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T3_NORTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T3_SOUTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T3_SOUTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T3_SOUTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T3_SOUTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T3_SOUTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T3_WEST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T3_WEST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T3_WEST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T3_WEST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T3_WEST_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T4_EAST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T4_EAST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T4_EAST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T4_EAST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T4_EAST_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T4_NORTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T4_NORTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T4_NORTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T4_NORTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T4_NORTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T4_SOUTH_SB_IN_B17_enable_value_O;
wire [0:0] SB_T4_SOUTH_SB_IN_B17_fan_in_O;
wire [0:0] SB_T4_SOUTH_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T4_SOUTH_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T4_SOUTH_SB_OUT_B17_sel_value_O;
wire [0:0] SB_T4_WEST_SB_IN_B17_enable_value_O;
wire [0:0] SB_T4_WEST_SB_IN_B17_fan_in_O;
wire [0:0] SB_T4_WEST_SB_OUT_B17_FANOUT_O;
wire [0:0] SB_T4_WEST_SB_OUT_B17_enable_value_O;
wire [2:0] SB_T4_WEST_SB_OUT_B17_sel_value_O;
wire [16:0] WIRE_SB_T0_EAST_SB_IN_B17_O;
wire WIRE_SB_T0_EAST_SB_IN_B17_ready_out;
wire WIRE_SB_T0_EAST_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T0_NORTH_SB_IN_B17_O;
wire WIRE_SB_T0_NORTH_SB_IN_B17_ready_out;
wire WIRE_SB_T0_NORTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T0_SOUTH_SB_IN_B17_O;
wire WIRE_SB_T0_SOUTH_SB_IN_B17_ready_out;
wire WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T0_WEST_SB_IN_B17_O;
wire WIRE_SB_T0_WEST_SB_IN_B17_ready_out;
wire WIRE_SB_T0_WEST_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T1_EAST_SB_IN_B17_O;
wire WIRE_SB_T1_EAST_SB_IN_B17_ready_out;
wire WIRE_SB_T1_EAST_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T1_NORTH_SB_IN_B17_O;
wire WIRE_SB_T1_NORTH_SB_IN_B17_ready_out;
wire WIRE_SB_T1_NORTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T1_SOUTH_SB_IN_B17_O;
wire WIRE_SB_T1_SOUTH_SB_IN_B17_ready_out;
wire WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T1_WEST_SB_IN_B17_O;
wire WIRE_SB_T1_WEST_SB_IN_B17_ready_out;
wire WIRE_SB_T1_WEST_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T2_EAST_SB_IN_B17_O;
wire WIRE_SB_T2_EAST_SB_IN_B17_ready_out;
wire WIRE_SB_T2_EAST_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T2_NORTH_SB_IN_B17_O;
wire WIRE_SB_T2_NORTH_SB_IN_B17_ready_out;
wire WIRE_SB_T2_NORTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T2_SOUTH_SB_IN_B17_O;
wire WIRE_SB_T2_SOUTH_SB_IN_B17_ready_out;
wire WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T2_WEST_SB_IN_B17_O;
wire WIRE_SB_T2_WEST_SB_IN_B17_ready_out;
wire WIRE_SB_T2_WEST_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T3_EAST_SB_IN_B17_O;
wire WIRE_SB_T3_EAST_SB_IN_B17_ready_out;
wire WIRE_SB_T3_EAST_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T3_NORTH_SB_IN_B17_O;
wire WIRE_SB_T3_NORTH_SB_IN_B17_ready_out;
wire WIRE_SB_T3_NORTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T3_SOUTH_SB_IN_B17_O;
wire WIRE_SB_T3_SOUTH_SB_IN_B17_ready_out;
wire WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T3_WEST_SB_IN_B17_O;
wire WIRE_SB_T3_WEST_SB_IN_B17_ready_out;
wire WIRE_SB_T3_WEST_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T4_EAST_SB_IN_B17_O;
wire WIRE_SB_T4_EAST_SB_IN_B17_ready_out;
wire WIRE_SB_T4_EAST_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T4_NORTH_SB_IN_B17_O;
wire WIRE_SB_T4_NORTH_SB_IN_B17_ready_out;
wire WIRE_SB_T4_NORTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T4_SOUTH_SB_IN_B17_O;
wire WIRE_SB_T4_SOUTH_SB_IN_B17_ready_out;
wire WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out;
wire [16:0] WIRE_SB_T4_WEST_SB_IN_B17_O;
wire WIRE_SB_T4_WEST_SB_IN_B17_ready_out;
wire WIRE_SB_T4_WEST_SB_IN_B17_valid_out;
wire ZextWrapper_23_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_23_32_inst0$self_O_in;
wire ZextWrapper_30_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_30_32_inst0$self_O_in;
wire ZextWrapper_31_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_31_32_inst0$self_O_in;
wire [0:0] and1_inst0_out;
wire [0:0] and1_inst1_out;
wire [0:0] and1_inst10_out;
wire [0:0] and1_inst11_out;
wire [0:0] and1_inst12_out;
wire [0:0] and1_inst13_out;
wire [0:0] and1_inst14_out;
wire [0:0] and1_inst15_out;
wire [0:0] and1_inst16_out;
wire [0:0] and1_inst17_out;
wire [0:0] and1_inst18_out;
wire [0:0] and1_inst19_out;
wire [0:0] and1_inst2_out;
wire [0:0] and1_inst3_out;
wire [0:0] and1_inst4_out;
wire [0:0] and1_inst5_out;
wire [0:0] and1_inst6_out;
wire [0:0] and1_inst7_out;
wire [0:0] and1_inst8_out;
wire [0:0] and1_inst9_out;
wire [31:0] config_reg_0_O;
wire [31:0] config_reg_1_O;
wire [31:0] config_reg_2_O;
wire [30:0] config_reg_3_O;
wire [29:0] config_reg_4_O;
wire [22:0] config_reg_5_O;
wire [0:0] const_1_1_out;
wire coreir_eq_1_inst0_out;
wire coreir_eq_1_inst1_out;
wire coreir_eq_1_inst10_out;
wire coreir_eq_1_inst11_out;
wire coreir_eq_1_inst12_out;
wire coreir_eq_1_inst13_out;
wire coreir_eq_1_inst14_out;
wire coreir_eq_1_inst15_out;
wire coreir_eq_1_inst16_out;
wire coreir_eq_1_inst17_out;
wire coreir_eq_1_inst18_out;
wire coreir_eq_1_inst19_out;
wire coreir_eq_1_inst2_out;
wire coreir_eq_1_inst3_out;
wire coreir_eq_1_inst4_out;
wire coreir_eq_1_inst5_out;
wire coreir_eq_1_inst6_out;
wire coreir_eq_1_inst7_out;
wire coreir_eq_1_inst8_out;
wire coreir_eq_1_inst9_out;
wire [31:0] mux_aoi_6_32_inst0_O;
wire [7:0] mux_aoi_6_32_inst0_out_sel;
wire [7:0] self_config_config_addr_out;
FanoutHash_E70AF988E4250F5 CB_MEM_output_width_17_num_0_fan_in (
    .S13(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
    .E13(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
    .S6(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
    .E2(SB_T0_EAST_SB_OUT_B17_enable_value_O),
    .E12(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
    .E7(SB_T1_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
    .E18(SB_T4_EAST_SB_OUT_B17_enable_value_O),
    .I3(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
    .E19(SB_T4_WEST_SB_OUT_B17_enable_value_O),
    .I14(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
    .S14(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
    .I9(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
    .S12(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
    .S17(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
    .I13(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
    .S9(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
    .E10(SB_T2_EAST_SB_OUT_B17_enable_value_O),
    .E15(SB_T3_WEST_SB_OUT_B17_enable_value_O),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
    .E5(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
    .S10(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
    .E8(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
    .I11(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
    .I6(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
    .S15(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
    .I7(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
    .E14(SB_T3_EAST_SB_OUT_B17_enable_value_O),
    .I2(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
    .E11(SB_T2_WEST_SB_OUT_B17_enable_value_O),
    .S3(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
    .S8(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
    .I10(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
    .S16(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
    .E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
    .E16(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
    .E3(SB_T0_WEST_SB_OUT_B17_enable_value_O),
    .S18(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
    .S19(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
    .S2(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
    .S4(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
    .E9(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
    .I16(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
    .I12(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
    .S11(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
    .I17(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
    .I19(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
    .I18(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
    .S7(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
    .E4(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
    .E17(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
    .S5(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
    .I1(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
    .I5(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
    .E6(SB_T1_EAST_SB_OUT_B17_enable_value_O),
    .I4(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
    .I8(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
    .O(CB_MEM_output_width_17_num_0_fan_in_O),
    .E1(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
    .I15(MUX_SB_T3_WEST_SB_OUT_B17_ready_out)
);
FanoutHash_82899D6851EDC11 CB_MEM_output_width_17_num_1_fan_in (
    .S13(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
    .E13(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
    .S6(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
    .E2(SB_T0_EAST_SB_OUT_B17_enable_value_O),
    .E12(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
    .E7(SB_T1_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
    .E18(SB_T4_EAST_SB_OUT_B17_enable_value_O),
    .I3(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
    .E19(SB_T4_WEST_SB_OUT_B17_enable_value_O),
    .I14(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
    .S14(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
    .I9(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
    .S12(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
    .S17(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
    .I13(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
    .S9(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
    .E10(SB_T2_EAST_SB_OUT_B17_enable_value_O),
    .E15(SB_T3_WEST_SB_OUT_B17_enable_value_O),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
    .E5(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
    .S10(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
    .E8(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
    .I11(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
    .I6(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
    .S15(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
    .I7(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
    .E14(SB_T3_EAST_SB_OUT_B17_enable_value_O),
    .I2(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
    .E11(SB_T2_WEST_SB_OUT_B17_enable_value_O),
    .S3(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
    .S8(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
    .I10(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
    .S16(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
    .E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
    .E16(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
    .E3(SB_T0_WEST_SB_OUT_B17_enable_value_O),
    .S18(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
    .S19(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
    .S2(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
    .S4(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
    .E9(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
    .I16(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
    .I12(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
    .S11(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
    .I17(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
    .I19(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
    .I18(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
    .S7(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
    .E4(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
    .E17(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
    .S5(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
    .I1(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
    .I5(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
    .E6(SB_T1_EAST_SB_OUT_B17_enable_value_O),
    .I4(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
    .I8(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
    .O(CB_MEM_output_width_17_num_1_fan_in_O),
    .E1(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
    .I15(MUX_SB_T3_WEST_SB_OUT_B17_ready_out)
);
FanoutHash_CE1AA874B742213 CB_MEM_output_width_17_num_2_fan_in (
    .S13(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
    .E13(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
    .S6(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
    .E2(SB_T0_EAST_SB_OUT_B17_enable_value_O),
    .E12(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
    .E7(SB_T1_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
    .E18(SB_T4_EAST_SB_OUT_B17_enable_value_O),
    .I3(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
    .E19(SB_T4_WEST_SB_OUT_B17_enable_value_O),
    .I14(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
    .S14(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
    .I9(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
    .S12(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
    .S17(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
    .I13(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
    .S9(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
    .E10(SB_T2_EAST_SB_OUT_B17_enable_value_O),
    .E15(SB_T3_WEST_SB_OUT_B17_enable_value_O),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
    .E5(SB_T1_SOUTH_SB_OUT_B17_enable_value_O),
    .S10(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
    .E8(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
    .I11(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
    .I6(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
    .S15(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
    .I7(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
    .E14(SB_T3_EAST_SB_OUT_B17_enable_value_O),
    .I2(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
    .E11(SB_T2_WEST_SB_OUT_B17_enable_value_O),
    .S3(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
    .S8(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
    .I10(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
    .S16(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
    .E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
    .E16(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
    .E3(SB_T0_WEST_SB_OUT_B17_enable_value_O),
    .S18(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
    .S19(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
    .S2(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
    .S4(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
    .E9(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
    .I16(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
    .I12(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
    .S11(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
    .I17(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
    .I19(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
    .I18(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
    .S7(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
    .E4(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
    .E17(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
    .S5(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
    .I1(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
    .I5(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
    .E6(SB_T1_EAST_SB_OUT_B17_enable_value_O),
    .I4(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
    .I8(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
    .O(CB_MEM_output_width_17_num_2_fan_in_O),
    .E1(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
    .I15(MUX_SB_T3_WEST_SB_OUT_B17_ready_out)
);
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(stall),
    .out(Invert1_inst0_out)
);
wire [16:0] MUX_SB_T0_EAST_SB_OUT_B17_I [5:0];
assign MUX_SB_T0_EAST_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T0_EAST_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T0_EAST_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T0_EAST_SB_OUT_B17_I[2] = WIRE_SB_T4_NORTH_SB_IN_B17_O;
assign MUX_SB_T0_EAST_SB_OUT_B17_I[1] = WIRE_SB_T3_SOUTH_SB_IN_B17_O;
assign MUX_SB_T0_EAST_SB_OUT_B17_I[0] = WIRE_SB_T0_WEST_SB_IN_B17_O;
wire [5:0] MUX_SB_T0_EAST_SB_OUT_B17_valid_in;
assign MUX_SB_T0_EAST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T4_NORTH_SB_IN_B17_valid_out,WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T0_WEST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T0_EAST_SB_OUT_B17 (
    .I(MUX_SB_T0_EAST_SB_OUT_B17_I),
    .O(MUX_SB_T0_EAST_SB_OUT_B17_O),
    .ready_in(SB_T0_EAST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T0_EAST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T0_EAST_SB_OUT_B17_valid_out),
    .S(SB_T0_EAST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T0_EAST_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T0_NORTH_SB_OUT_B17_I [5:0];
assign MUX_SB_T0_NORTH_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T0_NORTH_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T0_NORTH_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T0_NORTH_SB_OUT_B17_I[2] = WIRE_SB_T0_SOUTH_SB_IN_B17_O;
assign MUX_SB_T0_NORTH_SB_OUT_B17_I[1] = WIRE_SB_T1_EAST_SB_IN_B17_O;
assign MUX_SB_T0_NORTH_SB_OUT_B17_I[0] = WIRE_SB_T0_WEST_SB_IN_B17_O;
wire [5:0] MUX_SB_T0_NORTH_SB_OUT_B17_valid_in;
assign MUX_SB_T0_NORTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T1_EAST_SB_IN_B17_valid_out,WIRE_SB_T0_WEST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T0_NORTH_SB_OUT_B17 (
    .I(MUX_SB_T0_NORTH_SB_OUT_B17_I),
    .O(MUX_SB_T0_NORTH_SB_OUT_B17_O),
    .ready_in(SB_T0_NORTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T0_NORTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T0_NORTH_SB_OUT_B17_valid_out),
    .S(SB_T0_NORTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T0_SOUTH_SB_OUT_B17_I [5:0];
assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[2] = WIRE_SB_T1_WEST_SB_IN_B17_O;
assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[1] = WIRE_SB_T0_NORTH_SB_IN_B17_O;
assign MUX_SB_T0_SOUTH_SB_OUT_B17_I[0] = WIRE_SB_T3_EAST_SB_IN_B17_O;
wire [5:0] MUX_SB_T0_SOUTH_SB_OUT_B17_valid_in;
assign MUX_SB_T0_SOUTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T1_WEST_SB_IN_B17_valid_out,WIRE_SB_T0_NORTH_SB_IN_B17_valid_out,WIRE_SB_T3_EAST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T0_SOUTH_SB_OUT_B17 (
    .I(MUX_SB_T0_SOUTH_SB_OUT_B17_I),
    .O(MUX_SB_T0_SOUTH_SB_OUT_B17_O),
    .ready_in(SB_T0_SOUTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T0_SOUTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T0_SOUTH_SB_OUT_B17_valid_out),
    .S(SB_T0_SOUTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T0_WEST_SB_OUT_B17_I [5:0];
assign MUX_SB_T0_WEST_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T0_WEST_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T0_WEST_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T0_WEST_SB_OUT_B17_I[2] = WIRE_SB_T0_EAST_SB_IN_B17_O;
assign MUX_SB_T0_WEST_SB_OUT_B17_I[1] = WIRE_SB_T4_SOUTH_SB_IN_B17_O;
assign MUX_SB_T0_WEST_SB_OUT_B17_I[0] = WIRE_SB_T0_NORTH_SB_IN_B17_O;
wire [5:0] MUX_SB_T0_WEST_SB_OUT_B17_valid_in;
assign MUX_SB_T0_WEST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T0_EAST_SB_IN_B17_valid_out,WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T0_NORTH_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T0_WEST_SB_OUT_B17 (
    .I(MUX_SB_T0_WEST_SB_OUT_B17_I),
    .O(MUX_SB_T0_WEST_SB_OUT_B17_O),
    .ready_in(SB_T0_WEST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T0_WEST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T0_WEST_SB_OUT_B17_valid_out),
    .S(SB_T0_WEST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T0_WEST_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T1_EAST_SB_OUT_B17_I [5:0];
assign MUX_SB_T1_EAST_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T1_EAST_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T1_EAST_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T1_EAST_SB_OUT_B17_I[2] = WIRE_SB_T2_SOUTH_SB_IN_B17_O;
assign MUX_SB_T1_EAST_SB_OUT_B17_I[1] = WIRE_SB_T1_WEST_SB_IN_B17_O;
assign MUX_SB_T1_EAST_SB_OUT_B17_I[0] = WIRE_SB_T0_NORTH_SB_IN_B17_O;
wire [5:0] MUX_SB_T1_EAST_SB_OUT_B17_valid_in;
assign MUX_SB_T1_EAST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T1_WEST_SB_IN_B17_valid_out,WIRE_SB_T0_NORTH_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T1_EAST_SB_OUT_B17 (
    .I(MUX_SB_T1_EAST_SB_OUT_B17_I),
    .O(MUX_SB_T1_EAST_SB_OUT_B17_O),
    .ready_in(SB_T1_EAST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T1_EAST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T1_EAST_SB_OUT_B17_valid_out),
    .S(SB_T1_EAST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T1_EAST_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T1_NORTH_SB_OUT_B17_I [5:0];
assign MUX_SB_T1_NORTH_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T1_NORTH_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T1_NORTH_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T1_NORTH_SB_OUT_B17_I[2] = WIRE_SB_T4_WEST_SB_IN_B17_O;
assign MUX_SB_T1_NORTH_SB_OUT_B17_I[1] = WIRE_SB_T1_SOUTH_SB_IN_B17_O;
assign MUX_SB_T1_NORTH_SB_OUT_B17_I[0] = WIRE_SB_T2_EAST_SB_IN_B17_O;
wire [5:0] MUX_SB_T1_NORTH_SB_OUT_B17_valid_in;
assign MUX_SB_T1_NORTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T4_WEST_SB_IN_B17_valid_out,WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T2_EAST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T1_NORTH_SB_OUT_B17 (
    .I(MUX_SB_T1_NORTH_SB_OUT_B17_I),
    .O(MUX_SB_T1_NORTH_SB_OUT_B17_O),
    .ready_in(SB_T1_NORTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T1_NORTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T1_NORTH_SB_OUT_B17_valid_out),
    .S(SB_T1_NORTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T1_SOUTH_SB_OUT_B17_I [5:0];
assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[2] = WIRE_SB_T2_WEST_SB_IN_B17_O;
assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[1] = WIRE_SB_T1_NORTH_SB_IN_B17_O;
assign MUX_SB_T1_SOUTH_SB_OUT_B17_I[0] = WIRE_SB_T2_EAST_SB_IN_B17_O;
wire [5:0] MUX_SB_T1_SOUTH_SB_OUT_B17_valid_in;
assign MUX_SB_T1_SOUTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T2_WEST_SB_IN_B17_valid_out,WIRE_SB_T1_NORTH_SB_IN_B17_valid_out,WIRE_SB_T2_EAST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T1_SOUTH_SB_OUT_B17 (
    .I(MUX_SB_T1_SOUTH_SB_OUT_B17_I),
    .O(MUX_SB_T1_SOUTH_SB_OUT_B17_O),
    .ready_in(SB_T1_SOUTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T1_SOUTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T1_SOUTH_SB_OUT_B17_valid_out),
    .S(SB_T1_SOUTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T1_WEST_SB_OUT_B17_I [5:0];
assign MUX_SB_T1_WEST_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T1_WEST_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T1_WEST_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T1_WEST_SB_OUT_B17_I[2] = WIRE_SB_T1_EAST_SB_IN_B17_O;
assign MUX_SB_T1_WEST_SB_OUT_B17_I[1] = WIRE_SB_T0_SOUTH_SB_IN_B17_O;
assign MUX_SB_T1_WEST_SB_OUT_B17_I[0] = WIRE_SB_T4_NORTH_SB_IN_B17_O;
wire [5:0] MUX_SB_T1_WEST_SB_OUT_B17_valid_in;
assign MUX_SB_T1_WEST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T1_EAST_SB_IN_B17_valid_out,WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T4_NORTH_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T1_WEST_SB_OUT_B17 (
    .I(MUX_SB_T1_WEST_SB_OUT_B17_I),
    .O(MUX_SB_T1_WEST_SB_OUT_B17_O),
    .ready_in(SB_T1_WEST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T1_WEST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T1_WEST_SB_OUT_B17_valid_out),
    .S(SB_T1_WEST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T1_WEST_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T2_EAST_SB_OUT_B17_I [5:0];
assign MUX_SB_T2_EAST_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T2_EAST_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T2_EAST_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T2_EAST_SB_OUT_B17_I[2] = WIRE_SB_T2_WEST_SB_IN_B17_O;
assign MUX_SB_T2_EAST_SB_OUT_B17_I[1] = WIRE_SB_T1_SOUTH_SB_IN_B17_O;
assign MUX_SB_T2_EAST_SB_OUT_B17_I[0] = WIRE_SB_T1_NORTH_SB_IN_B17_O;
wire [5:0] MUX_SB_T2_EAST_SB_OUT_B17_valid_in;
assign MUX_SB_T2_EAST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T2_WEST_SB_IN_B17_valid_out,WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T1_NORTH_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T2_EAST_SB_OUT_B17 (
    .I(MUX_SB_T2_EAST_SB_OUT_B17_I),
    .O(MUX_SB_T2_EAST_SB_OUT_B17_O),
    .ready_in(SB_T2_EAST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T2_EAST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T2_EAST_SB_OUT_B17_valid_out),
    .S(SB_T2_EAST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T2_EAST_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T2_NORTH_SB_OUT_B17_I [5:0];
assign MUX_SB_T2_NORTH_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T2_NORTH_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T2_NORTH_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T2_NORTH_SB_OUT_B17_I[2] = WIRE_SB_T3_WEST_SB_IN_B17_O;
assign MUX_SB_T2_NORTH_SB_OUT_B17_I[1] = WIRE_SB_T2_SOUTH_SB_IN_B17_O;
assign MUX_SB_T2_NORTH_SB_OUT_B17_I[0] = WIRE_SB_T3_EAST_SB_IN_B17_O;
wire [5:0] MUX_SB_T2_NORTH_SB_OUT_B17_valid_in;
assign MUX_SB_T2_NORTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T3_WEST_SB_IN_B17_valid_out,WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T3_EAST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T2_NORTH_SB_OUT_B17 (
    .I(MUX_SB_T2_NORTH_SB_OUT_B17_I),
    .O(MUX_SB_T2_NORTH_SB_OUT_B17_O),
    .ready_in(SB_T2_NORTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T2_NORTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T2_NORTH_SB_OUT_B17_valid_out),
    .S(SB_T2_NORTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T2_SOUTH_SB_OUT_B17_I [5:0];
assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[2] = WIRE_SB_T3_WEST_SB_IN_B17_O;
assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[1] = WIRE_SB_T2_NORTH_SB_IN_B17_O;
assign MUX_SB_T2_SOUTH_SB_OUT_B17_I[0] = WIRE_SB_T1_EAST_SB_IN_B17_O;
wire [5:0] MUX_SB_T2_SOUTH_SB_OUT_B17_valid_in;
assign MUX_SB_T2_SOUTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T3_WEST_SB_IN_B17_valid_out,WIRE_SB_T2_NORTH_SB_IN_B17_valid_out,WIRE_SB_T1_EAST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T2_SOUTH_SB_OUT_B17 (
    .I(MUX_SB_T2_SOUTH_SB_OUT_B17_I),
    .O(MUX_SB_T2_SOUTH_SB_OUT_B17_O),
    .ready_in(SB_T2_SOUTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T2_SOUTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T2_SOUTH_SB_OUT_B17_valid_out),
    .S(SB_T2_SOUTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T2_WEST_SB_OUT_B17_I [5:0];
assign MUX_SB_T2_WEST_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T2_WEST_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T2_WEST_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T2_WEST_SB_OUT_B17_I[2] = WIRE_SB_T2_EAST_SB_IN_B17_O;
assign MUX_SB_T2_WEST_SB_OUT_B17_I[1] = WIRE_SB_T1_SOUTH_SB_IN_B17_O;
assign MUX_SB_T2_WEST_SB_OUT_B17_I[0] = WIRE_SB_T3_NORTH_SB_IN_B17_O;
wire [5:0] MUX_SB_T2_WEST_SB_OUT_B17_valid_in;
assign MUX_SB_T2_WEST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T2_EAST_SB_IN_B17_valid_out,WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T3_NORTH_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T2_WEST_SB_OUT_B17 (
    .I(MUX_SB_T2_WEST_SB_OUT_B17_I),
    .O(MUX_SB_T2_WEST_SB_OUT_B17_O),
    .ready_in(SB_T2_WEST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T2_WEST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T2_WEST_SB_OUT_B17_valid_out),
    .S(SB_T2_WEST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T2_WEST_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T3_EAST_SB_OUT_B17_I [5:0];
assign MUX_SB_T3_EAST_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T3_EAST_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T3_EAST_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T3_EAST_SB_OUT_B17_I[2] = WIRE_SB_T3_WEST_SB_IN_B17_O;
assign MUX_SB_T3_EAST_SB_OUT_B17_I[1] = WIRE_SB_T2_NORTH_SB_IN_B17_O;
assign MUX_SB_T3_EAST_SB_OUT_B17_I[0] = WIRE_SB_T0_SOUTH_SB_IN_B17_O;
wire [5:0] MUX_SB_T3_EAST_SB_OUT_B17_valid_in;
assign MUX_SB_T3_EAST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T3_WEST_SB_IN_B17_valid_out,WIRE_SB_T2_NORTH_SB_IN_B17_valid_out,WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T3_EAST_SB_OUT_B17 (
    .I(MUX_SB_T3_EAST_SB_OUT_B17_I),
    .O(MUX_SB_T3_EAST_SB_OUT_B17_O),
    .ready_in(SB_T3_EAST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T3_EAST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T3_EAST_SB_OUT_B17_valid_out),
    .S(SB_T3_EAST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T3_EAST_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T3_NORTH_SB_OUT_B17_I [5:0];
assign MUX_SB_T3_NORTH_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T3_NORTH_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T3_NORTH_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T3_NORTH_SB_OUT_B17_I[2] = WIRE_SB_T3_SOUTH_SB_IN_B17_O;
assign MUX_SB_T3_NORTH_SB_OUT_B17_I[1] = WIRE_SB_T4_EAST_SB_IN_B17_O;
assign MUX_SB_T3_NORTH_SB_OUT_B17_I[0] = WIRE_SB_T2_WEST_SB_IN_B17_O;
wire [5:0] MUX_SB_T3_NORTH_SB_OUT_B17_valid_in;
assign MUX_SB_T3_NORTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T4_EAST_SB_IN_B17_valid_out,WIRE_SB_T2_WEST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T3_NORTH_SB_OUT_B17 (
    .I(MUX_SB_T3_NORTH_SB_OUT_B17_I),
    .O(MUX_SB_T3_NORTH_SB_OUT_B17_O),
    .ready_in(SB_T3_NORTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T3_NORTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T3_NORTH_SB_OUT_B17_valid_out),
    .S(SB_T3_NORTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T3_SOUTH_SB_OUT_B17_I [5:0];
assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[2] = WIRE_SB_T4_WEST_SB_IN_B17_O;
assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[1] = WIRE_SB_T3_NORTH_SB_IN_B17_O;
assign MUX_SB_T3_SOUTH_SB_OUT_B17_I[0] = WIRE_SB_T0_EAST_SB_IN_B17_O;
wire [5:0] MUX_SB_T3_SOUTH_SB_OUT_B17_valid_in;
assign MUX_SB_T3_SOUTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T4_WEST_SB_IN_B17_valid_out,WIRE_SB_T3_NORTH_SB_IN_B17_valid_out,WIRE_SB_T0_EAST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T3_SOUTH_SB_OUT_B17 (
    .I(MUX_SB_T3_SOUTH_SB_OUT_B17_I),
    .O(MUX_SB_T3_SOUTH_SB_OUT_B17_O),
    .ready_in(SB_T3_SOUTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T3_SOUTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T3_SOUTH_SB_OUT_B17_valid_out),
    .S(SB_T3_SOUTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T3_WEST_SB_OUT_B17_I [5:0];
assign MUX_SB_T3_WEST_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T3_WEST_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T3_WEST_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T3_WEST_SB_OUT_B17_I[2] = WIRE_SB_T3_EAST_SB_IN_B17_O;
assign MUX_SB_T3_WEST_SB_OUT_B17_I[1] = WIRE_SB_T2_SOUTH_SB_IN_B17_O;
assign MUX_SB_T3_WEST_SB_OUT_B17_I[0] = WIRE_SB_T2_NORTH_SB_IN_B17_O;
wire [5:0] MUX_SB_T3_WEST_SB_OUT_B17_valid_in;
assign MUX_SB_T3_WEST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T3_EAST_SB_IN_B17_valid_out,WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T2_NORTH_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T3_WEST_SB_OUT_B17 (
    .I(MUX_SB_T3_WEST_SB_OUT_B17_I),
    .O(MUX_SB_T3_WEST_SB_OUT_B17_O),
    .ready_in(SB_T3_WEST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T3_WEST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T3_WEST_SB_OUT_B17_valid_out),
    .S(SB_T3_WEST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T3_WEST_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T4_EAST_SB_OUT_B17_I [5:0];
assign MUX_SB_T4_EAST_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T4_EAST_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T4_EAST_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T4_EAST_SB_OUT_B17_I[2] = WIRE_SB_T4_WEST_SB_IN_B17_O;
assign MUX_SB_T4_EAST_SB_OUT_B17_I[1] = WIRE_SB_T4_SOUTH_SB_IN_B17_O;
assign MUX_SB_T4_EAST_SB_OUT_B17_I[0] = WIRE_SB_T3_NORTH_SB_IN_B17_O;
wire [5:0] MUX_SB_T4_EAST_SB_OUT_B17_valid_in;
assign MUX_SB_T4_EAST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T4_WEST_SB_IN_B17_valid_out,WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T3_NORTH_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T4_EAST_SB_OUT_B17 (
    .I(MUX_SB_T4_EAST_SB_OUT_B17_I),
    .O(MUX_SB_T4_EAST_SB_OUT_B17_O),
    .ready_in(SB_T4_EAST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T4_EAST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T4_EAST_SB_OUT_B17_valid_out),
    .S(SB_T4_EAST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T4_EAST_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T4_NORTH_SB_OUT_B17_I [5:0];
assign MUX_SB_T4_NORTH_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T4_NORTH_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T4_NORTH_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T4_NORTH_SB_OUT_B17_I[2] = WIRE_SB_T4_SOUTH_SB_IN_B17_O;
assign MUX_SB_T4_NORTH_SB_OUT_B17_I[1] = WIRE_SB_T0_EAST_SB_IN_B17_O;
assign MUX_SB_T4_NORTH_SB_OUT_B17_I[0] = WIRE_SB_T1_WEST_SB_IN_B17_O;
wire [5:0] MUX_SB_T4_NORTH_SB_OUT_B17_valid_in;
assign MUX_SB_T4_NORTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T0_EAST_SB_IN_B17_valid_out,WIRE_SB_T1_WEST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T4_NORTH_SB_OUT_B17 (
    .I(MUX_SB_T4_NORTH_SB_OUT_B17_I),
    .O(MUX_SB_T4_NORTH_SB_OUT_B17_O),
    .ready_in(SB_T4_NORTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T4_NORTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T4_NORTH_SB_OUT_B17_valid_out),
    .S(SB_T4_NORTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T4_SOUTH_SB_OUT_B17_I [5:0];
assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[2] = WIRE_SB_T4_NORTH_SB_IN_B17_O;
assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[1] = WIRE_SB_T4_EAST_SB_IN_B17_O;
assign MUX_SB_T4_SOUTH_SB_OUT_B17_I[0] = WIRE_SB_T0_WEST_SB_IN_B17_O;
wire [5:0] MUX_SB_T4_SOUTH_SB_OUT_B17_valid_in;
assign MUX_SB_T4_SOUTH_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T4_NORTH_SB_IN_B17_valid_out,WIRE_SB_T4_EAST_SB_IN_B17_valid_out,WIRE_SB_T0_WEST_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T4_SOUTH_SB_OUT_B17 (
    .I(MUX_SB_T4_SOUTH_SB_OUT_B17_I),
    .O(MUX_SB_T4_SOUTH_SB_OUT_B17_O),
    .ready_in(SB_T4_SOUTH_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T4_SOUTH_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T4_SOUTH_SB_OUT_B17_valid_out),
    .S(SB_T4_SOUTH_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel)
);
wire [16:0] MUX_SB_T4_WEST_SB_OUT_B17_I [5:0];
assign MUX_SB_T4_WEST_SB_OUT_B17_I[5] = MEM_output_width_17_num_2;
assign MUX_SB_T4_WEST_SB_OUT_B17_I[4] = MEM_output_width_17_num_1;
assign MUX_SB_T4_WEST_SB_OUT_B17_I[3] = MEM_output_width_17_num_0;
assign MUX_SB_T4_WEST_SB_OUT_B17_I[2] = WIRE_SB_T4_EAST_SB_IN_B17_O;
assign MUX_SB_T4_WEST_SB_OUT_B17_I[1] = WIRE_SB_T3_SOUTH_SB_IN_B17_O;
assign MUX_SB_T4_WEST_SB_OUT_B17_I[0] = WIRE_SB_T1_NORTH_SB_IN_B17_O;
wire [5:0] MUX_SB_T4_WEST_SB_OUT_B17_valid_in;
assign MUX_SB_T4_WEST_SB_OUT_B17_valid_in = {MEM_output_width_17_num_2_valid,MEM_output_width_17_num_1_valid,MEM_output_width_17_num_0_valid,WIRE_SB_T4_EAST_SB_IN_B17_valid_out,WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out,WIRE_SB_T1_NORTH_SB_IN_B17_valid_out};
mux_aoi_ready_valid_6_17 MUX_SB_T4_WEST_SB_OUT_B17 (
    .I(MUX_SB_T4_WEST_SB_OUT_B17_I),
    .O(MUX_SB_T4_WEST_SB_OUT_B17_O),
    .ready_in(SB_T4_WEST_SB_OUT_B17_FANOUT_O[0]),
    .ready_out(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
    .valid_in(MUX_SB_T4_WEST_SB_OUT_B17_valid_in),
    .valid_out(MUX_SB_T4_WEST_SB_OUT_B17_valid_out),
    .S(SB_T4_WEST_SB_OUT_B17_sel_value_O),
    .out_sel(MUX_SB_T4_WEST_SB_OUT_B17_out_sel)
);
SplitFifo_17 REG_T0_EAST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T0_EAST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T0_EAST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T0_EAST_B17_fifo_value_O[0]),
    .end_fifo(REG_T0_EAST_B17_end_value_O[0]),
    .data_in(MUX_SB_T0_EAST_SB_OUT_B17_O),
    .ready1(RMUX_T0_EAST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T0_EAST_SB_OUT_B17_valid_out),
    .data_out(REG_T0_EAST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T0_EAST_B17_start_value_O[0]),
    .clk_en(and1_inst2_out[0])
);
SliceWrapper_32_0_1 REG_T0_EAST_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T0_EAST_B17_end_value_O)
);
SliceWrapper_32_1_2 REG_T0_EAST_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T0_EAST_B17_fifo_value_O)
);
SliceWrapper_32_2_3 REG_T0_EAST_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T0_EAST_B17_start_value_O)
);
SplitFifo_17 REG_T0_NORTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T0_NORTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T0_NORTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T0_NORTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T0_NORTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T0_NORTH_SB_OUT_B17_O),
    .ready1(RMUX_T0_NORTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T0_NORTH_SB_OUT_B17_valid_out),
    .data_out(REG_T0_NORTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T0_NORTH_B17_start_value_O[0]),
    .clk_en(and1_inst0_out[0])
);
SliceWrapper_32_3_4 REG_T0_NORTH_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T0_NORTH_B17_end_value_O)
);
SliceWrapper_32_4_5 REG_T0_NORTH_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T0_NORTH_B17_fifo_value_O)
);
SliceWrapper_32_5_6 REG_T0_NORTH_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T0_NORTH_B17_start_value_O)
);
SplitFifo_17 REG_T0_SOUTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T0_SOUTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T0_SOUTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T0_SOUTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T0_SOUTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T0_SOUTH_SB_OUT_B17_O),
    .ready1(RMUX_T0_SOUTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T0_SOUTH_SB_OUT_B17_valid_out),
    .data_out(REG_T0_SOUTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T0_SOUTH_B17_start_value_O[0]),
    .clk_en(and1_inst1_out[0])
);
SliceWrapper_32_6_7 REG_T0_SOUTH_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T0_SOUTH_B17_end_value_O)
);
SliceWrapper_32_7_8 REG_T0_SOUTH_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T0_SOUTH_B17_fifo_value_O)
);
SliceWrapper_32_8_9 REG_T0_SOUTH_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T0_SOUTH_B17_start_value_O)
);
SplitFifo_17 REG_T0_WEST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T0_WEST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T0_WEST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T0_WEST_B17_fifo_value_O[0]),
    .end_fifo(REG_T0_WEST_B17_end_value_O[0]),
    .data_in(MUX_SB_T0_WEST_SB_OUT_B17_O),
    .ready1(RMUX_T0_WEST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T0_WEST_SB_OUT_B17_valid_out),
    .data_out(REG_T0_WEST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T0_WEST_B17_start_value_O[0]),
    .clk_en(and1_inst3_out[0])
);
SliceWrapper_32_9_10 REG_T0_WEST_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T0_WEST_B17_end_value_O)
);
SliceWrapper_32_10_11 REG_T0_WEST_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T0_WEST_B17_fifo_value_O)
);
SliceWrapper_32_11_12 REG_T0_WEST_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T0_WEST_B17_start_value_O)
);
SplitFifo_17 REG_T1_EAST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T1_EAST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T1_EAST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T1_EAST_B17_fifo_value_O[0]),
    .end_fifo(REG_T1_EAST_B17_end_value_O[0]),
    .data_in(MUX_SB_T1_EAST_SB_OUT_B17_O),
    .ready1(RMUX_T1_EAST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T1_EAST_SB_OUT_B17_valid_out),
    .data_out(REG_T1_EAST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T1_EAST_B17_start_value_O[0]),
    .clk_en(and1_inst6_out[0])
);
SliceWrapper_32_12_13 REG_T1_EAST_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T1_EAST_B17_end_value_O)
);
SliceWrapper_32_13_14 REG_T1_EAST_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T1_EAST_B17_fifo_value_O)
);
SliceWrapper_32_14_15 REG_T1_EAST_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T1_EAST_B17_start_value_O)
);
SplitFifo_17 REG_T1_NORTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T1_NORTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T1_NORTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T1_NORTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T1_NORTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T1_NORTH_SB_OUT_B17_O),
    .ready1(RMUX_T1_NORTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T1_NORTH_SB_OUT_B17_valid_out),
    .data_out(REG_T1_NORTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T1_NORTH_B17_start_value_O[0]),
    .clk_en(and1_inst4_out[0])
);
SliceWrapper_32_15_16 REG_T1_NORTH_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T1_NORTH_B17_end_value_O)
);
SliceWrapper_32_16_17 REG_T1_NORTH_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T1_NORTH_B17_fifo_value_O)
);
SliceWrapper_32_17_18 REG_T1_NORTH_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T1_NORTH_B17_start_value_O)
);
SplitFifo_17 REG_T1_SOUTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T1_SOUTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T1_SOUTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T1_SOUTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T1_SOUTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T1_SOUTH_SB_OUT_B17_O),
    .ready1(RMUX_T1_SOUTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T1_SOUTH_SB_OUT_B17_valid_out),
    .data_out(REG_T1_SOUTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T1_SOUTH_B17_start_value_O[0]),
    .clk_en(and1_inst5_out[0])
);
SliceWrapper_32_18_19 REG_T1_SOUTH_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T1_SOUTH_B17_end_value_O)
);
SliceWrapper_32_19_20 REG_T1_SOUTH_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T1_SOUTH_B17_fifo_value_O)
);
SliceWrapper_32_20_21 REG_T1_SOUTH_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T1_SOUTH_B17_start_value_O)
);
SplitFifo_17 REG_T1_WEST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T1_WEST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T1_WEST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T1_WEST_B17_fifo_value_O[0]),
    .end_fifo(REG_T1_WEST_B17_end_value_O[0]),
    .data_in(MUX_SB_T1_WEST_SB_OUT_B17_O),
    .ready1(RMUX_T1_WEST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T1_WEST_SB_OUT_B17_valid_out),
    .data_out(REG_T1_WEST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T1_WEST_B17_start_value_O[0]),
    .clk_en(and1_inst7_out[0])
);
SliceWrapper_32_21_22 REG_T1_WEST_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T1_WEST_B17_end_value_O)
);
SliceWrapper_32_22_23 REG_T1_WEST_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T1_WEST_B17_fifo_value_O)
);
SliceWrapper_32_23_24 REG_T1_WEST_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T1_WEST_B17_start_value_O)
);
SplitFifo_17 REG_T2_EAST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T2_EAST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T2_EAST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T2_EAST_B17_fifo_value_O[0]),
    .end_fifo(REG_T2_EAST_B17_end_value_O[0]),
    .data_in(MUX_SB_T2_EAST_SB_OUT_B17_O),
    .ready1(RMUX_T2_EAST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T2_EAST_SB_OUT_B17_valid_out),
    .data_out(REG_T2_EAST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T2_EAST_B17_start_value_O[0]),
    .clk_en(and1_inst10_out[0])
);
SliceWrapper_32_24_25 REG_T2_EAST_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T2_EAST_B17_end_value_O)
);
SliceWrapper_32_25_26 REG_T2_EAST_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T2_EAST_B17_fifo_value_O)
);
SliceWrapper_32_26_27 REG_T2_EAST_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T2_EAST_B17_start_value_O)
);
SplitFifo_17 REG_T2_NORTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T2_NORTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T2_NORTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T2_NORTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T2_NORTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T2_NORTH_SB_OUT_B17_O),
    .ready1(RMUX_T2_NORTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T2_NORTH_SB_OUT_B17_valid_out),
    .data_out(REG_T2_NORTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T2_NORTH_B17_start_value_O[0]),
    .clk_en(and1_inst8_out[0])
);
SliceWrapper_32_27_28 REG_T2_NORTH_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T2_NORTH_B17_end_value_O)
);
SliceWrapper_32_28_29 REG_T2_NORTH_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T2_NORTH_B17_fifo_value_O)
);
SliceWrapper_32_29_30 REG_T2_NORTH_B17_start_value (
    .I(config_reg_0_O),
    .O(REG_T2_NORTH_B17_start_value_O)
);
SplitFifo_17 REG_T2_SOUTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T2_SOUTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T2_SOUTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T2_SOUTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T2_SOUTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T2_SOUTH_SB_OUT_B17_O),
    .ready1(RMUX_T2_SOUTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T2_SOUTH_SB_OUT_B17_valid_out),
    .data_out(REG_T2_SOUTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T2_SOUTH_B17_start_value_O[0]),
    .clk_en(and1_inst9_out[0])
);
SliceWrapper_32_30_31 REG_T2_SOUTH_B17_end_value (
    .I(config_reg_0_O),
    .O(REG_T2_SOUTH_B17_end_value_O)
);
SliceWrapper_32_31_32 REG_T2_SOUTH_B17_fifo_value (
    .I(config_reg_0_O),
    .O(REG_T2_SOUTH_B17_fifo_value_O)
);
SliceWrapper_32_0_1 REG_T2_SOUTH_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T2_SOUTH_B17_start_value_O)
);
SplitFifo_17 REG_T2_WEST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T2_WEST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T2_WEST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T2_WEST_B17_fifo_value_O[0]),
    .end_fifo(REG_T2_WEST_B17_end_value_O[0]),
    .data_in(MUX_SB_T2_WEST_SB_OUT_B17_O),
    .ready1(RMUX_T2_WEST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T2_WEST_SB_OUT_B17_valid_out),
    .data_out(REG_T2_WEST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T2_WEST_B17_start_value_O[0]),
    .clk_en(and1_inst11_out[0])
);
SliceWrapper_32_1_2 REG_T2_WEST_B17_end_value (
    .I(config_reg_1_O),
    .O(REG_T2_WEST_B17_end_value_O)
);
SliceWrapper_32_2_3 REG_T2_WEST_B17_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T2_WEST_B17_fifo_value_O)
);
SliceWrapper_32_3_4 REG_T2_WEST_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T2_WEST_B17_start_value_O)
);
SplitFifo_17 REG_T3_EAST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T3_EAST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T3_EAST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T3_EAST_B17_fifo_value_O[0]),
    .end_fifo(REG_T3_EAST_B17_end_value_O[0]),
    .data_in(MUX_SB_T3_EAST_SB_OUT_B17_O),
    .ready1(RMUX_T3_EAST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T3_EAST_SB_OUT_B17_valid_out),
    .data_out(REG_T3_EAST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T3_EAST_B17_start_value_O[0]),
    .clk_en(and1_inst14_out[0])
);
SliceWrapper_32_4_5 REG_T3_EAST_B17_end_value (
    .I(config_reg_1_O),
    .O(REG_T3_EAST_B17_end_value_O)
);
SliceWrapper_32_5_6 REG_T3_EAST_B17_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T3_EAST_B17_fifo_value_O)
);
SliceWrapper_32_6_7 REG_T3_EAST_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T3_EAST_B17_start_value_O)
);
SplitFifo_17 REG_T3_NORTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T3_NORTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T3_NORTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T3_NORTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T3_NORTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T3_NORTH_SB_OUT_B17_O),
    .ready1(RMUX_T3_NORTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T3_NORTH_SB_OUT_B17_valid_out),
    .data_out(REG_T3_NORTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T3_NORTH_B17_start_value_O[0]),
    .clk_en(and1_inst12_out[0])
);
SliceWrapper_32_7_8 REG_T3_NORTH_B17_end_value (
    .I(config_reg_1_O),
    .O(REG_T3_NORTH_B17_end_value_O)
);
SliceWrapper_32_8_9 REG_T3_NORTH_B17_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T3_NORTH_B17_fifo_value_O)
);
SliceWrapper_32_9_10 REG_T3_NORTH_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T3_NORTH_B17_start_value_O)
);
SplitFifo_17 REG_T3_SOUTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T3_SOUTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T3_SOUTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T3_SOUTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T3_SOUTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T3_SOUTH_SB_OUT_B17_O),
    .ready1(RMUX_T3_SOUTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T3_SOUTH_SB_OUT_B17_valid_out),
    .data_out(REG_T3_SOUTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T3_SOUTH_B17_start_value_O[0]),
    .clk_en(and1_inst13_out[0])
);
SliceWrapper_32_10_11 REG_T3_SOUTH_B17_end_value (
    .I(config_reg_1_O),
    .O(REG_T3_SOUTH_B17_end_value_O)
);
SliceWrapper_32_11_12 REG_T3_SOUTH_B17_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T3_SOUTH_B17_fifo_value_O)
);
SliceWrapper_32_12_13 REG_T3_SOUTH_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T3_SOUTH_B17_start_value_O)
);
SplitFifo_17 REG_T3_WEST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T3_WEST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T3_WEST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T3_WEST_B17_fifo_value_O[0]),
    .end_fifo(REG_T3_WEST_B17_end_value_O[0]),
    .data_in(MUX_SB_T3_WEST_SB_OUT_B17_O),
    .ready1(RMUX_T3_WEST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T3_WEST_SB_OUT_B17_valid_out),
    .data_out(REG_T3_WEST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T3_WEST_B17_start_value_O[0]),
    .clk_en(and1_inst15_out[0])
);
SliceWrapper_32_13_14 REG_T3_WEST_B17_end_value (
    .I(config_reg_1_O),
    .O(REG_T3_WEST_B17_end_value_O)
);
SliceWrapper_32_14_15 REG_T3_WEST_B17_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T3_WEST_B17_fifo_value_O)
);
SliceWrapper_32_15_16 REG_T3_WEST_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T3_WEST_B17_start_value_O)
);
SplitFifo_17 REG_T4_EAST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T4_EAST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T4_EAST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T4_EAST_B17_fifo_value_O[0]),
    .end_fifo(REG_T4_EAST_B17_end_value_O[0]),
    .data_in(MUX_SB_T4_EAST_SB_OUT_B17_O),
    .ready1(RMUX_T4_EAST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T4_EAST_SB_OUT_B17_valid_out),
    .data_out(REG_T4_EAST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T4_EAST_B17_start_value_O[0]),
    .clk_en(and1_inst18_out[0])
);
SliceWrapper_32_16_17 REG_T4_EAST_B17_end_value (
    .I(config_reg_1_O),
    .O(REG_T4_EAST_B17_end_value_O)
);
SliceWrapper_32_17_18 REG_T4_EAST_B17_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T4_EAST_B17_fifo_value_O)
);
SliceWrapper_32_18_19 REG_T4_EAST_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T4_EAST_B17_start_value_O)
);
SplitFifo_17 REG_T4_NORTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T4_NORTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T4_NORTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T4_NORTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T4_NORTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T4_NORTH_SB_OUT_B17_O),
    .ready1(RMUX_T4_NORTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T4_NORTH_SB_OUT_B17_valid_out),
    .data_out(REG_T4_NORTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T4_NORTH_B17_start_value_O[0]),
    .clk_en(and1_inst16_out[0])
);
SliceWrapper_32_19_20 REG_T4_NORTH_B17_end_value (
    .I(config_reg_1_O),
    .O(REG_T4_NORTH_B17_end_value_O)
);
SliceWrapper_32_20_21 REG_T4_NORTH_B17_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T4_NORTH_B17_fifo_value_O)
);
SliceWrapper_32_21_22 REG_T4_NORTH_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T4_NORTH_B17_start_value_O)
);
SplitFifo_17 REG_T4_SOUTH_B17$SplitFifo_17_inst0 (
    .ready0(REG_T4_SOUTH_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T4_SOUTH_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T4_SOUTH_B17_fifo_value_O[0]),
    .end_fifo(REG_T4_SOUTH_B17_end_value_O[0]),
    .data_in(MUX_SB_T4_SOUTH_SB_OUT_B17_O),
    .ready1(RMUX_T4_SOUTH_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T4_SOUTH_SB_OUT_B17_valid_out),
    .data_out(REG_T4_SOUTH_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T4_SOUTH_B17_start_value_O[0]),
    .clk_en(and1_inst17_out[0])
);
SliceWrapper_32_22_23 REG_T4_SOUTH_B17_end_value (
    .I(config_reg_1_O),
    .O(REG_T4_SOUTH_B17_end_value_O)
);
SliceWrapper_32_23_24 REG_T4_SOUTH_B17_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T4_SOUTH_B17_fifo_value_O)
);
SliceWrapper_32_24_25 REG_T4_SOUTH_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T4_SOUTH_B17_start_value_O)
);
SplitFifo_17 REG_T4_WEST_B17$SplitFifo_17_inst0 (
    .ready0(REG_T4_WEST_B17$SplitFifo_17_inst0_ready0),
    .rst(reset),
    .valid1(REG_T4_WEST_B17$SplitFifo_17_inst0_valid1),
    .fifo_en(REG_T4_WEST_B17_fifo_value_O[0]),
    .end_fifo(REG_T4_WEST_B17_end_value_O[0]),
    .data_in(MUX_SB_T4_WEST_SB_OUT_B17_O),
    .ready1(RMUX_T4_WEST_B17_ready_out),
    .clk(clk),
    .valid0(MUX_SB_T4_WEST_SB_OUT_B17_valid_out),
    .data_out(REG_T4_WEST_B17$SplitFifo_17_inst0_data_out),
    .start_fifo(REG_T4_WEST_B17_start_value_O[0]),
    .clk_en(and1_inst19_out[0])
);
SliceWrapper_32_25_26 REG_T4_WEST_B17_end_value (
    .I(config_reg_1_O),
    .O(REG_T4_WEST_B17_end_value_O)
);
SliceWrapper_32_26_27 REG_T4_WEST_B17_fifo_value (
    .I(config_reg_1_O),
    .O(REG_T4_WEST_B17_fifo_value_O)
);
SliceWrapper_32_27_28 REG_T4_WEST_B17_start_value (
    .I(config_reg_1_O),
    .O(REG_T4_WEST_B17_start_value_O)
);
wire [16:0] RMUX_T0_EAST_B17_I [1:0];
assign RMUX_T0_EAST_B17_I[1] = REG_T0_EAST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T0_EAST_B17_I[0] = MUX_SB_T0_EAST_SB_OUT_B17_O;
wire [1:0] RMUX_T0_EAST_B17_valid_in;
assign RMUX_T0_EAST_B17_valid_in = {REG_T0_EAST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T0_EAST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T0_EAST_B17 (
    .I(RMUX_T0_EAST_B17_I),
    .O(RMUX_T0_EAST_B17_O),
    .ready_in(SB_T0_EAST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T0_EAST_B17_ready_out),
    .valid_in(RMUX_T0_EAST_B17_valid_in),
    .valid_out(RMUX_T0_EAST_B17_valid_out),
    .S(RMUX_T0_EAST_B17_sel_value_O),
    .out_sel(RMUX_T0_EAST_B17_out_sel)
);
SliceWrapper_32_28_29 RMUX_T0_EAST_B17_sel_value (
    .I(config_reg_1_O),
    .O(RMUX_T0_EAST_B17_sel_value_O)
);
wire [16:0] RMUX_T0_NORTH_B17_I [1:0];
assign RMUX_T0_NORTH_B17_I[1] = REG_T0_NORTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T0_NORTH_B17_I[0] = MUX_SB_T0_NORTH_SB_OUT_B17_O;
wire [1:0] RMUX_T0_NORTH_B17_valid_in;
assign RMUX_T0_NORTH_B17_valid_in = {REG_T0_NORTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T0_NORTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T0_NORTH_B17 (
    .I(RMUX_T0_NORTH_B17_I),
    .O(RMUX_T0_NORTH_B17_O),
    .ready_in(SB_T0_NORTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T0_NORTH_B17_ready_out),
    .valid_in(RMUX_T0_NORTH_B17_valid_in),
    .valid_out(RMUX_T0_NORTH_B17_valid_out),
    .S(RMUX_T0_NORTH_B17_sel_value_O),
    .out_sel(RMUX_T0_NORTH_B17_out_sel)
);
SliceWrapper_32_29_30 RMUX_T0_NORTH_B17_sel_value (
    .I(config_reg_1_O),
    .O(RMUX_T0_NORTH_B17_sel_value_O)
);
wire [16:0] RMUX_T0_SOUTH_B17_I [1:0];
assign RMUX_T0_SOUTH_B17_I[1] = REG_T0_SOUTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T0_SOUTH_B17_I[0] = MUX_SB_T0_SOUTH_SB_OUT_B17_O;
wire [1:0] RMUX_T0_SOUTH_B17_valid_in;
assign RMUX_T0_SOUTH_B17_valid_in = {REG_T0_SOUTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T0_SOUTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T0_SOUTH_B17 (
    .I(RMUX_T0_SOUTH_B17_I),
    .O(RMUX_T0_SOUTH_B17_O),
    .ready_in(SB_T0_SOUTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T0_SOUTH_B17_ready_out),
    .valid_in(RMUX_T0_SOUTH_B17_valid_in),
    .valid_out(RMUX_T0_SOUTH_B17_valid_out),
    .S(RMUX_T0_SOUTH_B17_sel_value_O),
    .out_sel(RMUX_T0_SOUTH_B17_out_sel)
);
SliceWrapper_32_30_31 RMUX_T0_SOUTH_B17_sel_value (
    .I(config_reg_1_O),
    .O(RMUX_T0_SOUTH_B17_sel_value_O)
);
wire [16:0] RMUX_T0_WEST_B17_I [1:0];
assign RMUX_T0_WEST_B17_I[1] = REG_T0_WEST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T0_WEST_B17_I[0] = MUX_SB_T0_WEST_SB_OUT_B17_O;
wire [1:0] RMUX_T0_WEST_B17_valid_in;
assign RMUX_T0_WEST_B17_valid_in = {REG_T0_WEST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T0_WEST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T0_WEST_B17 (
    .I(RMUX_T0_WEST_B17_I),
    .O(RMUX_T0_WEST_B17_O),
    .ready_in(SB_T0_WEST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T0_WEST_B17_ready_out),
    .valid_in(RMUX_T0_WEST_B17_valid_in),
    .valid_out(RMUX_T0_WEST_B17_valid_out),
    .S(RMUX_T0_WEST_B17_sel_value_O),
    .out_sel(RMUX_T0_WEST_B17_out_sel)
);
SliceWrapper_32_31_32 RMUX_T0_WEST_B17_sel_value (
    .I(config_reg_1_O),
    .O(RMUX_T0_WEST_B17_sel_value_O)
);
wire [16:0] RMUX_T1_EAST_B17_I [1:0];
assign RMUX_T1_EAST_B17_I[1] = REG_T1_EAST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T1_EAST_B17_I[0] = MUX_SB_T1_EAST_SB_OUT_B17_O;
wire [1:0] RMUX_T1_EAST_B17_valid_in;
assign RMUX_T1_EAST_B17_valid_in = {REG_T1_EAST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T1_EAST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T1_EAST_B17 (
    .I(RMUX_T1_EAST_B17_I),
    .O(RMUX_T1_EAST_B17_O),
    .ready_in(SB_T1_EAST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T1_EAST_B17_ready_out),
    .valid_in(RMUX_T1_EAST_B17_valid_in),
    .valid_out(RMUX_T1_EAST_B17_valid_out),
    .S(RMUX_T1_EAST_B17_sel_value_O),
    .out_sel(RMUX_T1_EAST_B17_out_sel)
);
SliceWrapper_32_0_1 RMUX_T1_EAST_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T1_EAST_B17_sel_value_O)
);
wire [16:0] RMUX_T1_NORTH_B17_I [1:0];
assign RMUX_T1_NORTH_B17_I[1] = REG_T1_NORTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T1_NORTH_B17_I[0] = MUX_SB_T1_NORTH_SB_OUT_B17_O;
wire [1:0] RMUX_T1_NORTH_B17_valid_in;
assign RMUX_T1_NORTH_B17_valid_in = {REG_T1_NORTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T1_NORTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T1_NORTH_B17 (
    .I(RMUX_T1_NORTH_B17_I),
    .O(RMUX_T1_NORTH_B17_O),
    .ready_in(SB_T1_NORTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T1_NORTH_B17_ready_out),
    .valid_in(RMUX_T1_NORTH_B17_valid_in),
    .valid_out(RMUX_T1_NORTH_B17_valid_out),
    .S(RMUX_T1_NORTH_B17_sel_value_O),
    .out_sel(RMUX_T1_NORTH_B17_out_sel)
);
SliceWrapper_32_1_2 RMUX_T1_NORTH_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T1_NORTH_B17_sel_value_O)
);
wire [16:0] RMUX_T1_SOUTH_B17_I [1:0];
assign RMUX_T1_SOUTH_B17_I[1] = REG_T1_SOUTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T1_SOUTH_B17_I[0] = MUX_SB_T1_SOUTH_SB_OUT_B17_O;
wire [1:0] RMUX_T1_SOUTH_B17_valid_in;
assign RMUX_T1_SOUTH_B17_valid_in = {REG_T1_SOUTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T1_SOUTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T1_SOUTH_B17 (
    .I(RMUX_T1_SOUTH_B17_I),
    .O(RMUX_T1_SOUTH_B17_O),
    .ready_in(SB_T1_SOUTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T1_SOUTH_B17_ready_out),
    .valid_in(RMUX_T1_SOUTH_B17_valid_in),
    .valid_out(RMUX_T1_SOUTH_B17_valid_out),
    .S(RMUX_T1_SOUTH_B17_sel_value_O),
    .out_sel(RMUX_T1_SOUTH_B17_out_sel)
);
SliceWrapper_32_2_3 RMUX_T1_SOUTH_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T1_SOUTH_B17_sel_value_O)
);
wire [16:0] RMUX_T1_WEST_B17_I [1:0];
assign RMUX_T1_WEST_B17_I[1] = REG_T1_WEST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T1_WEST_B17_I[0] = MUX_SB_T1_WEST_SB_OUT_B17_O;
wire [1:0] RMUX_T1_WEST_B17_valid_in;
assign RMUX_T1_WEST_B17_valid_in = {REG_T1_WEST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T1_WEST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T1_WEST_B17 (
    .I(RMUX_T1_WEST_B17_I),
    .O(RMUX_T1_WEST_B17_O),
    .ready_in(SB_T1_WEST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T1_WEST_B17_ready_out),
    .valid_in(RMUX_T1_WEST_B17_valid_in),
    .valid_out(RMUX_T1_WEST_B17_valid_out),
    .S(RMUX_T1_WEST_B17_sel_value_O),
    .out_sel(RMUX_T1_WEST_B17_out_sel)
);
SliceWrapper_32_3_4 RMUX_T1_WEST_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T1_WEST_B17_sel_value_O)
);
wire [16:0] RMUX_T2_EAST_B17_I [1:0];
assign RMUX_T2_EAST_B17_I[1] = REG_T2_EAST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T2_EAST_B17_I[0] = MUX_SB_T2_EAST_SB_OUT_B17_O;
wire [1:0] RMUX_T2_EAST_B17_valid_in;
assign RMUX_T2_EAST_B17_valid_in = {REG_T2_EAST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T2_EAST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T2_EAST_B17 (
    .I(RMUX_T2_EAST_B17_I),
    .O(RMUX_T2_EAST_B17_O),
    .ready_in(SB_T2_EAST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T2_EAST_B17_ready_out),
    .valid_in(RMUX_T2_EAST_B17_valid_in),
    .valid_out(RMUX_T2_EAST_B17_valid_out),
    .S(RMUX_T2_EAST_B17_sel_value_O),
    .out_sel(RMUX_T2_EAST_B17_out_sel)
);
SliceWrapper_32_4_5 RMUX_T2_EAST_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T2_EAST_B17_sel_value_O)
);
wire [16:0] RMUX_T2_NORTH_B17_I [1:0];
assign RMUX_T2_NORTH_B17_I[1] = REG_T2_NORTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T2_NORTH_B17_I[0] = MUX_SB_T2_NORTH_SB_OUT_B17_O;
wire [1:0] RMUX_T2_NORTH_B17_valid_in;
assign RMUX_T2_NORTH_B17_valid_in = {REG_T2_NORTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T2_NORTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T2_NORTH_B17 (
    .I(RMUX_T2_NORTH_B17_I),
    .O(RMUX_T2_NORTH_B17_O),
    .ready_in(SB_T2_NORTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T2_NORTH_B17_ready_out),
    .valid_in(RMUX_T2_NORTH_B17_valid_in),
    .valid_out(RMUX_T2_NORTH_B17_valid_out),
    .S(RMUX_T2_NORTH_B17_sel_value_O),
    .out_sel(RMUX_T2_NORTH_B17_out_sel)
);
SliceWrapper_32_5_6 RMUX_T2_NORTH_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T2_NORTH_B17_sel_value_O)
);
wire [16:0] RMUX_T2_SOUTH_B17_I [1:0];
assign RMUX_T2_SOUTH_B17_I[1] = REG_T2_SOUTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T2_SOUTH_B17_I[0] = MUX_SB_T2_SOUTH_SB_OUT_B17_O;
wire [1:0] RMUX_T2_SOUTH_B17_valid_in;
assign RMUX_T2_SOUTH_B17_valid_in = {REG_T2_SOUTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T2_SOUTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T2_SOUTH_B17 (
    .I(RMUX_T2_SOUTH_B17_I),
    .O(RMUX_T2_SOUTH_B17_O),
    .ready_in(SB_T2_SOUTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T2_SOUTH_B17_ready_out),
    .valid_in(RMUX_T2_SOUTH_B17_valid_in),
    .valid_out(RMUX_T2_SOUTH_B17_valid_out),
    .S(RMUX_T2_SOUTH_B17_sel_value_O),
    .out_sel(RMUX_T2_SOUTH_B17_out_sel)
);
SliceWrapper_32_6_7 RMUX_T2_SOUTH_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T2_SOUTH_B17_sel_value_O)
);
wire [16:0] RMUX_T2_WEST_B17_I [1:0];
assign RMUX_T2_WEST_B17_I[1] = REG_T2_WEST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T2_WEST_B17_I[0] = MUX_SB_T2_WEST_SB_OUT_B17_O;
wire [1:0] RMUX_T2_WEST_B17_valid_in;
assign RMUX_T2_WEST_B17_valid_in = {REG_T2_WEST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T2_WEST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T2_WEST_B17 (
    .I(RMUX_T2_WEST_B17_I),
    .O(RMUX_T2_WEST_B17_O),
    .ready_in(SB_T2_WEST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T2_WEST_B17_ready_out),
    .valid_in(RMUX_T2_WEST_B17_valid_in),
    .valid_out(RMUX_T2_WEST_B17_valid_out),
    .S(RMUX_T2_WEST_B17_sel_value_O),
    .out_sel(RMUX_T2_WEST_B17_out_sel)
);
SliceWrapper_32_7_8 RMUX_T2_WEST_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T2_WEST_B17_sel_value_O)
);
wire [16:0] RMUX_T3_EAST_B17_I [1:0];
assign RMUX_T3_EAST_B17_I[1] = REG_T3_EAST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T3_EAST_B17_I[0] = MUX_SB_T3_EAST_SB_OUT_B17_O;
wire [1:0] RMUX_T3_EAST_B17_valid_in;
assign RMUX_T3_EAST_B17_valid_in = {REG_T3_EAST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T3_EAST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T3_EAST_B17 (
    .I(RMUX_T3_EAST_B17_I),
    .O(RMUX_T3_EAST_B17_O),
    .ready_in(SB_T3_EAST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T3_EAST_B17_ready_out),
    .valid_in(RMUX_T3_EAST_B17_valid_in),
    .valid_out(RMUX_T3_EAST_B17_valid_out),
    .S(RMUX_T3_EAST_B17_sel_value_O),
    .out_sel(RMUX_T3_EAST_B17_out_sel)
);
SliceWrapper_32_8_9 RMUX_T3_EAST_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T3_EAST_B17_sel_value_O)
);
wire [16:0] RMUX_T3_NORTH_B17_I [1:0];
assign RMUX_T3_NORTH_B17_I[1] = REG_T3_NORTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T3_NORTH_B17_I[0] = MUX_SB_T3_NORTH_SB_OUT_B17_O;
wire [1:0] RMUX_T3_NORTH_B17_valid_in;
assign RMUX_T3_NORTH_B17_valid_in = {REG_T3_NORTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T3_NORTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T3_NORTH_B17 (
    .I(RMUX_T3_NORTH_B17_I),
    .O(RMUX_T3_NORTH_B17_O),
    .ready_in(SB_T3_NORTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T3_NORTH_B17_ready_out),
    .valid_in(RMUX_T3_NORTH_B17_valid_in),
    .valid_out(RMUX_T3_NORTH_B17_valid_out),
    .S(RMUX_T3_NORTH_B17_sel_value_O),
    .out_sel(RMUX_T3_NORTH_B17_out_sel)
);
SliceWrapper_32_9_10 RMUX_T3_NORTH_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T3_NORTH_B17_sel_value_O)
);
wire [16:0] RMUX_T3_SOUTH_B17_I [1:0];
assign RMUX_T3_SOUTH_B17_I[1] = REG_T3_SOUTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T3_SOUTH_B17_I[0] = MUX_SB_T3_SOUTH_SB_OUT_B17_O;
wire [1:0] RMUX_T3_SOUTH_B17_valid_in;
assign RMUX_T3_SOUTH_B17_valid_in = {REG_T3_SOUTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T3_SOUTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T3_SOUTH_B17 (
    .I(RMUX_T3_SOUTH_B17_I),
    .O(RMUX_T3_SOUTH_B17_O),
    .ready_in(SB_T3_SOUTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T3_SOUTH_B17_ready_out),
    .valid_in(RMUX_T3_SOUTH_B17_valid_in),
    .valid_out(RMUX_T3_SOUTH_B17_valid_out),
    .S(RMUX_T3_SOUTH_B17_sel_value_O),
    .out_sel(RMUX_T3_SOUTH_B17_out_sel)
);
SliceWrapper_32_10_11 RMUX_T3_SOUTH_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T3_SOUTH_B17_sel_value_O)
);
wire [16:0] RMUX_T3_WEST_B17_I [1:0];
assign RMUX_T3_WEST_B17_I[1] = REG_T3_WEST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T3_WEST_B17_I[0] = MUX_SB_T3_WEST_SB_OUT_B17_O;
wire [1:0] RMUX_T3_WEST_B17_valid_in;
assign RMUX_T3_WEST_B17_valid_in = {REG_T3_WEST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T3_WEST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T3_WEST_B17 (
    .I(RMUX_T3_WEST_B17_I),
    .O(RMUX_T3_WEST_B17_O),
    .ready_in(SB_T3_WEST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T3_WEST_B17_ready_out),
    .valid_in(RMUX_T3_WEST_B17_valid_in),
    .valid_out(RMUX_T3_WEST_B17_valid_out),
    .S(RMUX_T3_WEST_B17_sel_value_O),
    .out_sel(RMUX_T3_WEST_B17_out_sel)
);
SliceWrapper_32_11_12 RMUX_T3_WEST_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T3_WEST_B17_sel_value_O)
);
wire [16:0] RMUX_T4_EAST_B17_I [1:0];
assign RMUX_T4_EAST_B17_I[1] = REG_T4_EAST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T4_EAST_B17_I[0] = MUX_SB_T4_EAST_SB_OUT_B17_O;
wire [1:0] RMUX_T4_EAST_B17_valid_in;
assign RMUX_T4_EAST_B17_valid_in = {REG_T4_EAST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T4_EAST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T4_EAST_B17 (
    .I(RMUX_T4_EAST_B17_I),
    .O(RMUX_T4_EAST_B17_O),
    .ready_in(SB_T4_EAST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T4_EAST_B17_ready_out),
    .valid_in(RMUX_T4_EAST_B17_valid_in),
    .valid_out(RMUX_T4_EAST_B17_valid_out),
    .S(RMUX_T4_EAST_B17_sel_value_O),
    .out_sel(RMUX_T4_EAST_B17_out_sel)
);
SliceWrapper_32_12_13 RMUX_T4_EAST_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T4_EAST_B17_sel_value_O)
);
wire [16:0] RMUX_T4_NORTH_B17_I [1:0];
assign RMUX_T4_NORTH_B17_I[1] = REG_T4_NORTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T4_NORTH_B17_I[0] = MUX_SB_T4_NORTH_SB_OUT_B17_O;
wire [1:0] RMUX_T4_NORTH_B17_valid_in;
assign RMUX_T4_NORTH_B17_valid_in = {REG_T4_NORTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T4_NORTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T4_NORTH_B17 (
    .I(RMUX_T4_NORTH_B17_I),
    .O(RMUX_T4_NORTH_B17_O),
    .ready_in(SB_T4_NORTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T4_NORTH_B17_ready_out),
    .valid_in(RMUX_T4_NORTH_B17_valid_in),
    .valid_out(RMUX_T4_NORTH_B17_valid_out),
    .S(RMUX_T4_NORTH_B17_sel_value_O),
    .out_sel(RMUX_T4_NORTH_B17_out_sel)
);
SliceWrapper_32_13_14 RMUX_T4_NORTH_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T4_NORTH_B17_sel_value_O)
);
wire [16:0] RMUX_T4_SOUTH_B17_I [1:0];
assign RMUX_T4_SOUTH_B17_I[1] = REG_T4_SOUTH_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T4_SOUTH_B17_I[0] = MUX_SB_T4_SOUTH_SB_OUT_B17_O;
wire [1:0] RMUX_T4_SOUTH_B17_valid_in;
assign RMUX_T4_SOUTH_B17_valid_in = {REG_T4_SOUTH_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T4_SOUTH_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T4_SOUTH_B17 (
    .I(RMUX_T4_SOUTH_B17_I),
    .O(RMUX_T4_SOUTH_B17_O),
    .ready_in(SB_T4_SOUTH_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T4_SOUTH_B17_ready_out),
    .valid_in(RMUX_T4_SOUTH_B17_valid_in),
    .valid_out(RMUX_T4_SOUTH_B17_valid_out),
    .S(RMUX_T4_SOUTH_B17_sel_value_O),
    .out_sel(RMUX_T4_SOUTH_B17_out_sel)
);
SliceWrapper_32_14_15 RMUX_T4_SOUTH_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T4_SOUTH_B17_sel_value_O)
);
wire [16:0] RMUX_T4_WEST_B17_I [1:0];
assign RMUX_T4_WEST_B17_I[1] = REG_T4_WEST_B17$SplitFifo_17_inst0_data_out;
assign RMUX_T4_WEST_B17_I[0] = MUX_SB_T4_WEST_SB_OUT_B17_O;
wire [1:0] RMUX_T4_WEST_B17_valid_in;
assign RMUX_T4_WEST_B17_valid_in = {REG_T4_WEST_B17$SplitFifo_17_inst0_valid1[0],MUX_SB_T4_WEST_SB_OUT_B17_valid_out};
mux_aoi_ready_valid_2_17 RMUX_T4_WEST_B17 (
    .I(RMUX_T4_WEST_B17_I),
    .O(RMUX_T4_WEST_B17_O),
    .ready_in(SB_T4_WEST_SB_OUT_B17_ready_in),
    .ready_out(RMUX_T4_WEST_B17_ready_out),
    .valid_in(RMUX_T4_WEST_B17_valid_in),
    .valid_out(RMUX_T4_WEST_B17_valid_out),
    .S(RMUX_T4_WEST_B17_sel_value_O),
    .out_sel(RMUX_T4_WEST_B17_out_sel)
);
SliceWrapper_32_15_16 RMUX_T4_WEST_B17_sel_value (
    .I(config_reg_2_O),
    .O(RMUX_T4_WEST_B17_sel_value_O)
);
SliceWrapper_32_16_17 SB_T0_EAST_SB_IN_B17_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_EAST_SB_IN_B17_enable_value_O)
);
FanoutHash_302974B49BE3F0C4 SB_T0_EAST_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T0_WEST_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T0_EAST_SB_IN_B17_fan_in_O),
    .E1(SB_T3_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T0_EAST_SB_OUT_B17_FANOUT_I;
assign SB_T0_EAST_SB_OUT_B17_FANOUT_I = {REG_T0_EAST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T0_EAST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T0_EAST_SB_OUT_B17_FANOUT (
    .S(RMUX_T0_EAST_B17_out_sel),
    .O(SB_T0_EAST_SB_OUT_B17_FANOUT_O),
    .I(SB_T0_EAST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_32_17_18 SB_T0_EAST_SB_OUT_B17_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_EAST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_32_18_21 SB_T0_EAST_SB_OUT_B17_sel_value (
    .I(config_reg_2_O),
    .O(SB_T0_EAST_SB_OUT_B17_sel_value_O)
);
SliceWrapper_32_21_22 SB_T0_NORTH_SB_IN_B17_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_NORTH_SB_IN_B17_enable_value_O)
);
FanoutHash_47712AAC902ADA2 SB_T0_NORTH_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T0_WEST_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T0_NORTH_SB_IN_B17_fan_in_O),
    .E1(SB_T1_EAST_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T0_NORTH_SB_OUT_B17_FANOUT_I;
assign SB_T0_NORTH_SB_OUT_B17_FANOUT_I = {REG_T0_NORTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T0_NORTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T0_NORTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T0_NORTH_B17_out_sel),
    .O(SB_T0_NORTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T0_NORTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_32_22_23 SB_T0_NORTH_SB_OUT_B17_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_NORTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_32_23_26 SB_T0_NORTH_SB_OUT_B17_sel_value (
    .I(config_reg_2_O),
    .O(SB_T0_NORTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_32_26_27 SB_T0_SOUTH_SB_IN_B17_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_SOUTH_SB_IN_B17_enable_value_O)
);
FanoutHash_2785CE916183C5C SB_T0_SOUTH_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T1_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T3_EAST_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T0_SOUTH_SB_IN_B17_fan_in_O),
    .E1(SB_T0_NORTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T0_SOUTH_SB_OUT_B17_FANOUT_I;
assign SB_T0_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T0_SOUTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T0_SOUTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T0_SOUTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T0_SOUTH_B17_out_sel),
    .O(SB_T0_SOUTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T0_SOUTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_32_27_28 SB_T0_SOUTH_SB_OUT_B17_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_SOUTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_32_28_31 SB_T0_SOUTH_SB_OUT_B17_sel_value (
    .I(config_reg_2_O),
    .O(SB_T0_SOUTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_32_31_32 SB_T0_WEST_SB_IN_B17_enable_value (
    .I(config_reg_2_O),
    .O(SB_T0_WEST_SB_IN_B17_enable_value_O)
);
FanoutHash_65A468071775C7BB SB_T0_WEST_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T0_EAST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T0_WEST_SB_IN_B17_fan_in_O),
    .E1(SB_T4_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T0_WEST_SB_OUT_B17_FANOUT_I;
assign SB_T0_WEST_SB_OUT_B17_FANOUT_I = {REG_T0_WEST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T0_WEST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T0_WEST_SB_OUT_B17_FANOUT (
    .S(RMUX_T0_WEST_B17_out_sel),
    .O(SB_T0_WEST_SB_OUT_B17_FANOUT_O),
    .I(SB_T0_WEST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_31_0_1 SB_T0_WEST_SB_OUT_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T0_WEST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_31_1_4 SB_T0_WEST_SB_OUT_B17_sel_value (
    .I(config_reg_3_O),
    .O(SB_T0_WEST_SB_OUT_B17_sel_value_O)
);
SliceWrapper_31_4_5 SB_T1_EAST_SB_IN_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_EAST_SB_IN_B17_enable_value_O)
);
FanoutHash_4F83851A40824F89 SB_T1_EAST_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T2_SOUTH_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T0_NORTH_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T0_NORTH_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T0_NORTH_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T1_EAST_SB_IN_B17_fan_in_O),
    .E1(SB_T1_WEST_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T1_EAST_SB_OUT_B17_FANOUT_I;
assign SB_T1_EAST_SB_OUT_B17_FANOUT_I = {REG_T1_EAST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T1_EAST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T1_EAST_SB_OUT_B17_FANOUT (
    .S(RMUX_T1_EAST_B17_out_sel),
    .O(SB_T1_EAST_SB_OUT_B17_FANOUT_O),
    .I(SB_T1_EAST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_31_5_6 SB_T1_EAST_SB_OUT_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_EAST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_31_6_9 SB_T1_EAST_SB_OUT_B17_sel_value (
    .I(config_reg_3_O),
    .O(SB_T1_EAST_SB_OUT_B17_sel_value_O)
);
SliceWrapper_31_9_10 SB_T1_NORTH_SB_IN_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_NORTH_SB_IN_B17_enable_value_O)
);
FanoutHash_4FADDC8F90390680 SB_T1_NORTH_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T4_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T2_EAST_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T1_NORTH_SB_IN_B17_fan_in_O),
    .E1(SB_T1_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T1_NORTH_SB_OUT_B17_FANOUT_I;
assign SB_T1_NORTH_SB_OUT_B17_FANOUT_I = {REG_T1_NORTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T1_NORTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T1_NORTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T1_NORTH_B17_out_sel),
    .O(SB_T1_NORTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T1_NORTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_31_10_11 SB_T1_NORTH_SB_OUT_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_NORTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_31_11_14 SB_T1_NORTH_SB_OUT_B17_sel_value (
    .I(config_reg_3_O),
    .O(SB_T1_NORTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_31_14_15 SB_T1_SOUTH_SB_IN_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_SOUTH_SB_IN_B17_enable_value_O)
);
FanoutHash_466EB88CFD0CAD7B SB_T1_SOUTH_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T2_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T2_EAST_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T1_SOUTH_SB_IN_B17_fan_in_O),
    .E1(SB_T1_NORTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T1_SOUTH_SB_OUT_B17_FANOUT_I;
assign SB_T1_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T1_SOUTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T1_SOUTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T1_SOUTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T1_SOUTH_B17_out_sel),
    .O(SB_T1_SOUTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T1_SOUTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_31_15_16 SB_T1_SOUTH_SB_OUT_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_SOUTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_31_16_19 SB_T1_SOUTH_SB_OUT_B17_sel_value (
    .I(config_reg_3_O),
    .O(SB_T1_SOUTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_31_19_20 SB_T1_WEST_SB_IN_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_WEST_SB_IN_B17_enable_value_O)
);
FanoutHash_7ED1C80229B84786 SB_T1_WEST_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T1_EAST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T1_WEST_SB_IN_B17_fan_in_O),
    .E1(SB_T0_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T1_WEST_SB_OUT_B17_FANOUT_I;
assign SB_T1_WEST_SB_OUT_B17_FANOUT_I = {REG_T1_WEST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T1_WEST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T1_WEST_SB_OUT_B17_FANOUT (
    .S(RMUX_T1_WEST_B17_out_sel),
    .O(SB_T1_WEST_SB_OUT_B17_FANOUT_O),
    .I(SB_T1_WEST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_31_20_21 SB_T1_WEST_SB_OUT_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T1_WEST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_31_21_24 SB_T1_WEST_SB_OUT_B17_sel_value (
    .I(config_reg_3_O),
    .O(SB_T1_WEST_SB_OUT_B17_sel_value_O)
);
SliceWrapper_31_24_25 SB_T2_EAST_SB_IN_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T2_EAST_SB_IN_B17_enable_value_O)
);
FanoutHash_7F4660D1463D9234 SB_T2_EAST_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T2_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T2_EAST_SB_IN_B17_fan_in_O),
    .E1(SB_T1_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T2_EAST_SB_OUT_B17_FANOUT_I;
assign SB_T2_EAST_SB_OUT_B17_FANOUT_I = {REG_T2_EAST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T2_EAST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T2_EAST_SB_OUT_B17_FANOUT (
    .S(RMUX_T2_EAST_B17_out_sel),
    .O(SB_T2_EAST_SB_OUT_B17_FANOUT_O),
    .I(SB_T2_EAST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_31_25_26 SB_T2_EAST_SB_OUT_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T2_EAST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_31_26_29 SB_T2_EAST_SB_OUT_B17_sel_value (
    .I(config_reg_3_O),
    .O(SB_T2_EAST_SB_OUT_B17_sel_value_O)
);
SliceWrapper_31_29_30 SB_T2_NORTH_SB_IN_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T2_NORTH_SB_IN_B17_enable_value_O)
);
FanoutHash_3B67229CB02928BA SB_T2_NORTH_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T3_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T3_EAST_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T2_NORTH_SB_IN_B17_fan_in_O),
    .E1(SB_T2_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T2_NORTH_SB_OUT_B17_FANOUT_I;
assign SB_T2_NORTH_SB_OUT_B17_FANOUT_I = {REG_T2_NORTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T2_NORTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T2_NORTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T2_NORTH_B17_out_sel),
    .O(SB_T2_NORTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T2_NORTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_31_30_31 SB_T2_NORTH_SB_OUT_B17_enable_value (
    .I(config_reg_3_O),
    .O(SB_T2_NORTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_30_0_3 SB_T2_NORTH_SB_OUT_B17_sel_value (
    .I(config_reg_4_O),
    .O(SB_T2_NORTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_30_3_4 SB_T2_SOUTH_SB_IN_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T2_SOUTH_SB_IN_B17_enable_value_O)
);
FanoutHash_28125A548B305607 SB_T2_SOUTH_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T3_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T1_EAST_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T1_EAST_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T1_EAST_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T2_SOUTH_SB_IN_B17_fan_in_O),
    .E1(SB_T2_NORTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T2_SOUTH_SB_OUT_B17_FANOUT_I;
assign SB_T2_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T2_SOUTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T2_SOUTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T2_SOUTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T2_SOUTH_B17_out_sel),
    .O(SB_T2_SOUTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T2_SOUTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_30_4_5 SB_T2_SOUTH_SB_OUT_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T2_SOUTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_30_5_8 SB_T2_SOUTH_SB_OUT_B17_sel_value (
    .I(config_reg_4_O),
    .O(SB_T2_SOUTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_30_8_9 SB_T2_WEST_SB_IN_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T2_WEST_SB_IN_B17_enable_value_O)
);
FanoutHash_752C11B748DD905C SB_T2_WEST_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T2_EAST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T1_SOUTH_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T2_EAST_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T2_EAST_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T1_SOUTH_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T2_WEST_SB_IN_B17_fan_in_O),
    .E1(SB_T1_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T2_WEST_SB_OUT_B17_FANOUT_I;
assign SB_T2_WEST_SB_OUT_B17_FANOUT_I = {REG_T2_WEST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T2_WEST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T2_WEST_SB_OUT_B17_FANOUT (
    .S(RMUX_T2_WEST_B17_out_sel),
    .O(SB_T2_WEST_SB_OUT_B17_FANOUT_O),
    .I(SB_T2_WEST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_30_9_10 SB_T2_WEST_SB_OUT_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T2_WEST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_30_10_13 SB_T2_WEST_SB_OUT_B17_sel_value (
    .I(config_reg_4_O),
    .O(SB_T2_WEST_SB_OUT_B17_sel_value_O)
);
SliceWrapper_30_13_14 SB_T3_EAST_SB_IN_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_EAST_SB_IN_B17_enable_value_O)
);
FanoutHash_43D5C80ABD816837 SB_T3_EAST_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T3_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T0_SOUTH_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T3_WEST_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T3_WEST_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T0_SOUTH_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T0_SOUTH_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T3_EAST_SB_IN_B17_fan_in_O),
    .E1(SB_T2_NORTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T3_EAST_SB_OUT_B17_FANOUT_I;
assign SB_T3_EAST_SB_OUT_B17_FANOUT_I = {REG_T3_EAST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T3_EAST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T3_EAST_SB_OUT_B17_FANOUT (
    .S(RMUX_T3_EAST_B17_out_sel),
    .O(SB_T3_EAST_SB_OUT_B17_FANOUT_O),
    .I(SB_T3_EAST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_30_14_15 SB_T3_EAST_SB_OUT_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_EAST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_30_15_18 SB_T3_EAST_SB_OUT_B17_sel_value (
    .I(config_reg_4_O),
    .O(SB_T3_EAST_SB_OUT_B17_sel_value_O)
);
SliceWrapper_30_18_19 SB_T3_NORTH_SB_IN_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_NORTH_SB_IN_B17_enable_value_O)
);
FanoutHash_69376833A2418E2 SB_T3_NORTH_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T3_SOUTH_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T2_WEST_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T2_WEST_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T2_WEST_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T3_NORTH_SB_IN_B17_fan_in_O),
    .E1(SB_T4_EAST_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T3_NORTH_SB_OUT_B17_FANOUT_I;
assign SB_T3_NORTH_SB_OUT_B17_FANOUT_I = {REG_T3_NORTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T3_NORTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T3_NORTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T3_NORTH_B17_out_sel),
    .O(SB_T3_NORTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T3_NORTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_30_19_20 SB_T3_NORTH_SB_OUT_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_NORTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_30_20_23 SB_T3_NORTH_SB_OUT_B17_sel_value (
    .I(config_reg_4_O),
    .O(SB_T3_NORTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_30_23_24 SB_T3_SOUTH_SB_IN_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_SOUTH_SB_IN_B17_enable_value_O)
);
FanoutHash_66A75CC8494A4D6B SB_T3_SOUTH_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T4_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T0_EAST_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T3_SOUTH_SB_IN_B17_fan_in_O),
    .E1(SB_T3_NORTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T3_SOUTH_SB_OUT_B17_FANOUT_I;
assign SB_T3_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T3_SOUTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T3_SOUTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T3_SOUTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T3_SOUTH_B17_out_sel),
    .O(SB_T3_SOUTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T3_SOUTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_30_24_25 SB_T3_SOUTH_SB_OUT_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_SOUTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_30_25_28 SB_T3_SOUTH_SB_OUT_B17_sel_value (
    .I(config_reg_4_O),
    .O(SB_T3_SOUTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_30_28_29 SB_T3_WEST_SB_IN_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_WEST_SB_IN_B17_enable_value_O)
);
FanoutHash_31AE65CCDD94603 SB_T3_WEST_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T3_EAST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T2_SOUTH_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T2_NORTH_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T3_EAST_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T3_EAST_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T2_NORTH_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T2_NORTH_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T2_SOUTH_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T3_WEST_SB_IN_B17_fan_in_O),
    .E1(SB_T2_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T3_WEST_SB_OUT_B17_FANOUT_I;
assign SB_T3_WEST_SB_OUT_B17_FANOUT_I = {REG_T3_WEST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T3_WEST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T3_WEST_SB_OUT_B17_FANOUT (
    .S(RMUX_T3_WEST_B17_out_sel),
    .O(SB_T3_WEST_SB_OUT_B17_FANOUT_O),
    .I(SB_T3_WEST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_30_29_30 SB_T3_WEST_SB_OUT_B17_enable_value (
    .I(config_reg_4_O),
    .O(SB_T3_WEST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_23_0_3 SB_T3_WEST_SB_OUT_B17_sel_value (
    .I(config_reg_5_O),
    .O(SB_T3_WEST_SB_OUT_B17_sel_value_O)
);
SliceWrapper_23_3_4 SB_T4_EAST_SB_IN_B17_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_EAST_SB_IN_B17_enable_value_O)
);
FanoutHash_5D7AEC1255CDC1CC SB_T4_EAST_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T4_WEST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T3_NORTH_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T4_WEST_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T4_WEST_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T3_NORTH_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T3_NORTH_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T4_EAST_SB_IN_B17_fan_in_O),
    .E1(SB_T4_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T4_EAST_SB_OUT_B17_FANOUT_I;
assign SB_T4_EAST_SB_OUT_B17_FANOUT_I = {REG_T4_EAST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T4_EAST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T4_EAST_SB_OUT_B17_FANOUT (
    .S(RMUX_T4_EAST_B17_out_sel),
    .O(SB_T4_EAST_SB_OUT_B17_FANOUT_O),
    .I(SB_T4_EAST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_23_4_5 SB_T4_EAST_SB_OUT_B17_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_EAST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_23_5_8 SB_T4_EAST_SB_OUT_B17_sel_value (
    .I(config_reg_5_O),
    .O(SB_T4_EAST_SB_OUT_B17_sel_value_O)
);
SliceWrapper_23_8_9 SB_T4_NORTH_SB_IN_B17_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_NORTH_SB_IN_B17_enable_value_O)
);
FanoutHash_184DFC10DAF19BE9 SB_T4_NORTH_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T4_SOUTH_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T0_EAST_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T1_WEST_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T4_SOUTH_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T4_SOUTH_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T1_WEST_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T1_WEST_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T0_EAST_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T4_NORTH_SB_IN_B17_fan_in_O),
    .E1(SB_T0_EAST_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T4_NORTH_SB_OUT_B17_FANOUT_I;
assign SB_T4_NORTH_SB_OUT_B17_FANOUT_I = {REG_T4_NORTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T4_NORTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T4_NORTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T4_NORTH_B17_out_sel),
    .O(SB_T4_NORTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T4_NORTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_23_9_10 SB_T4_NORTH_SB_OUT_B17_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_NORTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_23_10_13 SB_T4_NORTH_SB_OUT_B17_sel_value (
    .I(config_reg_5_O),
    .O(SB_T4_NORTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_23_13_14 SB_T4_SOUTH_SB_IN_B17_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_SOUTH_SB_IN_B17_enable_value_O)
);
FanoutHash_26B6474864379B6A SB_T4_SOUTH_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T4_NORTH_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T0_WEST_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T4_NORTH_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T4_NORTH_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T0_WEST_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T0_WEST_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T4_SOUTH_SB_IN_B17_fan_in_O),
    .E1(SB_T4_EAST_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T4_SOUTH_SB_OUT_B17_FANOUT_I;
assign SB_T4_SOUTH_SB_OUT_B17_FANOUT_I = {REG_T4_SOUTH_B17$SplitFifo_17_inst0_ready0[0],RMUX_T4_SOUTH_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T4_SOUTH_SB_OUT_B17_FANOUT (
    .S(RMUX_T4_SOUTH_B17_out_sel),
    .O(SB_T4_SOUTH_SB_OUT_B17_FANOUT_O),
    .I(SB_T4_SOUTH_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_23_14_15 SB_T4_SOUTH_SB_OUT_B17_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_SOUTH_SB_OUT_B17_enable_value_O)
);
SliceWrapper_23_15_18 SB_T4_SOUTH_SB_OUT_B17_sel_value (
    .I(config_reg_5_O),
    .O(SB_T4_SOUTH_SB_OUT_B17_sel_value_O)
);
SliceWrapper_23_18_19 SB_T4_WEST_SB_IN_B17_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_WEST_SB_IN_B17_enable_value_O)
);
FanoutHash_1816466D6957000 SB_T4_WEST_SB_IN_B17_fan_in (
    .S6(MEM_input_width_17_num_3_out_sel),
    .E2(SB_T4_EAST_SB_OUT_B17_enable_value_O),
    .S1(MUX_SB_T3_SOUTH_SB_OUT_B17_out_sel),
    .I3(MEM_input_width_17_num_0_ready),
    .S0(MUX_SB_T1_NORTH_SB_OUT_B17_out_sel),
    .E5(MEM_input_width_17_num_2_enable),
    .I6(MEM_input_width_17_num_3_ready),
    .I2(MUX_SB_T4_EAST_SB_OUT_B17_ready_out),
    .S3(MEM_input_width_17_num_0_out_sel),
    .S2(MUX_SB_T4_EAST_SB_OUT_B17_out_sel),
    .E3(MEM_input_width_17_num_0_enable),
    .E0(SB_T1_NORTH_SB_OUT_B17_enable_value_O),
    .S4(MEM_input_width_17_num_1_out_sel),
    .I0(MUX_SB_T1_NORTH_SB_OUT_B17_ready_out),
    .E4(MEM_input_width_17_num_1_enable),
    .S5(MEM_input_width_17_num_2_out_sel),
    .I1(MUX_SB_T3_SOUTH_SB_OUT_B17_ready_out),
    .I5(MEM_input_width_17_num_2_ready),
    .E6(MEM_input_width_17_num_3_enable),
    .I4(MEM_input_width_17_num_1_ready),
    .O(SB_T4_WEST_SB_IN_B17_fan_in_O),
    .E1(SB_T3_SOUTH_SB_OUT_B17_enable_value_O)
);
wire [1:0] SB_T4_WEST_SB_OUT_B17_FANOUT_I;
assign SB_T4_WEST_SB_OUT_B17_FANOUT_I = {REG_T4_WEST_B17$SplitFifo_17_inst0_ready0[0],RMUX_T4_WEST_B17_ready_out};
ExclusiveNodeFanout_H2 SB_T4_WEST_SB_OUT_B17_FANOUT (
    .S(RMUX_T4_WEST_B17_out_sel),
    .O(SB_T4_WEST_SB_OUT_B17_FANOUT_O),
    .I(SB_T4_WEST_SB_OUT_B17_FANOUT_I)
);
SliceWrapper_23_19_20 SB_T4_WEST_SB_OUT_B17_enable_value (
    .I(config_reg_5_O),
    .O(SB_T4_WEST_SB_OUT_B17_enable_value_O)
);
SliceWrapper_23_20_23 SB_T4_WEST_SB_OUT_B17_sel_value (
    .I(config_reg_5_O),
    .O(SB_T4_WEST_SB_OUT_B17_sel_value_O)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T0_EAST_SB_IN_B17 (
    .I(SB_T0_EAST_SB_IN_B17),
    .O(WIRE_SB_T0_EAST_SB_IN_B17_O),
    .ready_in(SB_T0_EAST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T0_EAST_SB_IN_B17_ready_out),
    .valid_in(SB_T0_EAST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T0_EAST_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T0_NORTH_SB_IN_B17 (
    .I(SB_T0_NORTH_SB_IN_B17),
    .O(WIRE_SB_T0_NORTH_SB_IN_B17_O),
    .ready_in(SB_T0_NORTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T0_NORTH_SB_IN_B17_ready_out),
    .valid_in(SB_T0_NORTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T0_NORTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T0_SOUTH_SB_IN_B17 (
    .I(SB_T0_SOUTH_SB_IN_B17),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B17_O),
    .ready_in(SB_T0_SOUTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T0_SOUTH_SB_IN_B17_ready_out),
    .valid_in(SB_T0_SOUTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T0_SOUTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T0_WEST_SB_IN_B17 (
    .I(SB_T0_WEST_SB_IN_B17),
    .O(WIRE_SB_T0_WEST_SB_IN_B17_O),
    .ready_in(SB_T0_WEST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T0_WEST_SB_IN_B17_ready_out),
    .valid_in(SB_T0_WEST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T0_WEST_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T1_EAST_SB_IN_B17 (
    .I(SB_T1_EAST_SB_IN_B17),
    .O(WIRE_SB_T1_EAST_SB_IN_B17_O),
    .ready_in(SB_T1_EAST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T1_EAST_SB_IN_B17_ready_out),
    .valid_in(SB_T1_EAST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T1_EAST_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T1_NORTH_SB_IN_B17 (
    .I(SB_T1_NORTH_SB_IN_B17),
    .O(WIRE_SB_T1_NORTH_SB_IN_B17_O),
    .ready_in(SB_T1_NORTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T1_NORTH_SB_IN_B17_ready_out),
    .valid_in(SB_T1_NORTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T1_NORTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T1_SOUTH_SB_IN_B17 (
    .I(SB_T1_SOUTH_SB_IN_B17),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B17_O),
    .ready_in(SB_T1_SOUTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T1_SOUTH_SB_IN_B17_ready_out),
    .valid_in(SB_T1_SOUTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T1_SOUTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T1_WEST_SB_IN_B17 (
    .I(SB_T1_WEST_SB_IN_B17),
    .O(WIRE_SB_T1_WEST_SB_IN_B17_O),
    .ready_in(SB_T1_WEST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T1_WEST_SB_IN_B17_ready_out),
    .valid_in(SB_T1_WEST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T1_WEST_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T2_EAST_SB_IN_B17 (
    .I(SB_T2_EAST_SB_IN_B17),
    .O(WIRE_SB_T2_EAST_SB_IN_B17_O),
    .ready_in(SB_T2_EAST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T2_EAST_SB_IN_B17_ready_out),
    .valid_in(SB_T2_EAST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T2_EAST_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T2_NORTH_SB_IN_B17 (
    .I(SB_T2_NORTH_SB_IN_B17),
    .O(WIRE_SB_T2_NORTH_SB_IN_B17_O),
    .ready_in(SB_T2_NORTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T2_NORTH_SB_IN_B17_ready_out),
    .valid_in(SB_T2_NORTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T2_NORTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T2_SOUTH_SB_IN_B17 (
    .I(SB_T2_SOUTH_SB_IN_B17),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B17_O),
    .ready_in(SB_T2_SOUTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T2_SOUTH_SB_IN_B17_ready_out),
    .valid_in(SB_T2_SOUTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T2_SOUTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T2_WEST_SB_IN_B17 (
    .I(SB_T2_WEST_SB_IN_B17),
    .O(WIRE_SB_T2_WEST_SB_IN_B17_O),
    .ready_in(SB_T2_WEST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T2_WEST_SB_IN_B17_ready_out),
    .valid_in(SB_T2_WEST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T2_WEST_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T3_EAST_SB_IN_B17 (
    .I(SB_T3_EAST_SB_IN_B17),
    .O(WIRE_SB_T3_EAST_SB_IN_B17_O),
    .ready_in(SB_T3_EAST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T3_EAST_SB_IN_B17_ready_out),
    .valid_in(SB_T3_EAST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T3_EAST_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T3_NORTH_SB_IN_B17 (
    .I(SB_T3_NORTH_SB_IN_B17),
    .O(WIRE_SB_T3_NORTH_SB_IN_B17_O),
    .ready_in(SB_T3_NORTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T3_NORTH_SB_IN_B17_ready_out),
    .valid_in(SB_T3_NORTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T3_NORTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T3_SOUTH_SB_IN_B17 (
    .I(SB_T3_SOUTH_SB_IN_B17),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B17_O),
    .ready_in(SB_T3_SOUTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T3_SOUTH_SB_IN_B17_ready_out),
    .valid_in(SB_T3_SOUTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T3_SOUTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T3_WEST_SB_IN_B17 (
    .I(SB_T3_WEST_SB_IN_B17),
    .O(WIRE_SB_T3_WEST_SB_IN_B17_O),
    .ready_in(SB_T3_WEST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T3_WEST_SB_IN_B17_ready_out),
    .valid_in(SB_T3_WEST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T3_WEST_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T4_EAST_SB_IN_B17 (
    .I(SB_T4_EAST_SB_IN_B17),
    .O(WIRE_SB_T4_EAST_SB_IN_B17_O),
    .ready_in(SB_T4_EAST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T4_EAST_SB_IN_B17_ready_out),
    .valid_in(SB_T4_EAST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T4_EAST_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T4_NORTH_SB_IN_B17 (
    .I(SB_T4_NORTH_SB_IN_B17),
    .O(WIRE_SB_T4_NORTH_SB_IN_B17_O),
    .ready_in(SB_T4_NORTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T4_NORTH_SB_IN_B17_ready_out),
    .valid_in(SB_T4_NORTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T4_NORTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T4_SOUTH_SB_IN_B17 (
    .I(SB_T4_SOUTH_SB_IN_B17),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B17_O),
    .ready_in(SB_T4_SOUTH_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T4_SOUTH_SB_IN_B17_ready_out),
    .valid_in(SB_T4_SOUTH_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T4_SOUTH_SB_IN_B17_valid_out)
);
MuxWrapperAOI_1_17_RegularReadyValid WIRE_SB_T4_WEST_SB_IN_B17 (
    .I(SB_T4_WEST_SB_IN_B17),
    .O(WIRE_SB_T4_WEST_SB_IN_B17_O),
    .ready_in(SB_T4_WEST_SB_IN_B17_fan_in_O[0]),
    .ready_out(WIRE_SB_T4_WEST_SB_IN_B17_ready_out),
    .valid_in(SB_T4_WEST_SB_IN_B17_valid_in),
    .valid_out(WIRE_SB_T4_WEST_SB_IN_B17_valid_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_23_32_inst0$bit_const_0_None (
    .out(ZextWrapper_23_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_23_32_inst0$self_O_out;
assign ZextWrapper_23_32_inst0$self_O_out = {ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,config_reg_5_O};
mantle_wire__typeBitIn32 ZextWrapper_23_32_inst0$self_O (
    .in(ZextWrapper_23_32_inst0$self_O_in),
    .out(ZextWrapper_23_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_30_32_inst0$bit_const_0_None (
    .out(ZextWrapper_30_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_30_32_inst0$self_O_out;
assign ZextWrapper_30_32_inst0$self_O_out = {ZextWrapper_30_32_inst0$bit_const_0_None_out,ZextWrapper_30_32_inst0$bit_const_0_None_out,config_reg_4_O};
mantle_wire__typeBitIn32 ZextWrapper_30_32_inst0$self_O (
    .in(ZextWrapper_30_32_inst0$self_O_in),
    .out(ZextWrapper_30_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_31_32_inst0$bit_const_0_None (
    .out(ZextWrapper_31_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_31_32_inst0$self_O_out;
assign ZextWrapper_31_32_inst0$self_O_out = {ZextWrapper_31_32_inst0$bit_const_0_None_out,config_reg_3_O};
mantle_wire__typeBitIn32 ZextWrapper_31_32_inst0$self_O (
    .in(ZextWrapper_31_32_inst0$self_O_in),
    .out(ZextWrapper_31_32_inst0$self_O_out)
);
coreir_and #(
    .width(1)
) and1_inst0 (
    .in0(coreir_eq_1_inst0_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst0_out)
);
coreir_and #(
    .width(1)
) and1_inst1 (
    .in0(coreir_eq_1_inst1_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst1_out)
);
coreir_and #(
    .width(1)
) and1_inst10 (
    .in0(coreir_eq_1_inst10_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst10_out)
);
coreir_and #(
    .width(1)
) and1_inst11 (
    .in0(coreir_eq_1_inst11_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst11_out)
);
coreir_and #(
    .width(1)
) and1_inst12 (
    .in0(coreir_eq_1_inst12_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst12_out)
);
coreir_and #(
    .width(1)
) and1_inst13 (
    .in0(coreir_eq_1_inst13_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst13_out)
);
coreir_and #(
    .width(1)
) and1_inst14 (
    .in0(coreir_eq_1_inst14_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst14_out)
);
coreir_and #(
    .width(1)
) and1_inst15 (
    .in0(coreir_eq_1_inst15_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst15_out)
);
coreir_and #(
    .width(1)
) and1_inst16 (
    .in0(coreir_eq_1_inst16_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst16_out)
);
coreir_and #(
    .width(1)
) and1_inst17 (
    .in0(coreir_eq_1_inst17_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst17_out)
);
coreir_and #(
    .width(1)
) and1_inst18 (
    .in0(coreir_eq_1_inst18_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst18_out)
);
coreir_and #(
    .width(1)
) and1_inst19 (
    .in0(coreir_eq_1_inst19_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst19_out)
);
coreir_and #(
    .width(1)
) and1_inst2 (
    .in0(coreir_eq_1_inst2_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst2_out)
);
coreir_and #(
    .width(1)
) and1_inst3 (
    .in0(coreir_eq_1_inst3_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst3_out)
);
coreir_and #(
    .width(1)
) and1_inst4 (
    .in0(coreir_eq_1_inst4_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst4_out)
);
coreir_and #(
    .width(1)
) and1_inst5 (
    .in0(coreir_eq_1_inst5_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst5_out)
);
coreir_and #(
    .width(1)
) and1_inst6 (
    .in0(coreir_eq_1_inst6_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst6_out)
);
coreir_and #(
    .width(1)
) and1_inst7 (
    .in0(coreir_eq_1_inst7_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst7_out)
);
coreir_and #(
    .width(1)
) and1_inst8 (
    .in0(coreir_eq_1_inst8_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst8_out)
);
coreir_and #(
    .width(1)
) and1_inst9 (
    .in0(coreir_eq_1_inst9_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst9_out)
);
wire [7:0] config_reg_0_config_addr;
assign config_reg_0_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_32_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_reg_0_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_1_config_addr;
assign config_reg_1_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_32_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_reg_1_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_2_config_addr;
assign config_reg_2_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_32_8_32_2 config_reg_2 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_2_O),
    .config_addr(config_reg_2_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_3_config_addr;
assign config_reg_3_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_31_8_32_3 config_reg_3 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_3_O),
    .config_addr(config_reg_3_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_4_config_addr;
assign config_reg_4_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_30_8_32_4 config_reg_4 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_4_O),
    .config_addr(config_reg_4_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_5_config_addr;
assign config_reg_5_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_23_8_32_5 config_reg_5 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_5_O),
    .config_addr(config_reg_5_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst0 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_NORTH_B17_sel_value_O),
    .out(coreir_eq_1_inst0_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst1 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_SOUTH_B17_sel_value_O),
    .out(coreir_eq_1_inst1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst10 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_EAST_B17_sel_value_O),
    .out(coreir_eq_1_inst10_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst11 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_WEST_B17_sel_value_O),
    .out(coreir_eq_1_inst11_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst12 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_NORTH_B17_sel_value_O),
    .out(coreir_eq_1_inst12_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst13 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_SOUTH_B17_sel_value_O),
    .out(coreir_eq_1_inst13_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst14 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_EAST_B17_sel_value_O),
    .out(coreir_eq_1_inst14_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst15 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_WEST_B17_sel_value_O),
    .out(coreir_eq_1_inst15_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst16 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_NORTH_B17_sel_value_O),
    .out(coreir_eq_1_inst16_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst17 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_SOUTH_B17_sel_value_O),
    .out(coreir_eq_1_inst17_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst18 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_EAST_B17_sel_value_O),
    .out(coreir_eq_1_inst18_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst19 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_WEST_B17_sel_value_O),
    .out(coreir_eq_1_inst19_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst2 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_EAST_B17_sel_value_O),
    .out(coreir_eq_1_inst2_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst3 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_WEST_B17_sel_value_O),
    .out(coreir_eq_1_inst3_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst4 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_NORTH_B17_sel_value_O),
    .out(coreir_eq_1_inst4_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst5 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_SOUTH_B17_sel_value_O),
    .out(coreir_eq_1_inst5_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst6 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_EAST_B17_sel_value_O),
    .out(coreir_eq_1_inst6_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst7 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_WEST_B17_sel_value_O),
    .out(coreir_eq_1_inst7_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst8 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_NORTH_B17_sel_value_O),
    .out(coreir_eq_1_inst8_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst9 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_SOUTH_B17_sel_value_O),
    .out(coreir_eq_1_inst9_out)
);
wire [31:0] mux_aoi_6_32_inst0_I [5:0];
assign mux_aoi_6_32_inst0_I[5] = ZextWrapper_23_32_inst0$self_O_in;
assign mux_aoi_6_32_inst0_I[4] = ZextWrapper_30_32_inst0$self_O_in;
assign mux_aoi_6_32_inst0_I[3] = ZextWrapper_31_32_inst0$self_O_in;
assign mux_aoi_6_32_inst0_I[2] = config_reg_2_O;
assign mux_aoi_6_32_inst0_I[1] = config_reg_1_O;
assign mux_aoi_6_32_inst0_I[0] = config_reg_0_O;
mux_aoi_6_32 mux_aoi_6_32_inst0 (
    .I(mux_aoi_6_32_inst0_I),
    .O(mux_aoi_6_32_inst0_O),
    .S(self_config_config_addr_out[2:0]),
    .out_sel(mux_aoi_6_32_inst0_out_sel)
);
mantle_wire__typeBit8 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
assign MEM_output_width_17_num_0_ready_out = CB_MEM_output_width_17_num_0_fan_in_O[0];
assign MEM_output_width_17_num_1_ready_out = CB_MEM_output_width_17_num_1_fan_in_O[0];
assign MEM_output_width_17_num_2_ready_out = CB_MEM_output_width_17_num_2_fan_in_O[0];
assign SB_T0_EAST_SB_IN_B17_enable = SB_T0_EAST_SB_IN_B17_enable_value_O[0];
assign SB_T0_EAST_SB_IN_B17_ready_out = WIRE_SB_T0_EAST_SB_IN_B17_ready_out;
assign SB_T0_EAST_SB_OUT_B17 = RMUX_T0_EAST_B17_O;
assign SB_T0_EAST_SB_OUT_B17_enable = SB_T0_EAST_SB_OUT_B17_enable_value_O[0];
assign SB_T0_EAST_SB_OUT_B17_valid_out = RMUX_T0_EAST_B17_valid_out;
assign SB_T0_NORTH_SB_IN_B17_enable = SB_T0_NORTH_SB_IN_B17_enable_value_O[0];
assign SB_T0_NORTH_SB_IN_B17_ready_out = WIRE_SB_T0_NORTH_SB_IN_B17_ready_out;
assign SB_T0_NORTH_SB_OUT_B17 = RMUX_T0_NORTH_B17_O;
assign SB_T0_NORTH_SB_OUT_B17_enable = SB_T0_NORTH_SB_OUT_B17_enable_value_O[0];
assign SB_T0_NORTH_SB_OUT_B17_valid_out = RMUX_T0_NORTH_B17_valid_out;
assign SB_T0_SOUTH_SB_IN_B17_enable = SB_T0_SOUTH_SB_IN_B17_enable_value_O[0];
assign SB_T0_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T0_SOUTH_SB_IN_B17_ready_out;
assign SB_T0_SOUTH_SB_OUT_B17 = RMUX_T0_SOUTH_B17_O;
assign SB_T0_SOUTH_SB_OUT_B17_enable = SB_T0_SOUTH_SB_OUT_B17_enable_value_O[0];
assign SB_T0_SOUTH_SB_OUT_B17_valid_out = RMUX_T0_SOUTH_B17_valid_out;
assign SB_T0_WEST_SB_IN_B17_enable = SB_T0_WEST_SB_IN_B17_enable_value_O[0];
assign SB_T0_WEST_SB_IN_B17_ready_out = WIRE_SB_T0_WEST_SB_IN_B17_ready_out;
assign SB_T0_WEST_SB_OUT_B17 = RMUX_T0_WEST_B17_O;
assign SB_T0_WEST_SB_OUT_B17_enable = SB_T0_WEST_SB_OUT_B17_enable_value_O[0];
assign SB_T0_WEST_SB_OUT_B17_valid_out = RMUX_T0_WEST_B17_valid_out;
assign SB_T1_EAST_SB_IN_B17_enable = SB_T1_EAST_SB_IN_B17_enable_value_O[0];
assign SB_T1_EAST_SB_IN_B17_ready_out = WIRE_SB_T1_EAST_SB_IN_B17_ready_out;
assign SB_T1_EAST_SB_OUT_B17 = RMUX_T1_EAST_B17_O;
assign SB_T1_EAST_SB_OUT_B17_enable = SB_T1_EAST_SB_OUT_B17_enable_value_O[0];
assign SB_T1_EAST_SB_OUT_B17_valid_out = RMUX_T1_EAST_B17_valid_out;
assign SB_T1_NORTH_SB_IN_B17_enable = SB_T1_NORTH_SB_IN_B17_enable_value_O[0];
assign SB_T1_NORTH_SB_IN_B17_ready_out = WIRE_SB_T1_NORTH_SB_IN_B17_ready_out;
assign SB_T1_NORTH_SB_OUT_B17 = RMUX_T1_NORTH_B17_O;
assign SB_T1_NORTH_SB_OUT_B17_enable = SB_T1_NORTH_SB_OUT_B17_enable_value_O[0];
assign SB_T1_NORTH_SB_OUT_B17_valid_out = RMUX_T1_NORTH_B17_valid_out;
assign SB_T1_SOUTH_SB_IN_B17_enable = SB_T1_SOUTH_SB_IN_B17_enable_value_O[0];
assign SB_T1_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T1_SOUTH_SB_IN_B17_ready_out;
assign SB_T1_SOUTH_SB_OUT_B17 = RMUX_T1_SOUTH_B17_O;
assign SB_T1_SOUTH_SB_OUT_B17_enable = SB_T1_SOUTH_SB_OUT_B17_enable_value_O[0];
assign SB_T1_SOUTH_SB_OUT_B17_valid_out = RMUX_T1_SOUTH_B17_valid_out;
assign SB_T1_WEST_SB_IN_B17_enable = SB_T1_WEST_SB_IN_B17_enable_value_O[0];
assign SB_T1_WEST_SB_IN_B17_ready_out = WIRE_SB_T1_WEST_SB_IN_B17_ready_out;
assign SB_T1_WEST_SB_OUT_B17 = RMUX_T1_WEST_B17_O;
assign SB_T1_WEST_SB_OUT_B17_enable = SB_T1_WEST_SB_OUT_B17_enable_value_O[0];
assign SB_T1_WEST_SB_OUT_B17_valid_out = RMUX_T1_WEST_B17_valid_out;
assign SB_T2_EAST_SB_IN_B17_enable = SB_T2_EAST_SB_IN_B17_enable_value_O[0];
assign SB_T2_EAST_SB_IN_B17_ready_out = WIRE_SB_T2_EAST_SB_IN_B17_ready_out;
assign SB_T2_EAST_SB_OUT_B17 = RMUX_T2_EAST_B17_O;
assign SB_T2_EAST_SB_OUT_B17_enable = SB_T2_EAST_SB_OUT_B17_enable_value_O[0];
assign SB_T2_EAST_SB_OUT_B17_valid_out = RMUX_T2_EAST_B17_valid_out;
assign SB_T2_NORTH_SB_IN_B17_enable = SB_T2_NORTH_SB_IN_B17_enable_value_O[0];
assign SB_T2_NORTH_SB_IN_B17_ready_out = WIRE_SB_T2_NORTH_SB_IN_B17_ready_out;
assign SB_T2_NORTH_SB_OUT_B17 = RMUX_T2_NORTH_B17_O;
assign SB_T2_NORTH_SB_OUT_B17_enable = SB_T2_NORTH_SB_OUT_B17_enable_value_O[0];
assign SB_T2_NORTH_SB_OUT_B17_valid_out = RMUX_T2_NORTH_B17_valid_out;
assign SB_T2_SOUTH_SB_IN_B17_enable = SB_T2_SOUTH_SB_IN_B17_enable_value_O[0];
assign SB_T2_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T2_SOUTH_SB_IN_B17_ready_out;
assign SB_T2_SOUTH_SB_OUT_B17 = RMUX_T2_SOUTH_B17_O;
assign SB_T2_SOUTH_SB_OUT_B17_enable = SB_T2_SOUTH_SB_OUT_B17_enable_value_O[0];
assign SB_T2_SOUTH_SB_OUT_B17_valid_out = RMUX_T2_SOUTH_B17_valid_out;
assign SB_T2_WEST_SB_IN_B17_enable = SB_T2_WEST_SB_IN_B17_enable_value_O[0];
assign SB_T2_WEST_SB_IN_B17_ready_out = WIRE_SB_T2_WEST_SB_IN_B17_ready_out;
assign SB_T2_WEST_SB_OUT_B17 = RMUX_T2_WEST_B17_O;
assign SB_T2_WEST_SB_OUT_B17_enable = SB_T2_WEST_SB_OUT_B17_enable_value_O[0];
assign SB_T2_WEST_SB_OUT_B17_valid_out = RMUX_T2_WEST_B17_valid_out;
assign SB_T3_EAST_SB_IN_B17_enable = SB_T3_EAST_SB_IN_B17_enable_value_O[0];
assign SB_T3_EAST_SB_IN_B17_ready_out = WIRE_SB_T3_EAST_SB_IN_B17_ready_out;
assign SB_T3_EAST_SB_OUT_B17 = RMUX_T3_EAST_B17_O;
assign SB_T3_EAST_SB_OUT_B17_enable = SB_T3_EAST_SB_OUT_B17_enable_value_O[0];
assign SB_T3_EAST_SB_OUT_B17_valid_out = RMUX_T3_EAST_B17_valid_out;
assign SB_T3_NORTH_SB_IN_B17_enable = SB_T3_NORTH_SB_IN_B17_enable_value_O[0];
assign SB_T3_NORTH_SB_IN_B17_ready_out = WIRE_SB_T3_NORTH_SB_IN_B17_ready_out;
assign SB_T3_NORTH_SB_OUT_B17 = RMUX_T3_NORTH_B17_O;
assign SB_T3_NORTH_SB_OUT_B17_enable = SB_T3_NORTH_SB_OUT_B17_enable_value_O[0];
assign SB_T3_NORTH_SB_OUT_B17_valid_out = RMUX_T3_NORTH_B17_valid_out;
assign SB_T3_SOUTH_SB_IN_B17_enable = SB_T3_SOUTH_SB_IN_B17_enable_value_O[0];
assign SB_T3_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T3_SOUTH_SB_IN_B17_ready_out;
assign SB_T3_SOUTH_SB_OUT_B17 = RMUX_T3_SOUTH_B17_O;
assign SB_T3_SOUTH_SB_OUT_B17_enable = SB_T3_SOUTH_SB_OUT_B17_enable_value_O[0];
assign SB_T3_SOUTH_SB_OUT_B17_valid_out = RMUX_T3_SOUTH_B17_valid_out;
assign SB_T3_WEST_SB_IN_B17_enable = SB_T3_WEST_SB_IN_B17_enable_value_O[0];
assign SB_T3_WEST_SB_IN_B17_ready_out = WIRE_SB_T3_WEST_SB_IN_B17_ready_out;
assign SB_T3_WEST_SB_OUT_B17 = RMUX_T3_WEST_B17_O;
assign SB_T3_WEST_SB_OUT_B17_enable = SB_T3_WEST_SB_OUT_B17_enable_value_O[0];
assign SB_T3_WEST_SB_OUT_B17_valid_out = RMUX_T3_WEST_B17_valid_out;
assign SB_T4_EAST_SB_IN_B17_enable = SB_T4_EAST_SB_IN_B17_enable_value_O[0];
assign SB_T4_EAST_SB_IN_B17_ready_out = WIRE_SB_T4_EAST_SB_IN_B17_ready_out;
assign SB_T4_EAST_SB_OUT_B17 = RMUX_T4_EAST_B17_O;
assign SB_T4_EAST_SB_OUT_B17_enable = SB_T4_EAST_SB_OUT_B17_enable_value_O[0];
assign SB_T4_EAST_SB_OUT_B17_valid_out = RMUX_T4_EAST_B17_valid_out;
assign SB_T4_NORTH_SB_IN_B17_enable = SB_T4_NORTH_SB_IN_B17_enable_value_O[0];
assign SB_T4_NORTH_SB_IN_B17_ready_out = WIRE_SB_T4_NORTH_SB_IN_B17_ready_out;
assign SB_T4_NORTH_SB_OUT_B17 = RMUX_T4_NORTH_B17_O;
assign SB_T4_NORTH_SB_OUT_B17_enable = SB_T4_NORTH_SB_OUT_B17_enable_value_O[0];
assign SB_T4_NORTH_SB_OUT_B17_valid_out = RMUX_T4_NORTH_B17_valid_out;
assign SB_T4_SOUTH_SB_IN_B17_enable = SB_T4_SOUTH_SB_IN_B17_enable_value_O[0];
assign SB_T4_SOUTH_SB_IN_B17_ready_out = WIRE_SB_T4_SOUTH_SB_IN_B17_ready_out;
assign SB_T4_SOUTH_SB_OUT_B17 = RMUX_T4_SOUTH_B17_O;
assign SB_T4_SOUTH_SB_OUT_B17_enable = SB_T4_SOUTH_SB_OUT_B17_enable_value_O[0];
assign SB_T4_SOUTH_SB_OUT_B17_valid_out = RMUX_T4_SOUTH_B17_valid_out;
assign SB_T4_WEST_SB_IN_B17_enable = SB_T4_WEST_SB_IN_B17_enable_value_O[0];
assign SB_T4_WEST_SB_IN_B17_ready_out = WIRE_SB_T4_WEST_SB_IN_B17_ready_out;
assign SB_T4_WEST_SB_OUT_B17 = RMUX_T4_WEST_B17_O;
assign SB_T4_WEST_SB_OUT_B17_enable = SB_T4_WEST_SB_OUT_B17_enable_value_O[0];
assign SB_T4_WEST_SB_OUT_B17_valid_out = RMUX_T4_WEST_B17_valid_out;
assign read_config_data = mux_aoi_6_32_inst0_O;
endmodule

module ConfigRegister_20_8_32_3 (
    input clk,
    input reset,
    output [19:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [19:0] Register_inst0_O;
wire [7:0] const_3_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq1 Register_inst0 (
    .I(config_data[19:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h03),
    .width(8)
) const_3_8 (
    .out(const_3_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_3_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module PE (
    input [16:0] PE_input_width_17_num_0,
    output [0:0] PE_input_width_17_num_0_ready,
    input [0:0] PE_input_width_17_num_0_valid,
    input [16:0] PE_input_width_17_num_1,
    output [0:0] PE_input_width_17_num_1_ready,
    input [0:0] PE_input_width_17_num_1_valid,
    input [16:0] PE_input_width_17_num_2,
    output [0:0] PE_input_width_17_num_2_ready,
    input [0:0] PE_input_width_17_num_2_valid,
    input [16:0] PE_input_width_17_num_3,
    output [0:0] PE_input_width_17_num_3_ready,
    input [0:0] PE_input_width_17_num_3_valid,
    input [0:0] PE_input_width_1_num_0,
    output PE_input_width_1_num_0_ready,
    input PE_input_width_1_num_0_valid,
    input [0:0] PE_input_width_1_num_1,
    output PE_input_width_1_num_1_ready,
    input PE_input_width_1_num_1_valid,
    input [0:0] PE_input_width_1_num_2,
    output PE_input_width_1_num_2_ready,
    input PE_input_width_1_num_2_valid,
    output [16:0] PE_output_width_17_num_0,
    input [0:0] PE_output_width_17_num_0_ready,
    output [0:0] PE_output_width_17_num_0_valid,
    output [16:0] PE_output_width_17_num_1,
    input [0:0] PE_output_width_17_num_1_ready,
    output [0:0] PE_output_width_17_num_1_valid,
    output [16:0] PE_output_width_17_num_2,
    input [0:0] PE_output_width_17_num_2_ready,
    output [0:0] PE_output_width_17_num_2_valid,
    output [0:0] PE_output_width_1_num_0,
    input PE_output_width_1_num_0_ready,
    output PE_output_width_1_num_0_valid,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    input [0:0] flush,
    input [0:0] flush_core,
    output [31:0] read_config_data,
    input reset,
    input [0:0] stall
);
wire [31:0] CONFIG_SPACE_0_value_O;
wire [31:0] CONFIG_SPACE_1_value_O;
wire [21:0] CONFIG_SPACE_2_value_O;
wire [0:0] Invert1_inst0_out;
wire [0:0] Invert1_inst1_out;
wire [15:0] PE_inner_W_inst0_PE_onyx_inst_onyxpeintf_O3;
wire [15:0] PE_inner_W_inst0_PE_onyx_inst_onyxpeintf_O4;
wire [0:0] PE_inner_W_inst0_PE_input_width_17_num_0_ready;
wire [16:0] PE_inner_W_inst0_PE_output_width_17_num_2;
wire [15:0] PE_inner_W_inst0_PE_onyx_inst_onyxpeintf_O2;
wire [0:0] PE_inner_W_inst0_PE_input_width_17_num_3_ready;
wire [0:0] PE_inner_W_inst0_PE_output_width_1_num_0;
wire [0:0] PE_inner_W_inst0_PE_output_width_17_num_2_valid;
wire [16:0] PE_inner_W_inst0_PE_output_width_17_num_1;
wire [0:0] PE_inner_W_inst0_PE_input_width_17_num_2_ready;
wire [0:0] PE_inner_W_inst0_PE_input_width_17_num_1_ready;
wire [0:0] PE_inner_W_inst0_PE_output_width_17_num_1_valid;
wire [16:0] PE_inner_W_inst0_PE_output_width_17_num_0;
wire [0:0] PE_inner_W_inst0_PE_output_width_17_num_0_valid;
wire [0:0] PE_input_width_17_num_0_dense_value_O;
wire [0:0] PE_input_width_17_num_0_valid_reg_sel_value_O;
wire [0:0] PE_input_width_17_num_0_valid_reg_value_value_O;
wire [0:0] PE_input_width_17_num_0_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_input_width_17_num_1_dense_value_O;
wire [0:0] PE_input_width_17_num_1_valid_reg_sel_value_O;
wire [0:0] PE_input_width_17_num_1_valid_reg_value_value_O;
wire [0:0] PE_input_width_17_num_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_input_width_17_num_2_valid_reg_sel_value_O;
wire [0:0] PE_input_width_17_num_2_valid_reg_value_value_O;
wire [0:0] PE_input_width_17_num_2_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_input_width_17_num_3_valid_reg_sel_value_O;
wire [0:0] PE_input_width_17_num_3_valid_reg_value_value_O;
wire [0:0] PE_input_width_17_num_3_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_input_width_1_num_0_reg_sel_value_O;
wire [0:0] PE_input_width_1_num_0_reg_value_value_O;
wire [0:0] PE_input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_input_width_1_num_1_reg_sel_value_O;
wire [0:0] PE_input_width_1_num_1_reg_value_value_O;
wire [0:0] PE_input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_input_width_1_num_2_reg_sel_value_O;
wire [0:0] PE_input_width_1_num_2_reg_value_value_O;
wire [0:0] PE_input_width_1_num_2_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [15:0] PE_onyx_inst_onyxpeintf_O2_value_O;
wire [15:0] PE_onyx_inst_onyxpeintf_O3_value_O;
wire [15:0] PE_onyx_inst_onyxpeintf_O4_value_O;
wire [0:0] PE_output_width_17_num_0_dense_value_O;
wire [0:0] PE_output_width_17_num_0_ready_reg_sel_value_O;
wire [0:0] PE_output_width_17_num_0_ready_reg_value_value_O;
wire [0:0] PE_output_width_17_num_0_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_output_width_17_num_1_ready_reg_sel_value_O;
wire [0:0] PE_output_width_17_num_1_ready_reg_value_value_O;
wire [0:0] PE_output_width_17_num_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_output_width_17_num_2_ready_reg_sel_value_O;
wire [0:0] PE_output_width_17_num_2_ready_reg_value_value_O;
wire [0:0] PE_output_width_17_num_2_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire ZextWrapper_16_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_16_32_inst0$self_O_in;
wire ZextWrapper_16_32_inst1$bit_const_0_None_out;
wire [31:0] ZextWrapper_16_32_inst1$self_O_in;
wire ZextWrapper_16_32_inst2$bit_const_0_None_out;
wire [31:0] ZextWrapper_16_32_inst2$self_O_in;
wire ZextWrapper_20_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_20_32_inst0$self_O_in;
wire bit_const_1_None_out;
wire [31:0] config_reg_0_O;
wire [31:0] config_reg_1_O;
wire [31:0] config_reg_2_O;
wire [19:0] config_reg_3_O;
wire coreir_wrapInAsyncReset_inst0_out;
wire coreir_wrapOutAsyncReset_inst0_out;
wire [0:0] flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] flush_mux_sel_value_O;
wire [0:0] flush_reg_sel_value_O;
wire [0:0] flush_reg_value_value_O;
wire [0:0] flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [2:0] mode_value_O;
wire [31:0] mux_aoi_7_32_inst0_O;
wire [7:0] mux_aoi_7_32_inst0_out_sel;
wire [7:0] self_config_config_addr_out;
wire [0:0] tile_en_value_O;
SliceWrapper_32_0_32 CONFIG_SPACE_0_value (
    .I(config_reg_0_O),
    .O(CONFIG_SPACE_0_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_1_value (
    .I(config_reg_1_O),
    .O(CONFIG_SPACE_1_value_O)
);
SliceWrapper_32_0_22 CONFIG_SPACE_2_value (
    .I(config_reg_2_O),
    .O(CONFIG_SPACE_2_value_O)
);
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(coreir_wrapInAsyncReset_inst0_out),
    .out(Invert1_inst0_out)
);
coreir_not #(
    .width(1)
) Invert1_inst1 (
    .in(stall),
    .out(Invert1_inst1_out)
);
PE_inner_W PE_inner_W_inst0 (
    .PE_onyx_inst_onyxpeintf_O3(PE_inner_W_inst0_PE_onyx_inst_onyxpeintf_O3),
    .PE_onyx_inst_onyxpeintf_O4(PE_inner_W_inst0_PE_onyx_inst_onyxpeintf_O4),
    .rst_n(coreir_wrapOutAsyncReset_inst0_out),
    .PE_output_width_17_num_0_dense(PE_output_width_17_num_0_dense_value_O),
    .mode(mode_value_O),
    .PE_input_width_17_num_0_ready(PE_inner_W_inst0_PE_input_width_17_num_0_ready),
    .CONFIG_SPACE_1(CONFIG_SPACE_1_value_O),
    .PE_output_width_17_num_2_ready(PE_output_width_17_num_2_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .PE_output_width_17_num_2(PE_inner_W_inst0_PE_output_width_17_num_2),
    .PE_input_width_17_num_0(PE_input_width_17_num_0),
    .PE_input_width_17_num_2(PE_input_width_17_num_2),
    .PE_onyx_inst_onyxpeintf_O2(PE_inner_W_inst0_PE_onyx_inst_onyxpeintf_O2),
    .PE_input_width_17_num_1_valid(PE_input_width_17_num_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .PE_input_width_1_num_0(PE_input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .tile_en(tile_en_value_O),
    .clk(clk),
    .PE_input_width_17_num_0_valid(PE_input_width_17_num_0_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .PE_input_width_17_num_3(PE_input_width_17_num_3),
    .PE_input_width_17_num_3_ready(PE_inner_W_inst0_PE_input_width_17_num_3_ready),
    .PE_output_width_1_num_0(PE_inner_W_inst0_PE_output_width_1_num_0),
    .PE_output_width_17_num_2_valid(PE_inner_W_inst0_PE_output_width_17_num_2_valid),
    .PE_input_width_17_num_1(PE_input_width_17_num_1),
    .PE_output_width_17_num_1(PE_inner_W_inst0_PE_output_width_17_num_1),
    .PE_input_width_17_num_2_valid(PE_input_width_17_num_2_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .PE_input_width_17_num_2_ready(PE_inner_W_inst0_PE_input_width_17_num_2_ready),
    .PE_input_width_1_num_2(PE_input_width_1_num_2_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .clk_en(Invert1_inst1_out),
    .PE_output_width_17_num_0_ready(PE_output_width_17_num_0_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .CONFIG_SPACE_2(CONFIG_SPACE_2_value_O),
    .PE_input_width_17_num_1_dense(PE_input_width_17_num_1_dense_value_O),
    .PE_input_width_17_num_1_ready(PE_inner_W_inst0_PE_input_width_17_num_1_ready),
    .PE_output_width_17_num_1_ready(PE_output_width_17_num_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .PE_output_width_17_num_1_valid(PE_inner_W_inst0_PE_output_width_17_num_1_valid),
    .PE_input_width_1_num_1(PE_input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .PE_input_width_17_num_0_dense(PE_input_width_17_num_0_dense_value_O),
    .PE_output_width_17_num_0(PE_inner_W_inst0_PE_output_width_17_num_0),
    .flush(flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .CONFIG_SPACE_0(CONFIG_SPACE_0_value_O),
    .PE_output_width_17_num_0_valid(PE_inner_W_inst0_PE_output_width_17_num_0_valid),
    .PE_input_width_17_num_3_valid(PE_input_width_17_num_3_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_32_22_23 PE_input_width_17_num_0_dense_value (
    .I(config_reg_2_O),
    .O(PE_input_width_17_num_0_dense_value_O)
);
SliceWrapper_32_23_24 PE_input_width_17_num_0_valid_reg_sel_value (
    .I(config_reg_2_O),
    .O(PE_input_width_17_num_0_valid_reg_sel_value_O)
);
SliceWrapper_32_24_25 PE_input_width_17_num_0_valid_reg_value_value (
    .I(config_reg_2_O),
    .O(PE_input_width_17_num_0_valid_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) PE_input_width_17_num_0_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(PE_input_width_17_num_0_valid),
    .in1(PE_input_width_17_num_0_valid_reg_value_value_O),
    .sel(PE_input_width_17_num_0_valid_reg_sel_value_O[0]),
    .out(PE_input_width_17_num_0_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_32_25_26 PE_input_width_17_num_1_dense_value (
    .I(config_reg_2_O),
    .O(PE_input_width_17_num_1_dense_value_O)
);
SliceWrapper_32_26_27 PE_input_width_17_num_1_valid_reg_sel_value (
    .I(config_reg_2_O),
    .O(PE_input_width_17_num_1_valid_reg_sel_value_O)
);
SliceWrapper_32_27_28 PE_input_width_17_num_1_valid_reg_value_value (
    .I(config_reg_2_O),
    .O(PE_input_width_17_num_1_valid_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) PE_input_width_17_num_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(PE_input_width_17_num_1_valid),
    .in1(PE_input_width_17_num_1_valid_reg_value_value_O),
    .sel(PE_input_width_17_num_1_valid_reg_sel_value_O[0]),
    .out(PE_input_width_17_num_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_32_28_29 PE_input_width_17_num_2_valid_reg_sel_value (
    .I(config_reg_2_O),
    .O(PE_input_width_17_num_2_valid_reg_sel_value_O)
);
SliceWrapper_32_29_30 PE_input_width_17_num_2_valid_reg_value_value (
    .I(config_reg_2_O),
    .O(PE_input_width_17_num_2_valid_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) PE_input_width_17_num_2_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(PE_input_width_17_num_2_valid),
    .in1(PE_input_width_17_num_2_valid_reg_value_value_O),
    .sel(PE_input_width_17_num_2_valid_reg_sel_value_O[0]),
    .out(PE_input_width_17_num_2_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_32_30_31 PE_input_width_17_num_3_valid_reg_sel_value (
    .I(config_reg_2_O),
    .O(PE_input_width_17_num_3_valid_reg_sel_value_O)
);
SliceWrapper_32_31_32 PE_input_width_17_num_3_valid_reg_value_value (
    .I(config_reg_2_O),
    .O(PE_input_width_17_num_3_valid_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) PE_input_width_17_num_3_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(PE_input_width_17_num_3_valid),
    .in1(PE_input_width_17_num_3_valid_reg_value_value_O),
    .sel(PE_input_width_17_num_3_valid_reg_sel_value_O[0]),
    .out(PE_input_width_17_num_3_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_20_0_1 PE_input_width_1_num_0_reg_sel_value (
    .I(config_reg_3_O),
    .O(PE_input_width_1_num_0_reg_sel_value_O)
);
SliceWrapper_20_1_2 PE_input_width_1_num_0_reg_value_value (
    .I(config_reg_3_O),
    .O(PE_input_width_1_num_0_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) PE_input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(PE_input_width_1_num_0),
    .in1(PE_input_width_1_num_0_reg_value_value_O),
    .sel(PE_input_width_1_num_0_reg_sel_value_O[0]),
    .out(PE_input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_20_2_3 PE_input_width_1_num_1_reg_sel_value (
    .I(config_reg_3_O),
    .O(PE_input_width_1_num_1_reg_sel_value_O)
);
SliceWrapper_20_3_4 PE_input_width_1_num_1_reg_value_value (
    .I(config_reg_3_O),
    .O(PE_input_width_1_num_1_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) PE_input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(PE_input_width_1_num_1),
    .in1(PE_input_width_1_num_1_reg_value_value_O),
    .sel(PE_input_width_1_num_1_reg_sel_value_O[0]),
    .out(PE_input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_20_4_5 PE_input_width_1_num_2_reg_sel_value (
    .I(config_reg_3_O),
    .O(PE_input_width_1_num_2_reg_sel_value_O)
);
SliceWrapper_20_5_6 PE_input_width_1_num_2_reg_value_value (
    .I(config_reg_3_O),
    .O(PE_input_width_1_num_2_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) PE_input_width_1_num_2_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(PE_input_width_1_num_2),
    .in1(PE_input_width_1_num_2_reg_value_value_O),
    .sel(PE_input_width_1_num_2_reg_sel_value_O[0]),
    .out(PE_input_width_1_num_2_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_16_0_16 PE_onyx_inst_onyxpeintf_O2_value (
    .I(PE_inner_W_inst0_PE_onyx_inst_onyxpeintf_O2),
    .O(PE_onyx_inst_onyxpeintf_O2_value_O)
);
SliceWrapper_16_0_16 PE_onyx_inst_onyxpeintf_O3_value (
    .I(PE_inner_W_inst0_PE_onyx_inst_onyxpeintf_O3),
    .O(PE_onyx_inst_onyxpeintf_O3_value_O)
);
SliceWrapper_16_0_16 PE_onyx_inst_onyxpeintf_O4_value (
    .I(PE_inner_W_inst0_PE_onyx_inst_onyxpeintf_O4),
    .O(PE_onyx_inst_onyxpeintf_O4_value_O)
);
SliceWrapper_20_6_7 PE_output_width_17_num_0_dense_value (
    .I(config_reg_3_O),
    .O(PE_output_width_17_num_0_dense_value_O)
);
SliceWrapper_20_7_8 PE_output_width_17_num_0_ready_reg_sel_value (
    .I(config_reg_3_O),
    .O(PE_output_width_17_num_0_ready_reg_sel_value_O)
);
SliceWrapper_20_8_9 PE_output_width_17_num_0_ready_reg_value_value (
    .I(config_reg_3_O),
    .O(PE_output_width_17_num_0_ready_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) PE_output_width_17_num_0_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(PE_output_width_17_num_0_ready),
    .in1(PE_output_width_17_num_0_ready_reg_value_value_O),
    .sel(PE_output_width_17_num_0_ready_reg_sel_value_O[0]),
    .out(PE_output_width_17_num_0_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_20_9_10 PE_output_width_17_num_1_ready_reg_sel_value (
    .I(config_reg_3_O),
    .O(PE_output_width_17_num_1_ready_reg_sel_value_O)
);
SliceWrapper_20_10_11 PE_output_width_17_num_1_ready_reg_value_value (
    .I(config_reg_3_O),
    .O(PE_output_width_17_num_1_ready_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) PE_output_width_17_num_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(PE_output_width_17_num_1_ready),
    .in1(PE_output_width_17_num_1_ready_reg_value_value_O),
    .sel(PE_output_width_17_num_1_ready_reg_sel_value_O[0]),
    .out(PE_output_width_17_num_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_20_11_12 PE_output_width_17_num_2_ready_reg_sel_value (
    .I(config_reg_3_O),
    .O(PE_output_width_17_num_2_ready_reg_sel_value_O)
);
SliceWrapper_20_12_13 PE_output_width_17_num_2_ready_reg_value_value (
    .I(config_reg_3_O),
    .O(PE_output_width_17_num_2_ready_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) PE_output_width_17_num_2_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(PE_output_width_17_num_2_ready),
    .in1(PE_output_width_17_num_2_ready_reg_value_value_O),
    .sel(PE_output_width_17_num_2_ready_reg_sel_value_O[0]),
    .out(PE_output_width_17_num_2_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_16_32_inst0$bit_const_0_None (
    .out(ZextWrapper_16_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_16_32_inst0$self_O_out;
assign ZextWrapper_16_32_inst0$self_O_out = {ZextWrapper_16_32_inst0$bit_const_0_None_out,ZextWrapper_16_32_inst0$bit_const_0_None_out,ZextWrapper_16_32_inst0$bit_const_0_None_out,ZextWrapper_16_32_inst0$bit_const_0_None_out,ZextWrapper_16_32_inst0$bit_const_0_None_out,ZextWrapper_16_32_inst0$bit_const_0_None_out,ZextWrapper_16_32_inst0$bit_const_0_None_out,ZextWrapper_16_32_inst0$bit_const_0_None_out,ZextWrapper_16_32_inst0$bit_const_0_None_out,ZextWrapper_16_32_inst0$bit_const_0_None_out,ZextWrapper_16_32_inst0$bit_const_0_None_out,ZextWrapper_16_32_inst0$bit_const_0_None_out,ZextWrapper_16_32_inst0$bit_const_0_None_out,ZextWrapper_16_32_inst0$bit_const_0_None_out,ZextWrapper_16_32_inst0$bit_const_0_None_out,ZextWrapper_16_32_inst0$bit_const_0_None_out,PE_onyx_inst_onyxpeintf_O3_value_O};
mantle_wire__typeBitIn32 ZextWrapper_16_32_inst0$self_O (
    .in(ZextWrapper_16_32_inst0$self_O_in),
    .out(ZextWrapper_16_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_16_32_inst1$bit_const_0_None (
    .out(ZextWrapper_16_32_inst1$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_16_32_inst1$self_O_out;
assign ZextWrapper_16_32_inst1$self_O_out = {ZextWrapper_16_32_inst1$bit_const_0_None_out,ZextWrapper_16_32_inst1$bit_const_0_None_out,ZextWrapper_16_32_inst1$bit_const_0_None_out,ZextWrapper_16_32_inst1$bit_const_0_None_out,ZextWrapper_16_32_inst1$bit_const_0_None_out,ZextWrapper_16_32_inst1$bit_const_0_None_out,ZextWrapper_16_32_inst1$bit_const_0_None_out,ZextWrapper_16_32_inst1$bit_const_0_None_out,ZextWrapper_16_32_inst1$bit_const_0_None_out,ZextWrapper_16_32_inst1$bit_const_0_None_out,ZextWrapper_16_32_inst1$bit_const_0_None_out,ZextWrapper_16_32_inst1$bit_const_0_None_out,ZextWrapper_16_32_inst1$bit_const_0_None_out,ZextWrapper_16_32_inst1$bit_const_0_None_out,ZextWrapper_16_32_inst1$bit_const_0_None_out,ZextWrapper_16_32_inst1$bit_const_0_None_out,PE_onyx_inst_onyxpeintf_O4_value_O};
mantle_wire__typeBitIn32 ZextWrapper_16_32_inst1$self_O (
    .in(ZextWrapper_16_32_inst1$self_O_in),
    .out(ZextWrapper_16_32_inst1$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_16_32_inst2$bit_const_0_None (
    .out(ZextWrapper_16_32_inst2$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_16_32_inst2$self_O_out;
assign ZextWrapper_16_32_inst2$self_O_out = {ZextWrapper_16_32_inst2$bit_const_0_None_out,ZextWrapper_16_32_inst2$bit_const_0_None_out,ZextWrapper_16_32_inst2$bit_const_0_None_out,ZextWrapper_16_32_inst2$bit_const_0_None_out,ZextWrapper_16_32_inst2$bit_const_0_None_out,ZextWrapper_16_32_inst2$bit_const_0_None_out,ZextWrapper_16_32_inst2$bit_const_0_None_out,ZextWrapper_16_32_inst2$bit_const_0_None_out,ZextWrapper_16_32_inst2$bit_const_0_None_out,ZextWrapper_16_32_inst2$bit_const_0_None_out,ZextWrapper_16_32_inst2$bit_const_0_None_out,ZextWrapper_16_32_inst2$bit_const_0_None_out,ZextWrapper_16_32_inst2$bit_const_0_None_out,ZextWrapper_16_32_inst2$bit_const_0_None_out,ZextWrapper_16_32_inst2$bit_const_0_None_out,ZextWrapper_16_32_inst2$bit_const_0_None_out,PE_onyx_inst_onyxpeintf_O2_value_O};
mantle_wire__typeBitIn32 ZextWrapper_16_32_inst2$self_O (
    .in(ZextWrapper_16_32_inst2$self_O_in),
    .out(ZextWrapper_16_32_inst2$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_20_32_inst0$bit_const_0_None (
    .out(ZextWrapper_20_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_20_32_inst0$self_O_out;
assign ZextWrapper_20_32_inst0$self_O_out = {ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,config_reg_3_O};
mantle_wire__typeBitIn32 ZextWrapper_20_32_inst0$self_O (
    .in(ZextWrapper_20_32_inst0$self_O_in),
    .out(ZextWrapper_20_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b1)
) bit_const_1_None (
    .out(bit_const_1_None_out)
);
wire [7:0] config_reg_0_config_addr;
assign config_reg_0_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_32_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_reg_0_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_1_config_addr;
assign config_reg_1_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_32_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_reg_1_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_2_config_addr;
assign config_reg_2_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_32_8_32_2 config_reg_2 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_2_O),
    .config_addr(config_reg_2_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_3_config_addr;
assign config_reg_3_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4],self_config_config_addr_out[3],self_config_config_addr_out[2:0]};
ConfigRegister_20_8_32_3 config_reg_3 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_3_O),
    .config_addr(config_reg_3_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_wrap coreir_wrapInAsyncReset_inst0 (
    .in(reset),
    .out(coreir_wrapInAsyncReset_inst0_out)
);
coreir_wrap coreir_wrapOutAsyncReset_inst0 (
    .in(Invert1_inst0_out[0]),
    .out(coreir_wrapOutAsyncReset_inst0_out)
);
coreir_mux #(
    .width(1)
) flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(flush_core),
    .in1(flush),
    .sel(flush_mux_sel_value_O[0]),
    .out(flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_20_13_14 flush_mux_sel_value (
    .I(config_reg_3_O),
    .O(flush_mux_sel_value_O)
);
SliceWrapper_20_14_15 flush_reg_sel_value (
    .I(config_reg_3_O),
    .O(flush_reg_sel_value_O)
);
SliceWrapper_20_15_16 flush_reg_value_value (
    .I(config_reg_3_O),
    .O(flush_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(flush),
    .in1(flush_reg_value_value_O),
    .sel(flush_reg_sel_value_O[0]),
    .out(flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_20_16_19 mode_value (
    .I(config_reg_3_O),
    .O(mode_value_O)
);
wire [31:0] mux_aoi_7_32_inst0_I [6:0];
assign mux_aoi_7_32_inst0_I[6] = ZextWrapper_16_32_inst2$self_O_in;
assign mux_aoi_7_32_inst0_I[5] = ZextWrapper_16_32_inst1$self_O_in;
assign mux_aoi_7_32_inst0_I[4] = ZextWrapper_16_32_inst0$self_O_in;
assign mux_aoi_7_32_inst0_I[3] = ZextWrapper_20_32_inst0$self_O_in;
assign mux_aoi_7_32_inst0_I[2] = config_reg_2_O;
assign mux_aoi_7_32_inst0_I[1] = config_reg_1_O;
assign mux_aoi_7_32_inst0_I[0] = config_reg_0_O;
mux_aoi_7_32 mux_aoi_7_32_inst0 (
    .I(mux_aoi_7_32_inst0_I),
    .O(mux_aoi_7_32_inst0_O),
    .S(self_config_config_addr_out[2:0]),
    .out_sel(mux_aoi_7_32_inst0_out_sel)
);
mantle_wire__typeBit8 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
SliceWrapper_20_19_20 tile_en_value (
    .I(config_reg_3_O),
    .O(tile_en_value_O)
);
assign PE_input_width_17_num_0_ready = PE_inner_W_inst0_PE_input_width_17_num_0_ready;
assign PE_input_width_17_num_1_ready = PE_inner_W_inst0_PE_input_width_17_num_1_ready;
assign PE_input_width_17_num_2_ready = PE_inner_W_inst0_PE_input_width_17_num_2_ready;
assign PE_input_width_17_num_3_ready = PE_inner_W_inst0_PE_input_width_17_num_3_ready;
assign PE_input_width_1_num_0_ready = bit_const_1_None_out;
assign PE_input_width_1_num_1_ready = bit_const_1_None_out;
assign PE_input_width_1_num_2_ready = bit_const_1_None_out;
assign PE_output_width_17_num_0 = PE_inner_W_inst0_PE_output_width_17_num_0;
assign PE_output_width_17_num_0_valid = PE_inner_W_inst0_PE_output_width_17_num_0_valid;
assign PE_output_width_17_num_1 = PE_inner_W_inst0_PE_output_width_17_num_1;
assign PE_output_width_17_num_1_valid = PE_inner_W_inst0_PE_output_width_17_num_1_valid;
assign PE_output_width_17_num_2 = PE_inner_W_inst0_PE_output_width_17_num_2;
assign PE_output_width_17_num_2_valid = PE_inner_W_inst0_PE_output_width_17_num_2_valid;
assign PE_output_width_1_num_0 = PE_inner_W_inst0_PE_output_width_1_num_0;
assign PE_output_width_1_num_0_valid = bit_const_1_None_out;
assign read_config_data = mux_aoi_7_32_inst0_O;
endmodule

module ConfigRegister_1_8_32_17 (
    input clk,
    input reset,
    output [0:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [0:0] Register_inst0_O;
wire [7:0] const_17_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq4 Register_inst0 (
    .I(config_data[0:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h11),
    .width(8)
) const_17_8 (
    .out(const_17_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_17_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module PondCore (
    input [16:0] PondTop_input_width_17_num_0,
    output PondTop_input_width_17_num_0_ready,
    input PondTop_input_width_17_num_0_valid,
    input [16:0] PondTop_input_width_17_num_1,
    output PondTop_input_width_17_num_1_ready,
    input PondTop_input_width_17_num_1_valid,
    output [16:0] PondTop_output_width_17_num_0,
    input PondTop_output_width_17_num_0_ready,
    output PondTop_output_width_17_num_0_valid,
    output [16:0] PondTop_output_width_17_num_1,
    input PondTop_output_width_17_num_1_ready,
    output PondTop_output_width_17_num_1_valid,
    output [0:0] PondTop_output_width_1_num_0,
    input PondTop_output_width_1_num_0_ready,
    output PondTop_output_width_1_num_0_valid,
    output [0:0] PondTop_output_width_1_num_1,
    input PondTop_output_width_1_num_1_ready,
    output PondTop_output_width_1_num_1_valid,
    input clk,
    input [7:0] config_1_config_addr,
    input [31:0] config_1_config_data,
    input [0:0] config_1_read,
    input [0:0] config_1_write,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input config_en_0,
    input [0:0] config_read,
    input [0:0] config_write,
    input [0:0] flush,
    input [0:0] flush_core,
    output [31:0] read_config_data,
    output [31:0] read_config_data_1,
    input reset,
    input [0:0] stall
);
wire [0:0] AND_CONFIG_EN_SRAM_0_out;
wire [31:0] CONFIG_SPACE_0_value_O;
wire [31:0] CONFIG_SPACE_10_value_O;
wire [31:0] CONFIG_SPACE_11_value_O;
wire [31:0] CONFIG_SPACE_12_value_O;
wire [31:0] CONFIG_SPACE_13_value_O;
wire [31:0] CONFIG_SPACE_14_value_O;
wire [31:0] CONFIG_SPACE_15_value_O;
wire [29:0] CONFIG_SPACE_16_value_O;
wire [31:0] CONFIG_SPACE_1_value_O;
wire [31:0] CONFIG_SPACE_2_value_O;
wire [31:0] CONFIG_SPACE_3_value_O;
wire [31:0] CONFIG_SPACE_4_value_O;
wire [31:0] CONFIG_SPACE_5_value_O;
wire [31:0] CONFIG_SPACE_6_value_O;
wire [31:0] CONFIG_SPACE_7_value_O;
wire [31:0] CONFIG_SPACE_8_value_O;
wire [31:0] CONFIG_SPACE_9_value_O;
wire [0:0] Invert1_inst0_out;
wire [0:0] Invert1_inst1_out;
wire [0:0] OR_CONFIG_EN_SRAM_0_out;
wire OR_CONFIG_RD_SRAM$orr_inst0_out;
wire OR_CONFIG_WR_SRAM$orr_inst0_out;
wire [7:0] OR_config_addr_FEATURE_out;
wire [31:0] OR_config_data_FEATURE_out;
wire [16:0] PondTop_W_inst0_PondTop_output_width_17_num_1;
wire [0:0] PondTop_W_inst0_PondTop_output_width_1_num_1;
wire [31:0] PondTop_W_inst0_config_data_out;
wire [0:0] PondTop_W_inst0_PondTop_output_width_1_num_0;
wire [16:0] PondTop_W_inst0_PondTop_output_width_17_num_0;
wire ZextWrapper_1_32_inst0$bit_const_0_None_out;
wire ZextWrapper_30_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_30_32_inst0$self_O_in;
wire bit_const_1_None_out;
wire [31:0] config_reg_0_O;
wire [31:0] config_reg_1_O;
wire [31:0] config_reg_10_O;
wire [31:0] config_reg_11_O;
wire [31:0] config_reg_12_O;
wire [31:0] config_reg_13_O;
wire [31:0] config_reg_14_O;
wire [31:0] config_reg_15_O;
wire [31:0] config_reg_16_O;
wire [0:0] config_reg_17_O;
wire [31:0] config_reg_2_O;
wire [31:0] config_reg_3_O;
wire [31:0] config_reg_4_O;
wire [31:0] config_reg_5_O;
wire [31:0] config_reg_6_O;
wire [31:0] config_reg_7_O;
wire [29:0] config_reg_8_O;
wire [31:0] config_reg_9_O;
wire coreir_wrapInAsyncReset_inst0_out;
wire coreir_wrapOutAsyncReset_inst0_out;
wire [31:0] mux_aoi_18_32_inst0_O;
wire [31:0] mux_aoi_18_32_inst0_out_sel;
wire [0:0] or1_inst0_out;
wire [7:0] self_config_config_addr_out;
wire [0:0] tile_en_value_O;
coreir_and #(
    .width(1)
) AND_CONFIG_EN_SRAM_0 (
    .in0(OR_CONFIG_EN_SRAM_0_out),
    .in1(config_en_0),
    .out(AND_CONFIG_EN_SRAM_0_out)
);
SliceWrapper_32_0_32 CONFIG_SPACE_0_value (
    .I(config_reg_0_O),
    .O(CONFIG_SPACE_0_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_10_value (
    .I(config_reg_2_O),
    .O(CONFIG_SPACE_10_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_11_value (
    .I(config_reg_3_O),
    .O(CONFIG_SPACE_11_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_12_value (
    .I(config_reg_4_O),
    .O(CONFIG_SPACE_12_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_13_value (
    .I(config_reg_5_O),
    .O(CONFIG_SPACE_13_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_14_value (
    .I(config_reg_6_O),
    .O(CONFIG_SPACE_14_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_15_value (
    .I(config_reg_7_O),
    .O(CONFIG_SPACE_15_value_O)
);
SliceWrapper_30_0_30 CONFIG_SPACE_16_value (
    .I(config_reg_8_O),
    .O(CONFIG_SPACE_16_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_1_value (
    .I(config_reg_1_O),
    .O(CONFIG_SPACE_1_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_2_value (
    .I(config_reg_9_O),
    .O(CONFIG_SPACE_2_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_3_value (
    .I(config_reg_10_O),
    .O(CONFIG_SPACE_3_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_4_value (
    .I(config_reg_11_O),
    .O(CONFIG_SPACE_4_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_5_value (
    .I(config_reg_12_O),
    .O(CONFIG_SPACE_5_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_6_value (
    .I(config_reg_13_O),
    .O(CONFIG_SPACE_6_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_7_value (
    .I(config_reg_14_O),
    .O(CONFIG_SPACE_7_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_8_value (
    .I(config_reg_15_O),
    .O(CONFIG_SPACE_8_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_9_value (
    .I(config_reg_16_O),
    .O(CONFIG_SPACE_9_value_O)
);
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(coreir_wrapInAsyncReset_inst0_out),
    .out(Invert1_inst0_out)
);
coreir_not #(
    .width(1)
) Invert1_inst1 (
    .in(stall),
    .out(Invert1_inst1_out)
);
coreir_or #(
    .width(1)
) OR_CONFIG_EN_SRAM_0 (
    .in0(config_1_write),
    .in1(config_1_read),
    .out(OR_CONFIG_EN_SRAM_0_out)
);
coreir_orr #(
    .width(1)
) OR_CONFIG_RD_SRAM$orr_inst0 (
    .in(config_1_write),
    .out(OR_CONFIG_RD_SRAM$orr_inst0_out)
);
coreir_orr #(
    .width(1)
) OR_CONFIG_WR_SRAM$orr_inst0 (
    .in(config_1_read),
    .out(OR_CONFIG_WR_SRAM$orr_inst0_out)
);
wire [7:0] OR_config_addr_FEATURE_in0;
assign OR_config_addr_FEATURE_in0 = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
coreir_or #(
    .width(8)
) OR_config_addr_FEATURE (
    .in0(OR_config_addr_FEATURE_in0),
    .in1(config_1_config_addr),
    .out(OR_config_addr_FEATURE_out)
);
coreir_or #(
    .width(32)
) OR_config_data_FEATURE (
    .in0(config_config_data),
    .in1(config_1_config_data),
    .out(OR_config_data_FEATURE_out)
);
PondTop_W PondTop_W_inst0 (
    .PondTop_output_width_17_num_1(PondTop_W_inst0_PondTop_output_width_17_num_1),
    .CONFIG_SPACE_5(CONFIG_SPACE_5_value_O),
    .config_data_in(OR_config_data_FEATURE_out),
    .config_en(AND_CONFIG_EN_SRAM_0_out),
    .PondTop_output_width_1_num_1(PondTop_W_inst0_PondTop_output_width_1_num_1),
    .CONFIG_SPACE_10(CONFIG_SPACE_10_value_O),
    .rst_n(coreir_wrapOutAsyncReset_inst0_out),
    .CONFIG_SPACE_11(CONFIG_SPACE_11_value_O),
    .CONFIG_SPACE_6(CONFIG_SPACE_6_value_O),
    .CONFIG_SPACE_15(CONFIG_SPACE_15_value_O),
    .config_data_out(PondTop_W_inst0_config_data_out),
    .CONFIG_SPACE_14(CONFIG_SPACE_14_value_O),
    .config_addr_in(OR_config_addr_FEATURE_out),
    .CONFIG_SPACE_1(CONFIG_SPACE_1_value_O),
    .CONFIG_SPACE_3(CONFIG_SPACE_3_value_O),
    .CONFIG_SPACE_13(CONFIG_SPACE_13_value_O),
    .CONFIG_SPACE_7(CONFIG_SPACE_7_value_O),
    .tile_en(tile_en_value_O),
    .config_read(OR_CONFIG_WR_SRAM$orr_inst0_out),
    .clk(clk),
    .CONFIG_SPACE_4(CONFIG_SPACE_4_value_O),
    .CONFIG_SPACE_9(CONFIG_SPACE_9_value_O),
    .CONFIG_SPACE_16(CONFIG_SPACE_16_value_O),
    .config_write(OR_CONFIG_RD_SRAM$orr_inst0_out),
    .PondTop_output_width_1_num_0(PondTop_W_inst0_PondTop_output_width_1_num_0),
    .PondTop_input_width_17_num_0(PondTop_input_width_17_num_0),
    .CONFIG_SPACE_12(CONFIG_SPACE_12_value_O),
    .clk_en(Invert1_inst1_out),
    .CONFIG_SPACE_2(CONFIG_SPACE_2_value_O),
    .PondTop_input_width_17_num_1(PondTop_input_width_17_num_1),
    .flush(or1_inst0_out),
    .PondTop_output_width_17_num_0(PondTop_W_inst0_PondTop_output_width_17_num_0),
    .CONFIG_SPACE_0(CONFIG_SPACE_0_value_O),
    .CONFIG_SPACE_8(CONFIG_SPACE_8_value_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_1_32_inst0$bit_const_0_None (
    .out(ZextWrapper_1_32_inst0$bit_const_0_None_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_30_32_inst0$bit_const_0_None (
    .out(ZextWrapper_30_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_30_32_inst0$self_O_out;
assign ZextWrapper_30_32_inst0$self_O_out = {ZextWrapper_30_32_inst0$bit_const_0_None_out,ZextWrapper_30_32_inst0$bit_const_0_None_out,config_reg_8_O};
mantle_wire__typeBitIn32 ZextWrapper_30_32_inst0$self_O (
    .in(ZextWrapper_30_32_inst0$self_O_in),
    .out(ZextWrapper_30_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b1)
) bit_const_1_None (
    .out(bit_const_1_None_out)
);
wire [7:0] config_reg_0_config_addr;
assign config_reg_0_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
ConfigRegister_32_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_reg_0_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_1_config_addr;
assign config_reg_1_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
ConfigRegister_32_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_reg_1_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_10_config_addr;
assign config_reg_10_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
ConfigRegister_32_8_32_10 config_reg_10 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_10_O),
    .config_addr(config_reg_10_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_11_config_addr;
assign config_reg_11_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
ConfigRegister_32_8_32_11 config_reg_11 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_11_O),
    .config_addr(config_reg_11_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_12_config_addr;
assign config_reg_12_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
ConfigRegister_32_8_32_12 config_reg_12 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_12_O),
    .config_addr(config_reg_12_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_13_config_addr;
assign config_reg_13_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
ConfigRegister_32_8_32_13 config_reg_13 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_13_O),
    .config_addr(config_reg_13_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_14_config_addr;
assign config_reg_14_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
ConfigRegister_32_8_32_14 config_reg_14 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_14_O),
    .config_addr(config_reg_14_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_15_config_addr;
assign config_reg_15_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
ConfigRegister_32_8_32_15 config_reg_15 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_15_O),
    .config_addr(config_reg_15_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_16_config_addr;
assign config_reg_16_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
ConfigRegister_32_8_32_16 config_reg_16 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_16_O),
    .config_addr(config_reg_16_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_17_config_addr;
assign config_reg_17_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
ConfigRegister_1_8_32_17 config_reg_17 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_17_O),
    .config_addr(config_reg_17_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_2_config_addr;
assign config_reg_2_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
ConfigRegister_32_8_32_2 config_reg_2 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_2_O),
    .config_addr(config_reg_2_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_3_config_addr;
assign config_reg_3_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
ConfigRegister_32_8_32_3 config_reg_3 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_3_O),
    .config_addr(config_reg_3_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_4_config_addr;
assign config_reg_4_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
ConfigRegister_32_8_32_4 config_reg_4 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_4_O),
    .config_addr(config_reg_4_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_5_config_addr;
assign config_reg_5_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
ConfigRegister_32_8_32_5 config_reg_5 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_5_O),
    .config_addr(config_reg_5_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_6_config_addr;
assign config_reg_6_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
ConfigRegister_32_8_32_6 config_reg_6 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_6_O),
    .config_addr(config_reg_6_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_7_config_addr;
assign config_reg_7_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
ConfigRegister_32_8_32_7 config_reg_7 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_7_O),
    .config_addr(config_reg_7_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_8_config_addr;
assign config_reg_8_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
ConfigRegister_30_8_32_8 config_reg_8 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_8_O),
    .config_addr(config_reg_8_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_9_config_addr;
assign config_reg_9_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5],self_config_config_addr_out[4:0]};
ConfigRegister_32_8_32_9 config_reg_9 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_9_O),
    .config_addr(config_reg_9_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_wrap coreir_wrapInAsyncReset_inst0 (
    .in(reset),
    .out(coreir_wrapInAsyncReset_inst0_out)
);
coreir_wrap coreir_wrapOutAsyncReset_inst0 (
    .in(Invert1_inst0_out[0]),
    .out(coreir_wrapOutAsyncReset_inst0_out)
);
wire [31:0] mux_aoi_18_32_inst0_I [17:0];
assign mux_aoi_18_32_inst0_I[17] = {ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,config_reg_17_O[0]};
assign mux_aoi_18_32_inst0_I[16] = config_reg_16_O;
assign mux_aoi_18_32_inst0_I[15] = config_reg_15_O;
assign mux_aoi_18_32_inst0_I[14] = config_reg_14_O;
assign mux_aoi_18_32_inst0_I[13] = config_reg_13_O;
assign mux_aoi_18_32_inst0_I[12] = config_reg_12_O;
assign mux_aoi_18_32_inst0_I[11] = config_reg_11_O;
assign mux_aoi_18_32_inst0_I[10] = config_reg_10_O;
assign mux_aoi_18_32_inst0_I[9] = config_reg_9_O;
assign mux_aoi_18_32_inst0_I[8] = ZextWrapper_30_32_inst0$self_O_in;
assign mux_aoi_18_32_inst0_I[7] = config_reg_7_O;
assign mux_aoi_18_32_inst0_I[6] = config_reg_6_O;
assign mux_aoi_18_32_inst0_I[5] = config_reg_5_O;
assign mux_aoi_18_32_inst0_I[4] = config_reg_4_O;
assign mux_aoi_18_32_inst0_I[3] = config_reg_3_O;
assign mux_aoi_18_32_inst0_I[2] = config_reg_2_O;
assign mux_aoi_18_32_inst0_I[1] = config_reg_1_O;
assign mux_aoi_18_32_inst0_I[0] = config_reg_0_O;
mux_aoi_18_32 mux_aoi_18_32_inst0 (
    .I(mux_aoi_18_32_inst0_I),
    .O(mux_aoi_18_32_inst0_O),
    .S(self_config_config_addr_out[4:0]),
    .out_sel(mux_aoi_18_32_inst0_out_sel)
);
coreir_or #(
    .width(1)
) or1_inst0 (
    .in0(flush_core),
    .in1(flush),
    .out(or1_inst0_out)
);
mantle_wire__typeBit8 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
SliceWrapper_1_0_1 tile_en_value (
    .I(config_reg_17_O),
    .O(tile_en_value_O)
);
assign PondTop_input_width_17_num_0_ready = bit_const_1_None_out;
assign PondTop_input_width_17_num_1_ready = bit_const_1_None_out;
assign PondTop_output_width_17_num_0 = PondTop_W_inst0_PondTop_output_width_17_num_0;
assign PondTop_output_width_17_num_0_valid = bit_const_1_None_out;
assign PondTop_output_width_17_num_1 = PondTop_W_inst0_PondTop_output_width_17_num_1;
assign PondTop_output_width_17_num_1_valid = bit_const_1_None_out;
assign PondTop_output_width_1_num_0 = PondTop_W_inst0_PondTop_output_width_1_num_0;
assign PondTop_output_width_1_num_0_valid = bit_const_1_None_out;
assign PondTop_output_width_1_num_1 = PondTop_W_inst0_PondTop_output_width_1_num_1;
assign PondTop_output_width_1_num_1_valid = bit_const_1_None_out;
assign read_config_data = mux_aoi_18_32_inst0_O;
assign read_config_data_1 = PondTop_W_inst0_config_data_out;
endmodule

module ConfigRegister_1_8_32_0 (
    input clk,
    input reset,
    output [0:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [0:0] Register_inst0_O;
wire [7:0] const_0_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq4 Register_inst0 (
    .I(config_data[0:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_0_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module PowerDomainConfigReg (
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [0:0] ps_en_out,
    output [31:0] read_config_data,
    input reset
);
wire ZextWrapper_1_32_inst0$bit_const_0_None_out;
wire [0:0] config_reg_0_O;
wire [0:0] ps_en_value_O;
corebit_const #(
    .value(1'b0)
) ZextWrapper_1_32_inst0$bit_const_0_None (
    .out(ZextWrapper_1_32_inst0$bit_const_0_None_out)
);
ConfigRegister_1_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
SliceWrapper_1_0_1 ps_en_value (
    .I(config_reg_0_O),
    .O(ps_en_value_O)
);
assign ps_en_out = ps_en_value_O;
assign read_config_data = {ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,ZextWrapper_1_32_inst0$bit_const_0_None_out,config_reg_0_O[0]};
endmodule

module ConfigRegister_19_8_32_40 (
    input clk,
    input reset,
    output [18:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [18:0] Register_inst0_O;
wire [7:0] const_40_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_unq7 Register_inst0 (
    .I(config_data[18:0]),
    .O(Register_inst0_O),
    .CE(magma_Bit_and_inst0_out),
    .CLK(clk),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h28),
    .width(8)
) const_40_8 (
    .out(const_40_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_40_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_inst0_O;
endmodule

module MemCore (
    input [16:0] MEM_input_width_17_num_0,
    output [0:0] MEM_input_width_17_num_0_ready,
    input [0:0] MEM_input_width_17_num_0_valid,
    input [16:0] MEM_input_width_17_num_1,
    output [0:0] MEM_input_width_17_num_1_ready,
    input [0:0] MEM_input_width_17_num_1_valid,
    input [16:0] MEM_input_width_17_num_2,
    output [0:0] MEM_input_width_17_num_2_ready,
    input [0:0] MEM_input_width_17_num_2_valid,
    input [16:0] MEM_input_width_17_num_3,
    output [0:0] MEM_input_width_17_num_3_ready,
    input [0:0] MEM_input_width_17_num_3_valid,
    input [0:0] MEM_input_width_1_num_0,
    output MEM_input_width_1_num_0_ready,
    input MEM_input_width_1_num_0_valid,
    input [0:0] MEM_input_width_1_num_1,
    output MEM_input_width_1_num_1_ready,
    input MEM_input_width_1_num_1_valid,
    output [16:0] MEM_output_width_17_num_0,
    input [0:0] MEM_output_width_17_num_0_ready,
    output [0:0] MEM_output_width_17_num_0_valid,
    output [16:0] MEM_output_width_17_num_1,
    input [0:0] MEM_output_width_17_num_1_ready,
    output [0:0] MEM_output_width_17_num_1_valid,
    output [16:0] MEM_output_width_17_num_2,
    input [0:0] MEM_output_width_17_num_2_ready,
    output [0:0] MEM_output_width_17_num_2_valid,
    output [0:0] MEM_output_width_1_num_0,
    input MEM_output_width_1_num_0_ready,
    output MEM_output_width_1_num_0_valid,
    output [0:0] MEM_output_width_1_num_1,
    input MEM_output_width_1_num_1_ready,
    output MEM_output_width_1_num_1_valid,
    output [0:0] MEM_output_width_1_num_2,
    input MEM_output_width_1_num_2_ready,
    output MEM_output_width_1_num_2_valid,
    input clk,
    input [7:0] config_1_config_addr,
    input [31:0] config_1_config_data,
    input [0:0] config_1_read,
    input [0:0] config_1_write,
    input [7:0] config_2_config_addr,
    input [31:0] config_2_config_data,
    input [0:0] config_2_read,
    input [0:0] config_2_write,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input config_en_0,
    input config_en_1,
    input [0:0] config_read,
    input [0:0] config_write,
    input [0:0] flush,
    input [0:0] flush_core,
    output [31:0] read_config_data,
    output [31:0] read_config_data_1,
    output [31:0] read_config_data_2,
    input reset,
    input [0:0] stall
);
wire [0:0] AND_CONFIG_EN_SRAM_0_out;
wire [0:0] AND_CONFIG_EN_SRAM_1_out;
wire [31:0] CONFIG_SPACE_0_value_O;
wire [31:0] CONFIG_SPACE_10_value_O;
wire [31:0] CONFIG_SPACE_11_value_O;
wire [31:0] CONFIG_SPACE_12_value_O;
wire [31:0] CONFIG_SPACE_13_value_O;
wire [31:0] CONFIG_SPACE_14_value_O;
wire [31:0] CONFIG_SPACE_15_value_O;
wire [31:0] CONFIG_SPACE_16_value_O;
wire [31:0] CONFIG_SPACE_17_value_O;
wire [31:0] CONFIG_SPACE_18_value_O;
wire [31:0] CONFIG_SPACE_19_value_O;
wire [31:0] CONFIG_SPACE_1_value_O;
wire [31:0] CONFIG_SPACE_20_value_O;
wire [31:0] CONFIG_SPACE_21_value_O;
wire [31:0] CONFIG_SPACE_22_value_O;
wire [31:0] CONFIG_SPACE_23_value_O;
wire [31:0] CONFIG_SPACE_24_value_O;
wire [31:0] CONFIG_SPACE_25_value_O;
wire [31:0] CONFIG_SPACE_26_value_O;
wire [31:0] CONFIG_SPACE_27_value_O;
wire [31:0] CONFIG_SPACE_28_value_O;
wire [31:0] CONFIG_SPACE_29_value_O;
wire [31:0] CONFIG_SPACE_2_value_O;
wire [31:0] CONFIG_SPACE_30_value_O;
wire [31:0] CONFIG_SPACE_31_value_O;
wire [31:0] CONFIG_SPACE_32_value_O;
wire [31:0] CONFIG_SPACE_33_value_O;
wire [31:0] CONFIG_SPACE_34_value_O;
wire [31:0] CONFIG_SPACE_35_value_O;
wire [31:0] CONFIG_SPACE_36_value_O;
wire [31:0] CONFIG_SPACE_37_value_O;
wire [31:0] CONFIG_SPACE_38_value_O;
wire [31:0] CONFIG_SPACE_39_value_O;
wire [31:0] CONFIG_SPACE_3_value_O;
wire [31:0] CONFIG_SPACE_40_value_O;
wire [31:0] CONFIG_SPACE_41_value_O;
wire [31:0] CONFIG_SPACE_42_value_O;
wire [31:0] CONFIG_SPACE_43_value_O;
wire [31:0] CONFIG_SPACE_44_value_O;
wire [18:0] CONFIG_SPACE_45_value_O;
wire [31:0] CONFIG_SPACE_4_value_O;
wire [31:0] CONFIG_SPACE_5_value_O;
wire [31:0] CONFIG_SPACE_6_value_O;
wire [31:0] CONFIG_SPACE_7_value_O;
wire [31:0] CONFIG_SPACE_8_value_O;
wire [31:0] CONFIG_SPACE_9_value_O;
wire [0:0] Invert1_inst0_out;
wire [0:0] Invert1_inst1_out;
wire [0:0] MEM_input_width_17_num_0_valid_reg_sel_value_O;
wire [0:0] MEM_input_width_17_num_0_valid_reg_value_value_O;
wire [0:0] MEM_input_width_17_num_0_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] MEM_input_width_17_num_1_valid_reg_sel_value_O;
wire [0:0] MEM_input_width_17_num_1_valid_reg_value_value_O;
wire [0:0] MEM_input_width_17_num_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] MEM_input_width_17_num_2_valid_reg_sel_value_O;
wire [0:0] MEM_input_width_17_num_2_valid_reg_value_value_O;
wire [0:0] MEM_input_width_17_num_2_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] MEM_input_width_17_num_3_valid_reg_sel_value_O;
wire [0:0] MEM_input_width_17_num_3_valid_reg_value_value_O;
wire [0:0] MEM_input_width_17_num_3_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] MEM_input_width_1_num_0_reg_sel_value_O;
wire [0:0] MEM_input_width_1_num_0_reg_value_value_O;
wire [0:0] MEM_input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] MEM_input_width_1_num_1_reg_sel_value_O;
wire [0:0] MEM_input_width_1_num_1_reg_value_value_O;
wire [0:0] MEM_input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] MEM_output_width_17_num_0_ready_reg_sel_value_O;
wire [0:0] MEM_output_width_17_num_0_ready_reg_value_value_O;
wire [0:0] MEM_output_width_17_num_0_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] MEM_output_width_17_num_1_ready_reg_sel_value_O;
wire [0:0] MEM_output_width_17_num_1_ready_reg_value_value_O;
wire [0:0] MEM_output_width_17_num_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] MEM_output_width_17_num_2_ready_reg_sel_value_O;
wire [0:0] MEM_output_width_17_num_2_ready_reg_value_value_O;
wire [0:0] MEM_output_width_17_num_2_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [31:0] MemCore_inner_W_inst0_config_data_out_1;
wire [0:0] MemCore_inner_W_inst0_MEM_output_width_1_num_1;
wire [0:0] MemCore_inner_W_inst0_MEM_output_width_17_num_1_valid;
wire [16:0] MemCore_inner_W_inst0_MEM_output_width_17_num_2;
wire [0:0] MemCore_inner_W_inst0_MEM_input_width_17_num_2_ready;
wire [0:0] MemCore_inner_W_inst0_MEM_output_width_17_num_0_valid;
wire [0:0] MemCore_inner_W_inst0_MEM_input_width_17_num_1_ready;
wire [0:0] MemCore_inner_W_inst0_MEM_input_width_17_num_0_ready;
wire [0:0] MemCore_inner_W_inst0_MEM_output_width_1_num_0;
wire [0:0] MemCore_inner_W_inst0_MEM_output_width_17_num_2_valid;
wire [16:0] MemCore_inner_W_inst0_MEM_output_width_17_num_1;
wire [16:0] MemCore_inner_W_inst0_MEM_output_width_17_num_0;
wire [0:0] MemCore_inner_W_inst0_MEM_output_width_1_num_2;
wire [31:0] MemCore_inner_W_inst0_config_data_out_0;
wire [0:0] MemCore_inner_W_inst0_MEM_input_width_17_num_3_ready;
wire [0:0] OR_CONFIG_EN_SRAM_0_out;
wire [0:0] OR_CONFIG_EN_SRAM_1_out;
wire [0:0] OR_CONFIG_RD_SRAM_out;
wire [0:0] OR_CONFIG_WR_SRAM_out;
wire [7:0] OR_config_addr_FEATURE_O;
wire [31:0] OR_config_data_FEATURE_O;
wire ZextWrapper_19_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_19_32_inst0$self_O_in;
wire ZextWrapper_25_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_25_32_inst0$self_O_in;
wire bit_const_1_None_out;
wire [31:0] config_reg_0_O;
wire [31:0] config_reg_1_O;
wire [31:0] config_reg_10_O;
wire [31:0] config_reg_11_O;
wire [31:0] config_reg_12_O;
wire [31:0] config_reg_13_O;
wire [31:0] config_reg_14_O;
wire [31:0] config_reg_15_O;
wire [31:0] config_reg_16_O;
wire [31:0] config_reg_17_O;
wire [31:0] config_reg_18_O;
wire [31:0] config_reg_19_O;
wire [31:0] config_reg_2_O;
wire [31:0] config_reg_20_O;
wire [31:0] config_reg_21_O;
wire [31:0] config_reg_22_O;
wire [31:0] config_reg_23_O;
wire [31:0] config_reg_24_O;
wire [31:0] config_reg_25_O;
wire [31:0] config_reg_26_O;
wire [31:0] config_reg_27_O;
wire [31:0] config_reg_28_O;
wire [31:0] config_reg_29_O;
wire [31:0] config_reg_3_O;
wire [31:0] config_reg_30_O;
wire [31:0] config_reg_31_O;
wire [31:0] config_reg_32_O;
wire [31:0] config_reg_33_O;
wire [31:0] config_reg_34_O;
wire [31:0] config_reg_35_O;
wire [31:0] config_reg_36_O;
wire [31:0] config_reg_37_O;
wire [31:0] config_reg_38_O;
wire [31:0] config_reg_39_O;
wire [31:0] config_reg_4_O;
wire [18:0] config_reg_40_O;
wire [31:0] config_reg_41_O;
wire [31:0] config_reg_42_O;
wire [31:0] config_reg_43_O;
wire [31:0] config_reg_44_O;
wire [31:0] config_reg_45_O;
wire [24:0] config_reg_46_O;
wire [31:0] config_reg_5_O;
wire [31:0] config_reg_6_O;
wire [31:0] config_reg_7_O;
wire [31:0] config_reg_8_O;
wire [31:0] config_reg_9_O;
wire coreir_wrapInAsyncReset_inst0_out;
wire coreir_wrapOutAsyncReset_inst0_out;
wire [0:0] flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] flush_mux_sel_value_O;
wire [0:0] flush_reg_sel_value_O;
wire [0:0] flush_reg_value_value_O;
wire [0:0] flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] mode_excl_value_O;
wire [1:0] mode_value_O;
wire [31:0] mux_aoi_47_32_inst0_O;
wire [63:0] mux_aoi_47_32_inst0_out_sel;
wire [7:0] self_config_config_addr_out;
wire [0:0] tile_en_value_O;
coreir_and #(
    .width(1)
) AND_CONFIG_EN_SRAM_0 (
    .in0(OR_CONFIG_EN_SRAM_0_out),
    .in1(config_en_0),
    .out(AND_CONFIG_EN_SRAM_0_out)
);
coreir_and #(
    .width(1)
) AND_CONFIG_EN_SRAM_1 (
    .in0(OR_CONFIG_EN_SRAM_1_out),
    .in1(config_en_1),
    .out(AND_CONFIG_EN_SRAM_1_out)
);
SliceWrapper_32_0_32 CONFIG_SPACE_0_value (
    .I(config_reg_0_O),
    .O(CONFIG_SPACE_0_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_10_value (
    .I(config_reg_2_O),
    .O(CONFIG_SPACE_10_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_11_value (
    .I(config_reg_3_O),
    .O(CONFIG_SPACE_11_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_12_value (
    .I(config_reg_4_O),
    .O(CONFIG_SPACE_12_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_13_value (
    .I(config_reg_5_O),
    .O(CONFIG_SPACE_13_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_14_value (
    .I(config_reg_6_O),
    .O(CONFIG_SPACE_14_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_15_value (
    .I(config_reg_7_O),
    .O(CONFIG_SPACE_15_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_16_value (
    .I(config_reg_8_O),
    .O(CONFIG_SPACE_16_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_17_value (
    .I(config_reg_9_O),
    .O(CONFIG_SPACE_17_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_18_value (
    .I(config_reg_10_O),
    .O(CONFIG_SPACE_18_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_19_value (
    .I(config_reg_11_O),
    .O(CONFIG_SPACE_19_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_1_value (
    .I(config_reg_1_O),
    .O(CONFIG_SPACE_1_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_20_value (
    .I(config_reg_13_O),
    .O(CONFIG_SPACE_20_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_21_value (
    .I(config_reg_14_O),
    .O(CONFIG_SPACE_21_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_22_value (
    .I(config_reg_15_O),
    .O(CONFIG_SPACE_22_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_23_value (
    .I(config_reg_16_O),
    .O(CONFIG_SPACE_23_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_24_value (
    .I(config_reg_17_O),
    .O(CONFIG_SPACE_24_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_25_value (
    .I(config_reg_18_O),
    .O(CONFIG_SPACE_25_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_26_value (
    .I(config_reg_19_O),
    .O(CONFIG_SPACE_26_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_27_value (
    .I(config_reg_20_O),
    .O(CONFIG_SPACE_27_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_28_value (
    .I(config_reg_21_O),
    .O(CONFIG_SPACE_28_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_29_value (
    .I(config_reg_22_O),
    .O(CONFIG_SPACE_29_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_2_value (
    .I(config_reg_12_O),
    .O(CONFIG_SPACE_2_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_30_value (
    .I(config_reg_24_O),
    .O(CONFIG_SPACE_30_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_31_value (
    .I(config_reg_25_O),
    .O(CONFIG_SPACE_31_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_32_value (
    .I(config_reg_26_O),
    .O(CONFIG_SPACE_32_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_33_value (
    .I(config_reg_27_O),
    .O(CONFIG_SPACE_33_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_34_value (
    .I(config_reg_28_O),
    .O(CONFIG_SPACE_34_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_35_value (
    .I(config_reg_29_O),
    .O(CONFIG_SPACE_35_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_36_value (
    .I(config_reg_30_O),
    .O(CONFIG_SPACE_36_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_37_value (
    .I(config_reg_31_O),
    .O(CONFIG_SPACE_37_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_38_value (
    .I(config_reg_32_O),
    .O(CONFIG_SPACE_38_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_39_value (
    .I(config_reg_33_O),
    .O(CONFIG_SPACE_39_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_3_value (
    .I(config_reg_23_O),
    .O(CONFIG_SPACE_3_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_40_value (
    .I(config_reg_35_O),
    .O(CONFIG_SPACE_40_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_41_value (
    .I(config_reg_36_O),
    .O(CONFIG_SPACE_41_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_42_value (
    .I(config_reg_37_O),
    .O(CONFIG_SPACE_42_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_43_value (
    .I(config_reg_38_O),
    .O(CONFIG_SPACE_43_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_44_value (
    .I(config_reg_39_O),
    .O(CONFIG_SPACE_44_value_O)
);
SliceWrapper_19_0_19 CONFIG_SPACE_45_value (
    .I(config_reg_40_O),
    .O(CONFIG_SPACE_45_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_4_value (
    .I(config_reg_34_O),
    .O(CONFIG_SPACE_4_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_5_value (
    .I(config_reg_41_O),
    .O(CONFIG_SPACE_5_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_6_value (
    .I(config_reg_42_O),
    .O(CONFIG_SPACE_6_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_7_value (
    .I(config_reg_43_O),
    .O(CONFIG_SPACE_7_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_8_value (
    .I(config_reg_44_O),
    .O(CONFIG_SPACE_8_value_O)
);
SliceWrapper_32_0_32 CONFIG_SPACE_9_value (
    .I(config_reg_45_O),
    .O(CONFIG_SPACE_9_value_O)
);
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(coreir_wrapInAsyncReset_inst0_out),
    .out(Invert1_inst0_out)
);
coreir_not #(
    .width(1)
) Invert1_inst1 (
    .in(stall),
    .out(Invert1_inst1_out)
);
SliceWrapper_25_0_1 MEM_input_width_17_num_0_valid_reg_sel_value (
    .I(config_reg_46_O),
    .O(MEM_input_width_17_num_0_valid_reg_sel_value_O)
);
SliceWrapper_25_1_2 MEM_input_width_17_num_0_valid_reg_value_value (
    .I(config_reg_46_O),
    .O(MEM_input_width_17_num_0_valid_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) MEM_input_width_17_num_0_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MEM_input_width_17_num_0_valid),
    .in1(MEM_input_width_17_num_0_valid_reg_value_value_O),
    .sel(MEM_input_width_17_num_0_valid_reg_sel_value_O[0]),
    .out(MEM_input_width_17_num_0_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_25_2_3 MEM_input_width_17_num_1_valid_reg_sel_value (
    .I(config_reg_46_O),
    .O(MEM_input_width_17_num_1_valid_reg_sel_value_O)
);
SliceWrapper_25_3_4 MEM_input_width_17_num_1_valid_reg_value_value (
    .I(config_reg_46_O),
    .O(MEM_input_width_17_num_1_valid_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) MEM_input_width_17_num_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MEM_input_width_17_num_1_valid),
    .in1(MEM_input_width_17_num_1_valid_reg_value_value_O),
    .sel(MEM_input_width_17_num_1_valid_reg_sel_value_O[0]),
    .out(MEM_input_width_17_num_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_25_4_5 MEM_input_width_17_num_2_valid_reg_sel_value (
    .I(config_reg_46_O),
    .O(MEM_input_width_17_num_2_valid_reg_sel_value_O)
);
SliceWrapper_25_5_6 MEM_input_width_17_num_2_valid_reg_value_value (
    .I(config_reg_46_O),
    .O(MEM_input_width_17_num_2_valid_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) MEM_input_width_17_num_2_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MEM_input_width_17_num_2_valid),
    .in1(MEM_input_width_17_num_2_valid_reg_value_value_O),
    .sel(MEM_input_width_17_num_2_valid_reg_sel_value_O[0]),
    .out(MEM_input_width_17_num_2_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_25_6_7 MEM_input_width_17_num_3_valid_reg_sel_value (
    .I(config_reg_46_O),
    .O(MEM_input_width_17_num_3_valid_reg_sel_value_O)
);
SliceWrapper_25_7_8 MEM_input_width_17_num_3_valid_reg_value_value (
    .I(config_reg_46_O),
    .O(MEM_input_width_17_num_3_valid_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) MEM_input_width_17_num_3_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MEM_input_width_17_num_3_valid),
    .in1(MEM_input_width_17_num_3_valid_reg_value_value_O),
    .sel(MEM_input_width_17_num_3_valid_reg_sel_value_O[0]),
    .out(MEM_input_width_17_num_3_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_25_8_9 MEM_input_width_1_num_0_reg_sel_value (
    .I(config_reg_46_O),
    .O(MEM_input_width_1_num_0_reg_sel_value_O)
);
SliceWrapper_25_9_10 MEM_input_width_1_num_0_reg_value_value (
    .I(config_reg_46_O),
    .O(MEM_input_width_1_num_0_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) MEM_input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MEM_input_width_1_num_0),
    .in1(MEM_input_width_1_num_0_reg_value_value_O),
    .sel(MEM_input_width_1_num_0_reg_sel_value_O[0]),
    .out(MEM_input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_25_10_11 MEM_input_width_1_num_1_reg_sel_value (
    .I(config_reg_46_O),
    .O(MEM_input_width_1_num_1_reg_sel_value_O)
);
SliceWrapper_25_11_12 MEM_input_width_1_num_1_reg_value_value (
    .I(config_reg_46_O),
    .O(MEM_input_width_1_num_1_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) MEM_input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MEM_input_width_1_num_1),
    .in1(MEM_input_width_1_num_1_reg_value_value_O),
    .sel(MEM_input_width_1_num_1_reg_sel_value_O[0]),
    .out(MEM_input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_25_12_13 MEM_output_width_17_num_0_ready_reg_sel_value (
    .I(config_reg_46_O),
    .O(MEM_output_width_17_num_0_ready_reg_sel_value_O)
);
SliceWrapper_25_13_14 MEM_output_width_17_num_0_ready_reg_value_value (
    .I(config_reg_46_O),
    .O(MEM_output_width_17_num_0_ready_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) MEM_output_width_17_num_0_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MEM_output_width_17_num_0_ready),
    .in1(MEM_output_width_17_num_0_ready_reg_value_value_O),
    .sel(MEM_output_width_17_num_0_ready_reg_sel_value_O[0]),
    .out(MEM_output_width_17_num_0_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_25_14_15 MEM_output_width_17_num_1_ready_reg_sel_value (
    .I(config_reg_46_O),
    .O(MEM_output_width_17_num_1_ready_reg_sel_value_O)
);
SliceWrapper_25_15_16 MEM_output_width_17_num_1_ready_reg_value_value (
    .I(config_reg_46_O),
    .O(MEM_output_width_17_num_1_ready_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) MEM_output_width_17_num_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MEM_output_width_17_num_1_ready),
    .in1(MEM_output_width_17_num_1_ready_reg_value_value_O),
    .sel(MEM_output_width_17_num_1_ready_reg_sel_value_O[0]),
    .out(MEM_output_width_17_num_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_25_16_17 MEM_output_width_17_num_2_ready_reg_sel_value (
    .I(config_reg_46_O),
    .O(MEM_output_width_17_num_2_ready_reg_sel_value_O)
);
SliceWrapper_25_17_18 MEM_output_width_17_num_2_ready_reg_value_value (
    .I(config_reg_46_O),
    .O(MEM_output_width_17_num_2_ready_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) MEM_output_width_17_num_2_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MEM_output_width_17_num_2_ready),
    .in1(MEM_output_width_17_num_2_ready_reg_value_value_O),
    .sel(MEM_output_width_17_num_2_ready_reg_sel_value_O[0]),
    .out(MEM_output_width_17_num_2_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
wire [1:0] MemCore_inner_W_inst0_config_en;
assign MemCore_inner_W_inst0_config_en = {AND_CONFIG_EN_SRAM_1_out[0],AND_CONFIG_EN_SRAM_0_out[0]};
MemCore_inner_W MemCore_inner_W_inst0 (
    .CONFIG_SPACE_5(CONFIG_SPACE_5_value_O),
    .mode(mode_value_O),
    .CONFIG_SPACE_35(CONFIG_SPACE_35_value_O),
    .config_data_out_1(MemCore_inner_W_inst0_config_data_out_1),
    .MEM_input_width_1_num_0(MEM_input_width_1_num_0_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .CONFIG_SPACE_41(CONFIG_SPACE_41_value_O),
    .CONFIG_SPACE_3(CONFIG_SPACE_3_value_O),
    .CONFIG_SPACE_26(CONFIG_SPACE_26_value_O),
    .tile_en(tile_en_value_O),
    .config_read(OR_CONFIG_WR_SRAM_out),
    .clk(clk),
    .CONFIG_SPACE_28(CONFIG_SPACE_28_value_O),
    .CONFIG_SPACE_18(CONFIG_SPACE_18_value_O),
    .MEM_input_width_17_num_2(MEM_input_width_17_num_2),
    .config_write(OR_CONFIG_RD_SRAM_out),
    .MEM_output_width_1_num_1(MemCore_inner_W_inst0_MEM_output_width_1_num_1),
    .CONFIG_SPACE_29(CONFIG_SPACE_29_value_O),
    .clk_en(Invert1_inst1_out),
    .CONFIG_SPACE_17(CONFIG_SPACE_17_value_O),
    .CONFIG_SPACE_2(CONFIG_SPACE_2_value_O),
    .CONFIG_SPACE_23(CONFIG_SPACE_23_value_O),
    .CONFIG_SPACE_21(CONFIG_SPACE_21_value_O),
    .MEM_output_width_17_num_1_valid(MemCore_inner_W_inst0_MEM_output_width_17_num_1_valid),
    .CONFIG_SPACE_10(CONFIG_SPACE_10_value_O),
    .rst_n(coreir_wrapOutAsyncReset_inst0_out),
    .MEM_output_width_17_num_2(MemCore_inner_W_inst0_MEM_output_width_17_num_2),
    .CONFIG_SPACE_15(CONFIG_SPACE_15_value_O),
    .MEM_input_width_17_num_3(MEM_input_width_17_num_3),
    .CONFIG_SPACE_31(CONFIG_SPACE_31_value_O),
    .CONFIG_SPACE_13(CONFIG_SPACE_13_value_O),
    .CONFIG_SPACE_36(CONFIG_SPACE_36_value_O),
    .CONFIG_SPACE_42(CONFIG_SPACE_42_value_O),
    .MEM_input_width_17_num_2_ready(MemCore_inner_W_inst0_MEM_input_width_17_num_2_ready),
    .CONFIG_SPACE_24(CONFIG_SPACE_24_value_O),
    .CONFIG_SPACE_12(CONFIG_SPACE_12_value_O),
    .CONFIG_SPACE_37(CONFIG_SPACE_37_value_O),
    .CONFIG_SPACE_30(CONFIG_SPACE_30_value_O),
    .CONFIG_SPACE_27(CONFIG_SPACE_27_value_O),
    .CONFIG_SPACE_45(CONFIG_SPACE_45_value_O),
    .CONFIG_SPACE_25(CONFIG_SPACE_25_value_O),
    .CONFIG_SPACE_38(CONFIG_SPACE_38_value_O),
    .MEM_output_width_17_num_0_valid(MemCore_inner_W_inst0_MEM_output_width_17_num_0_valid),
    .config_data_in(OR_config_data_FEATURE_O),
    .MEM_output_width_17_num_0_ready(MEM_output_width_17_num_0_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .config_en(MemCore_inner_W_inst0_config_en),
    .CONFIG_SPACE_11(CONFIG_SPACE_11_value_O),
    .CONFIG_SPACE_6(CONFIG_SPACE_6_value_O),
    .MEM_input_width_17_num_1_ready(MemCore_inner_W_inst0_MEM_input_width_17_num_1_ready),
    .MEM_input_width_17_num_2_valid(MEM_input_width_17_num_2_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .MEM_input_width_17_num_0_valid(MEM_input_width_17_num_0_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .MEM_input_width_17_num_0_ready(MemCore_inner_W_inst0_MEM_input_width_17_num_0_ready),
    .MEM_output_width_1_num_0(MemCore_inner_W_inst0_MEM_output_width_1_num_0),
    .MEM_output_width_17_num_2_valid(MemCore_inner_W_inst0_MEM_output_width_17_num_2_valid),
    .CONFIG_SPACE_9(CONFIG_SPACE_9_value_O),
    .CONFIG_SPACE_34(CONFIG_SPACE_34_value_O),
    .CONFIG_SPACE_44(CONFIG_SPACE_44_value_O),
    .MEM_output_width_17_num_2_ready(MEM_output_width_17_num_2_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .MEM_output_width_17_num_1(MemCore_inner_W_inst0_MEM_output_width_17_num_1),
    .CONFIG_SPACE_32(CONFIG_SPACE_32_value_O),
    .MEM_input_width_17_num_0(MEM_input_width_17_num_0),
    .MEM_input_width_17_num_1(MEM_input_width_17_num_1),
    .CONFIG_SPACE_39(CONFIG_SPACE_39_value_O),
    .CONFIG_SPACE_22(CONFIG_SPACE_22_value_O),
    .CONFIG_SPACE_0(CONFIG_SPACE_0_value_O),
    .CONFIG_SPACE_8(CONFIG_SPACE_8_value_O),
    .MEM_output_width_17_num_0(MemCore_inner_W_inst0_MEM_output_width_17_num_0),
    .CONFIG_SPACE_40(CONFIG_SPACE_40_value_O),
    .CONFIG_SPACE_14(CONFIG_SPACE_14_value_O),
    .config_addr_in(OR_config_addr_FEATURE_O),
    .MEM_input_width_1_num_1(MEM_input_width_1_num_1_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .CONFIG_SPACE_1(CONFIG_SPACE_1_value_O),
    .MEM_output_width_1_num_2(MemCore_inner_W_inst0_MEM_output_width_1_num_2),
    .CONFIG_SPACE_7(CONFIG_SPACE_7_value_O),
    .CONFIG_SPACE_4(CONFIG_SPACE_4_value_O),
    .CONFIG_SPACE_20(CONFIG_SPACE_20_value_O),
    .config_data_out_0(MemCore_inner_W_inst0_config_data_out_0),
    .CONFIG_SPACE_33(CONFIG_SPACE_33_value_O),
    .CONFIG_SPACE_16(CONFIG_SPACE_16_value_O),
    .CONFIG_SPACE_43(CONFIG_SPACE_43_value_O),
    .MEM_input_width_17_num_3_ready(MemCore_inner_W_inst0_MEM_input_width_17_num_3_ready),
    .MEM_output_width_17_num_1_ready(MEM_output_width_17_num_1_ready_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .CONFIG_SPACE_19(CONFIG_SPACE_19_value_O),
    .MEM_input_width_17_num_1_valid(MEM_input_width_17_num_1_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .mode_excl(mode_excl_value_O),
    .flush(flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .MEM_input_width_17_num_3_valid(MEM_input_width_17_num_3_valid_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_or #(
    .width(1)
) OR_CONFIG_EN_SRAM_0 (
    .in0(config_1_write),
    .in1(config_1_read),
    .out(OR_CONFIG_EN_SRAM_0_out)
);
coreir_or #(
    .width(1)
) OR_CONFIG_EN_SRAM_1 (
    .in0(config_2_write),
    .in1(config_2_read),
    .out(OR_CONFIG_EN_SRAM_1_out)
);
coreir_or #(
    .width(1)
) OR_CONFIG_RD_SRAM (
    .in0(config_1_write),
    .in1(config_2_write),
    .out(OR_CONFIG_RD_SRAM_out)
);
coreir_or #(
    .width(1)
) OR_CONFIG_WR_SRAM (
    .in0(config_1_read),
    .in1(config_2_read),
    .out(OR_CONFIG_WR_SRAM_out)
);
wire [7:0] OR_config_addr_FEATURE_I0;
assign OR_config_addr_FEATURE_I0 = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
Or3x8 OR_config_addr_FEATURE (
    .I0(OR_config_addr_FEATURE_I0),
    .I1(config_1_config_addr),
    .I2(config_2_config_addr),
    .O(OR_config_addr_FEATURE_O)
);
Or3x32 OR_config_data_FEATURE (
    .I0(config_config_data),
    .I1(config_1_config_data),
    .I2(config_2_config_data),
    .O(OR_config_data_FEATURE_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_19_32_inst0$bit_const_0_None (
    .out(ZextWrapper_19_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_19_32_inst0$self_O_out;
assign ZextWrapper_19_32_inst0$self_O_out = {ZextWrapper_19_32_inst0$bit_const_0_None_out,ZextWrapper_19_32_inst0$bit_const_0_None_out,ZextWrapper_19_32_inst0$bit_const_0_None_out,ZextWrapper_19_32_inst0$bit_const_0_None_out,ZextWrapper_19_32_inst0$bit_const_0_None_out,ZextWrapper_19_32_inst0$bit_const_0_None_out,ZextWrapper_19_32_inst0$bit_const_0_None_out,ZextWrapper_19_32_inst0$bit_const_0_None_out,ZextWrapper_19_32_inst0$bit_const_0_None_out,ZextWrapper_19_32_inst0$bit_const_0_None_out,ZextWrapper_19_32_inst0$bit_const_0_None_out,ZextWrapper_19_32_inst0$bit_const_0_None_out,ZextWrapper_19_32_inst0$bit_const_0_None_out,config_reg_40_O};
mantle_wire__typeBitIn32 ZextWrapper_19_32_inst0$self_O (
    .in(ZextWrapper_19_32_inst0$self_O_in),
    .out(ZextWrapper_19_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_25_32_inst0$bit_const_0_None (
    .out(ZextWrapper_25_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_25_32_inst0$self_O_out;
assign ZextWrapper_25_32_inst0$self_O_out = {ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$bit_const_0_None_out,config_reg_46_O};
mantle_wire__typeBitIn32 ZextWrapper_25_32_inst0$self_O (
    .in(ZextWrapper_25_32_inst0$self_O_in),
    .out(ZextWrapper_25_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b1)
) bit_const_1_None (
    .out(bit_const_1_None_out)
);
wire [7:0] config_reg_0_config_addr;
assign config_reg_0_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_reg_0_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_1_config_addr;
assign config_reg_1_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_reg_1_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_10_config_addr;
assign config_reg_10_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_10 config_reg_10 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_10_O),
    .config_addr(config_reg_10_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_11_config_addr;
assign config_reg_11_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_11 config_reg_11 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_11_O),
    .config_addr(config_reg_11_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_12_config_addr;
assign config_reg_12_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_12 config_reg_12 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_12_O),
    .config_addr(config_reg_12_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_13_config_addr;
assign config_reg_13_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_13 config_reg_13 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_13_O),
    .config_addr(config_reg_13_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_14_config_addr;
assign config_reg_14_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_14 config_reg_14 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_14_O),
    .config_addr(config_reg_14_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_15_config_addr;
assign config_reg_15_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_15 config_reg_15 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_15_O),
    .config_addr(config_reg_15_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_16_config_addr;
assign config_reg_16_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_16 config_reg_16 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_16_O),
    .config_addr(config_reg_16_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_17_config_addr;
assign config_reg_17_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_17 config_reg_17 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_17_O),
    .config_addr(config_reg_17_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_18_config_addr;
assign config_reg_18_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_18 config_reg_18 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_18_O),
    .config_addr(config_reg_18_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_19_config_addr;
assign config_reg_19_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_19 config_reg_19 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_19_O),
    .config_addr(config_reg_19_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_2_config_addr;
assign config_reg_2_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_2 config_reg_2 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_2_O),
    .config_addr(config_reg_2_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_20_config_addr;
assign config_reg_20_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_20 config_reg_20 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_20_O),
    .config_addr(config_reg_20_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_21_config_addr;
assign config_reg_21_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_21 config_reg_21 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_21_O),
    .config_addr(config_reg_21_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_22_config_addr;
assign config_reg_22_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_22 config_reg_22 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_22_O),
    .config_addr(config_reg_22_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_23_config_addr;
assign config_reg_23_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_23 config_reg_23 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_23_O),
    .config_addr(config_reg_23_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_24_config_addr;
assign config_reg_24_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_24 config_reg_24 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_24_O),
    .config_addr(config_reg_24_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_25_config_addr;
assign config_reg_25_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_25 config_reg_25 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_25_O),
    .config_addr(config_reg_25_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_26_config_addr;
assign config_reg_26_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_26 config_reg_26 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_26_O),
    .config_addr(config_reg_26_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_27_config_addr;
assign config_reg_27_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_27 config_reg_27 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_27_O),
    .config_addr(config_reg_27_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_28_config_addr;
assign config_reg_28_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_28 config_reg_28 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_28_O),
    .config_addr(config_reg_28_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_29_config_addr;
assign config_reg_29_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_29 config_reg_29 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_29_O),
    .config_addr(config_reg_29_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_3_config_addr;
assign config_reg_3_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_3 config_reg_3 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_3_O),
    .config_addr(config_reg_3_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_30_config_addr;
assign config_reg_30_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_30 config_reg_30 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_30_O),
    .config_addr(config_reg_30_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_31_config_addr;
assign config_reg_31_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_31 config_reg_31 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_31_O),
    .config_addr(config_reg_31_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_32_config_addr;
assign config_reg_32_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_32 config_reg_32 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_32_O),
    .config_addr(config_reg_32_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_33_config_addr;
assign config_reg_33_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_33 config_reg_33 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_33_O),
    .config_addr(config_reg_33_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_34_config_addr;
assign config_reg_34_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_34 config_reg_34 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_34_O),
    .config_addr(config_reg_34_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_35_config_addr;
assign config_reg_35_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_35 config_reg_35 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_35_O),
    .config_addr(config_reg_35_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_36_config_addr;
assign config_reg_36_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_36 config_reg_36 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_36_O),
    .config_addr(config_reg_36_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_37_config_addr;
assign config_reg_37_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_37 config_reg_37 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_37_O),
    .config_addr(config_reg_37_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_38_config_addr;
assign config_reg_38_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_38 config_reg_38 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_38_O),
    .config_addr(config_reg_38_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_39_config_addr;
assign config_reg_39_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_39 config_reg_39 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_39_O),
    .config_addr(config_reg_39_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_4_config_addr;
assign config_reg_4_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_4 config_reg_4 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_4_O),
    .config_addr(config_reg_4_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_40_config_addr;
assign config_reg_40_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_19_8_32_40 config_reg_40 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_40_O),
    .config_addr(config_reg_40_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_41_config_addr;
assign config_reg_41_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_41 config_reg_41 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_41_O),
    .config_addr(config_reg_41_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_42_config_addr;
assign config_reg_42_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_42 config_reg_42 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_42_O),
    .config_addr(config_reg_42_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_43_config_addr;
assign config_reg_43_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_43 config_reg_43 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_43_O),
    .config_addr(config_reg_43_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_44_config_addr;
assign config_reg_44_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_44 config_reg_44 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_44_O),
    .config_addr(config_reg_44_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_45_config_addr;
assign config_reg_45_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_45 config_reg_45 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_45_O),
    .config_addr(config_reg_45_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_46_config_addr;
assign config_reg_46_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_25_8_32_46 config_reg_46 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_46_O),
    .config_addr(config_reg_46_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_5_config_addr;
assign config_reg_5_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_5 config_reg_5 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_5_O),
    .config_addr(config_reg_5_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_6_config_addr;
assign config_reg_6_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_6 config_reg_6 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_6_O),
    .config_addr(config_reg_6_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_7_config_addr;
assign config_reg_7_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_7 config_reg_7 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_7_O),
    .config_addr(config_reg_7_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_8_config_addr;
assign config_reg_8_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_8 config_reg_8 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_8_O),
    .config_addr(config_reg_8_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
wire [7:0] config_reg_9_config_addr;
assign config_reg_9_config_addr = {self_config_config_addr_out[7],self_config_config_addr_out[6],self_config_config_addr_out[5:0]};
ConfigRegister_32_8_32_9 config_reg_9 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_9_O),
    .config_addr(config_reg_9_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_wrap coreir_wrapInAsyncReset_inst0 (
    .in(reset),
    .out(coreir_wrapInAsyncReset_inst0_out)
);
coreir_wrap coreir_wrapOutAsyncReset_inst0 (
    .in(Invert1_inst0_out[0]),
    .out(coreir_wrapOutAsyncReset_inst0_out)
);
coreir_mux #(
    .width(1)
) flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(flush_core),
    .in1(flush),
    .sel(flush_mux_sel_value_O[0]),
    .out(flush_mux$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_25_18_19 flush_mux_sel_value (
    .I(config_reg_46_O),
    .O(flush_mux_sel_value_O)
);
SliceWrapper_25_19_20 flush_reg_sel_value (
    .I(config_reg_46_O),
    .O(flush_reg_sel_value_O)
);
SliceWrapper_25_20_21 flush_reg_value_value (
    .I(config_reg_46_O),
    .O(flush_reg_value_value_O)
);
coreir_mux #(
    .width(1)
) flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(flush),
    .in1(flush_reg_value_value_O),
    .sel(flush_reg_sel_value_O[0]),
    .out(flush_sel$Mux2xBits1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
SliceWrapper_25_23_24 mode_excl_value (
    .I(config_reg_46_O),
    .O(mode_excl_value_O)
);
SliceWrapper_25_21_23 mode_value (
    .I(config_reg_46_O),
    .O(mode_value_O)
);
wire [31:0] mux_aoi_47_32_inst0_I [46:0];
assign mux_aoi_47_32_inst0_I[46] = ZextWrapper_25_32_inst0$self_O_in;
assign mux_aoi_47_32_inst0_I[45] = config_reg_45_O;
assign mux_aoi_47_32_inst0_I[44] = config_reg_44_O;
assign mux_aoi_47_32_inst0_I[43] = config_reg_43_O;
assign mux_aoi_47_32_inst0_I[42] = config_reg_42_O;
assign mux_aoi_47_32_inst0_I[41] = config_reg_41_O;
assign mux_aoi_47_32_inst0_I[40] = ZextWrapper_19_32_inst0$self_O_in;
assign mux_aoi_47_32_inst0_I[39] = config_reg_39_O;
assign mux_aoi_47_32_inst0_I[38] = config_reg_38_O;
assign mux_aoi_47_32_inst0_I[37] = config_reg_37_O;
assign mux_aoi_47_32_inst0_I[36] = config_reg_36_O;
assign mux_aoi_47_32_inst0_I[35] = config_reg_35_O;
assign mux_aoi_47_32_inst0_I[34] = config_reg_34_O;
assign mux_aoi_47_32_inst0_I[33] = config_reg_33_O;
assign mux_aoi_47_32_inst0_I[32] = config_reg_32_O;
assign mux_aoi_47_32_inst0_I[31] = config_reg_31_O;
assign mux_aoi_47_32_inst0_I[30] = config_reg_30_O;
assign mux_aoi_47_32_inst0_I[29] = config_reg_29_O;
assign mux_aoi_47_32_inst0_I[28] = config_reg_28_O;
assign mux_aoi_47_32_inst0_I[27] = config_reg_27_O;
assign mux_aoi_47_32_inst0_I[26] = config_reg_26_O;
assign mux_aoi_47_32_inst0_I[25] = config_reg_25_O;
assign mux_aoi_47_32_inst0_I[24] = config_reg_24_O;
assign mux_aoi_47_32_inst0_I[23] = config_reg_23_O;
assign mux_aoi_47_32_inst0_I[22] = config_reg_22_O;
assign mux_aoi_47_32_inst0_I[21] = config_reg_21_O;
assign mux_aoi_47_32_inst0_I[20] = config_reg_20_O;
assign mux_aoi_47_32_inst0_I[19] = config_reg_19_O;
assign mux_aoi_47_32_inst0_I[18] = config_reg_18_O;
assign mux_aoi_47_32_inst0_I[17] = config_reg_17_O;
assign mux_aoi_47_32_inst0_I[16] = config_reg_16_O;
assign mux_aoi_47_32_inst0_I[15] = config_reg_15_O;
assign mux_aoi_47_32_inst0_I[14] = config_reg_14_O;
assign mux_aoi_47_32_inst0_I[13] = config_reg_13_O;
assign mux_aoi_47_32_inst0_I[12] = config_reg_12_O;
assign mux_aoi_47_32_inst0_I[11] = config_reg_11_O;
assign mux_aoi_47_32_inst0_I[10] = config_reg_10_O;
assign mux_aoi_47_32_inst0_I[9] = config_reg_9_O;
assign mux_aoi_47_32_inst0_I[8] = config_reg_8_O;
assign mux_aoi_47_32_inst0_I[7] = config_reg_7_O;
assign mux_aoi_47_32_inst0_I[6] = config_reg_6_O;
assign mux_aoi_47_32_inst0_I[5] = config_reg_5_O;
assign mux_aoi_47_32_inst0_I[4] = config_reg_4_O;
assign mux_aoi_47_32_inst0_I[3] = config_reg_3_O;
assign mux_aoi_47_32_inst0_I[2] = config_reg_2_O;
assign mux_aoi_47_32_inst0_I[1] = config_reg_1_O;
assign mux_aoi_47_32_inst0_I[0] = config_reg_0_O;
mux_aoi_47_32 mux_aoi_47_32_inst0 (
    .I(mux_aoi_47_32_inst0_I),
    .O(mux_aoi_47_32_inst0_O),
    .S(self_config_config_addr_out[5:0]),
    .out_sel(mux_aoi_47_32_inst0_out_sel)
);
mantle_wire__typeBit8 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
SliceWrapper_25_24_25 tile_en_value (
    .I(config_reg_46_O),
    .O(tile_en_value_O)
);
assign MEM_input_width_17_num_0_ready = MemCore_inner_W_inst0_MEM_input_width_17_num_0_ready;
assign MEM_input_width_17_num_1_ready = MemCore_inner_W_inst0_MEM_input_width_17_num_1_ready;
assign MEM_input_width_17_num_2_ready = MemCore_inner_W_inst0_MEM_input_width_17_num_2_ready;
assign MEM_input_width_17_num_3_ready = MemCore_inner_W_inst0_MEM_input_width_17_num_3_ready;
assign MEM_input_width_1_num_0_ready = bit_const_1_None_out;
assign MEM_input_width_1_num_1_ready = bit_const_1_None_out;
assign MEM_output_width_17_num_0 = MemCore_inner_W_inst0_MEM_output_width_17_num_0;
assign MEM_output_width_17_num_0_valid = MemCore_inner_W_inst0_MEM_output_width_17_num_0_valid;
assign MEM_output_width_17_num_1 = MemCore_inner_W_inst0_MEM_output_width_17_num_1;
assign MEM_output_width_17_num_1_valid = MemCore_inner_W_inst0_MEM_output_width_17_num_1_valid;
assign MEM_output_width_17_num_2 = MemCore_inner_W_inst0_MEM_output_width_17_num_2;
assign MEM_output_width_17_num_2_valid = MemCore_inner_W_inst0_MEM_output_width_17_num_2_valid;
assign MEM_output_width_1_num_0 = MemCore_inner_W_inst0_MEM_output_width_1_num_0;
assign MEM_output_width_1_num_0_valid = bit_const_1_None_out;
assign MEM_output_width_1_num_1 = MemCore_inner_W_inst0_MEM_output_width_1_num_1;
assign MEM_output_width_1_num_1_valid = bit_const_1_None_out;
assign MEM_output_width_1_num_2 = MemCore_inner_W_inst0_MEM_output_width_1_num_2;
assign MEM_output_width_1_num_2_valid = bit_const_1_None_out;
assign read_config_data = mux_aoi_47_32_inst0_O;
assign read_config_data_1 = MemCore_inner_W_inst0_config_data_out_0;
assign read_config_data_2 = MemCore_inner_W_inst0_config_data_out_1;
endmodule

module CB_flush (
    input [0:0] I [19:0],
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output enable,
    output [31:0] out_sel,
    output [31:0] read_config_data,
    input ready_in,
    output ready_out,
    input reset,
    input [19:0] valid_in,
    output valid_out
);
wire [0:0] CB_flush_O;
wire CB_flush_ready_out;
wire CB_flush_valid_out;
wire [31:0] CB_flush_out_sel;
wire [0:0] CB_flush_enable_value_O;
wire [4:0] CB_flush_sel_value_O;
wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
wire [5:0] config_reg_0_O;
wire [0:0] CB_flush_I [19:0];
assign CB_flush_I[19] = I[19];
assign CB_flush_I[18] = I[18];
assign CB_flush_I[17] = I[17];
assign CB_flush_I[16] = I[16];
assign CB_flush_I[15] = I[15];
assign CB_flush_I[14] = I[14];
assign CB_flush_I[13] = I[13];
assign CB_flush_I[12] = I[12];
assign CB_flush_I[11] = I[11];
assign CB_flush_I[10] = I[10];
assign CB_flush_I[9] = I[9];
assign CB_flush_I[8] = I[8];
assign CB_flush_I[7] = I[7];
assign CB_flush_I[6] = I[6];
assign CB_flush_I[5] = I[5];
assign CB_flush_I[4] = I[4];
assign CB_flush_I[3] = I[3];
assign CB_flush_I[2] = I[2];
assign CB_flush_I[1] = I[1];
assign CB_flush_I[0] = I[0];
mux_aoi_ready_valid_const_20_1 CB_flush (
    .I(CB_flush_I),
    .O(CB_flush_O),
    .ready_in(ready_in),
    .ready_out(CB_flush_ready_out),
    .valid_in(valid_in),
    .valid_out(CB_flush_valid_out),
    .S(CB_flush_sel_value_O),
    .out_sel(CB_flush_out_sel)
);
SliceWrapper_6_0_1 CB_flush_enable_value (
    .I(config_reg_0_O),
    .O(CB_flush_enable_value_O)
);
SliceWrapper_6_1_6 CB_flush_sel_value (
    .I(config_reg_0_O),
    .O(CB_flush_sel_value_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_6_32_inst0$bit_const_0_None (
    .out(ZextWrapper_6_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O (
    .in(ZextWrapper_6_32_inst0$self_O_in),
    .out(ZextWrapper_6_32_inst0$self_O_out)
);
ConfigRegister_6_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_flush_O;
assign enable = CB_flush_enable_value_O[0];
assign out_sel = CB_flush_out_sel;
assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
assign ready_out = CB_flush_ready_out;
assign valid_out = CB_flush_valid_out;
endmodule

module CB_f2io_17 (
    output [16:0] O,
    input [16:0] I,
    input ready_in,
    output ready_out,
    input [0:0] valid_in,
    output valid_out,
    output [0:0] out_sel
);
wire [16:0] CB_f2io_17_O;
wire CB_f2io_17_ready_out;
wire CB_f2io_17_valid_out;
wire [0:0] const_0_1_out;
MuxWrapperAOI_1_17_ConstReadyValid CB_f2io_17 (
    .I(I),
    .O(CB_f2io_17_O),
    .ready_in(ready_in),
    .ready_out(CB_f2io_17_ready_out),
    .valid_in(valid_in[0]),
    .valid_out(CB_f2io_17_valid_out)
);
coreir_const #(
    .value(1'h0),
    .width(1)
) const_0_1 (
    .out(const_0_1_out)
);
assign O = CB_f2io_17_O;
assign ready_out = CB_f2io_17_ready_out;
assign valid_out = CB_f2io_17_valid_out;
assign out_sel = const_0_1_out;
endmodule

module CB_f2io_1 (
    output [0:0] O,
    input [0:0] I,
    input ready_in,
    output ready_out,
    input [0:0] valid_in,
    output valid_out,
    output [0:0] out_sel
);
wire [0:0] CB_f2io_1_O;
wire CB_f2io_1_ready_out;
wire CB_f2io_1_valid_out;
wire [0:0] const_0_1_out;
MuxWrapperAOI_1_1_ConstReadyValid CB_f2io_1 (
    .I(I),
    .O(CB_f2io_1_O),
    .ready_in(ready_in),
    .ready_out(CB_f2io_1_ready_out),
    .valid_in(valid_in[0]),
    .valid_out(CB_f2io_1_valid_out)
);
coreir_const #(
    .value(1'h0),
    .width(1)
) const_0_1 (
    .out(const_0_1_out)
);
assign O = CB_f2io_1_O;
assign ready_out = CB_f2io_1_ready_out;
assign valid_out = CB_f2io_1_valid_out;
assign out_sel = const_0_1_out;
endmodule

module Tile_IOCoreReadyValid (
    input clk,
    output clk_out,
    input [31:0] config_config_addr,
    input [31:0] config_config_data,
    output [31:0] config_out_config_addr,
    output [31:0] config_out_config_data,
    output [0:0] config_out_read,
    output [0:0] config_out_write,
    input [0:0] config_read,
    input [0:0] config_write,
    input [0:0] f2io_1,
    input [16:0] f2io_17,
    output f2io_17_ready,
    input f2io_17_valid,
    output f2io_1_ready,
    input f2io_1_valid,
    input [0:0] flush,
    output [0:0] flush_out,
    input [0:0] glb2io_1,
    input [16:0] glb2io_17,
    output glb2io_17_ready,
    input glb2io_17_valid,
    output glb2io_1_ready,
    input glb2io_1_valid,
    output [8:0] hi,
    output [0:0] io2f_1,
    output [16:0] io2f_17,
    input [4:0] io2f_17_ready,
    output io2f_17_valid,
    input [4:0] io2f_1_ready,
    output io2f_1_valid,
    output [0:0] io2glb_1,
    output [16:0] io2glb_17,
    input io2glb_17_ready,
    output io2glb_17_valid,
    input io2glb_1_ready,
    output io2glb_1_valid,
    output [7:0] lo,
    output [31:0] read_config_data,
    input [31:0] read_config_data_in,
    input reset,
    output reset_out,
    input [0:0] stall,
    output [0:0] stall_out,
    input [15:0] tile_id
);
wire [0:0] CB_f2io_1_O;
wire CB_f2io_1_ready_out;
wire CB_f2io_1_valid_out;
wire [0:0] CB_f2io_1_out_sel;
wire [16:0] CB_f2io_17_O;
wire CB_f2io_17_ready_out;
wire CB_f2io_17_valid_out;
wire [0:0] CB_f2io_17_out_sel;
wire DECODE_FEATURE_0_O;
wire DECODE_FEATURE_1_O;
wire DECODE_FEATURE_2_O;
wire DECODE_FEATURE_3_O;
wire DECODE_FEATURE_4_O;
wire DECODE_FEATURE_5_O;
wire FEATURE_AND_0_out;
wire FEATURE_AND_1_out;
wire FEATURE_AND_2_out;
wire FEATURE_AND_3_out;
wire FEATURE_AND_4_out;
wire FEATURE_AND_5_out;
wire [0:0] IOCoreReadyValid_inst0_f2io_17_ready;
wire [0:0] IOCoreReadyValid_inst0_f2io_1_ready;
wire [0:0] IOCoreReadyValid_inst0_glb2io_17_ready;
wire [0:0] IOCoreReadyValid_inst0_glb2io_1_ready;
wire [0:0] IOCoreReadyValid_inst0_io2f_1;
wire [16:0] IOCoreReadyValid_inst0_io2f_17;
wire [0:0] IOCoreReadyValid_inst0_io2f_17_valid;
wire [0:0] IOCoreReadyValid_inst0_io2f_1_valid;
wire [0:0] IOCoreReadyValid_inst0_io2glb_1;
wire [16:0] IOCoreReadyValid_inst0_io2glb_17;
wire [0:0] IOCoreReadyValid_inst0_io2glb_17_valid;
wire [0:0] IOCoreReadyValid_inst0_io2glb_1_valid;
wire [31:0] IOCoreReadyValid_inst0_read_config_data;
wire [0:0] PowerDomainConfigReg_inst0_ps_en_out;
wire [31:0] PowerDomainConfigReg_inst0_read_config_data;
wire [31:0] PowerDomainOR_O;
wire and_inst0_out;
wire and_inst1_out;
wire [31:0] const_0_32_out;
wire [7:0] const_0_8_out;
wire [8:0] const_511_9_out;
wire coreir_eq_16_inst0_out;
wire io2f_17_ready_merge$andr_inst0_out;
wire io2f_1_ready_merge$andr_inst0_out;
wire [31:0] read_data_mux_O;
wire [31:0] self_config_config_addr_out;
CB_f2io_1 CB_f2io_1 (
    .O(CB_f2io_1_O),
    .I(f2io_1),
    .ready_in(IOCoreReadyValid_inst0_f2io_1_ready[0]),
    .ready_out(CB_f2io_1_ready_out),
    .valid_in(f2io_1_valid),
    .valid_out(CB_f2io_1_valid_out),
    .out_sel(CB_f2io_1_out_sel)
);
CB_f2io_17 CB_f2io_17 (
    .O(CB_f2io_17_O),
    .I(f2io_17),
    .ready_in(IOCoreReadyValid_inst0_f2io_17_ready[0]),
    .ready_out(CB_f2io_17_ready_out),
    .valid_in(f2io_17_valid),
    .valid_out(CB_f2io_17_valid_out),
    .out_sel(CB_f2io_17_out_sel)
);
Decode08 DECODE_FEATURE_0 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_0_O)
);
Decode18 DECODE_FEATURE_1 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_1_O)
);
Decode28 DECODE_FEATURE_2 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_2_O)
);
Decode38 DECODE_FEATURE_3 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_3_O)
);
Decode48 DECODE_FEATURE_4 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_4_O)
);
Decode58 DECODE_FEATURE_5 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_5_O)
);
corebit_and FEATURE_AND_0 (
    .in0(DECODE_FEATURE_0_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_0_out)
);
corebit_and FEATURE_AND_1 (
    .in0(DECODE_FEATURE_1_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_1_out)
);
corebit_and FEATURE_AND_2 (
    .in0(DECODE_FEATURE_2_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_2_out)
);
corebit_and FEATURE_AND_3 (
    .in0(DECODE_FEATURE_3_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_3_out)
);
corebit_and FEATURE_AND_4 (
    .in0(DECODE_FEATURE_4_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_4_out)
);
corebit_and FEATURE_AND_5 (
    .in0(DECODE_FEATURE_5_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_5_out)
);
IOCoreReadyValid IOCoreReadyValid_inst0 (
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_0_out),
    .f2io_1(CB_f2io_1_O),
    .f2io_17(CB_f2io_17_O),
    .f2io_17_ready(IOCoreReadyValid_inst0_f2io_17_ready),
    .f2io_17_valid(CB_f2io_17_valid_out),
    .f2io_1_ready(IOCoreReadyValid_inst0_f2io_1_ready),
    .f2io_1_valid(CB_f2io_1_valid_out),
    .flush(flush),
    .flush_core(flush),
    .glb2io_1(glb2io_1),
    .glb2io_17(glb2io_17),
    .glb2io_17_ready(IOCoreReadyValid_inst0_glb2io_17_ready),
    .glb2io_17_valid(glb2io_17_valid),
    .glb2io_1_ready(IOCoreReadyValid_inst0_glb2io_1_ready),
    .glb2io_1_valid(glb2io_1_valid),
    .io2f_1(IOCoreReadyValid_inst0_io2f_1),
    .io2f_17(IOCoreReadyValid_inst0_io2f_17),
    .io2f_17_ready(io2f_17_ready_merge$andr_inst0_out),
    .io2f_17_valid(IOCoreReadyValid_inst0_io2f_17_valid),
    .io2f_1_ready(io2f_1_ready_merge$andr_inst0_out),
    .io2f_1_valid(IOCoreReadyValid_inst0_io2f_1_valid),
    .io2glb_1(IOCoreReadyValid_inst0_io2glb_1),
    .io2glb_17(IOCoreReadyValid_inst0_io2glb_17),
    .io2glb_17_ready(io2glb_17_ready),
    .io2glb_17_valid(IOCoreReadyValid_inst0_io2glb_17_valid),
    .io2glb_1_ready(io2glb_1_ready),
    .io2glb_1_valid(IOCoreReadyValid_inst0_io2glb_1_valid),
    .read_config_data(IOCoreReadyValid_inst0_read_config_data),
    .reset(reset),
    .stall(stall)
);
PowerDomainConfigReg PowerDomainConfigReg_inst0 (
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_5_out),
    .ps_en_out(PowerDomainConfigReg_inst0_ps_en_out),
    .read_config_data(PowerDomainConfigReg_inst0_read_config_data),
    .reset(reset)
);
PowerDomainOR PowerDomainOR (
    .I0(read_data_mux_O),
    .I1(read_config_data_in),
    .O(PowerDomainOR_O),
    .I_not(PowerDomainConfigReg_inst0_ps_en_out)
);
corebit_and and_inst0 (
    .in0(coreir_eq_16_inst0_out),
    .in1(config_read[0]),
    .out(and_inst0_out)
);
corebit_and and_inst1 (
    .in0(coreir_eq_16_inst0_out),
    .in1(config_write[0]),
    .out(and_inst1_out)
);
coreir_const #(
    .value(32'h00000000),
    .width(32)
) const_0_32 (
    .out(const_0_32_out)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
coreir_const #(
    .value(9'h1ff),
    .width(9)
) const_511_9 (
    .out(const_511_9_out)
);
coreir_eq #(
    .width(16)
) coreir_eq_16_inst0 (
    .in0(tile_id),
    .in1(self_config_config_addr_out[15:0]),
    .out(coreir_eq_16_inst0_out)
);
wire [4:0] io2f_17_ready_merge$andr_inst0_in;
assign io2f_17_ready_merge$andr_inst0_in = {io2f_17_ready[4],io2f_17_ready[3],io2f_17_ready[2],io2f_17_ready[1],io2f_17_ready[0]};
coreir_andr #(
    .width(5)
) io2f_17_ready_merge$andr_inst0 (
    .in(io2f_17_ready_merge$andr_inst0_in),
    .out(io2f_17_ready_merge$andr_inst0_out)
);
wire [4:0] io2f_1_ready_merge$andr_inst0_in;
assign io2f_1_ready_merge$andr_inst0_in = {io2f_1_ready[4],io2f_1_ready[3],io2f_1_ready[2],io2f_1_ready[1],io2f_1_ready[0]};
coreir_andr #(
    .width(5)
) io2f_1_ready_merge$andr_inst0 (
    .in(io2f_1_ready_merge$andr_inst0_in),
    .out(io2f_1_ready_merge$andr_inst0_out)
);
wire [31:0] read_data_mux_I [5:0];
assign read_data_mux_I[5] = PowerDomainConfigReg_inst0_read_config_data;
assign read_data_mux_I[4] = const_0_32_out;
assign read_data_mux_I[3] = const_0_32_out;
assign read_data_mux_I[2] = const_0_32_out;
assign read_data_mux_I[1] = const_0_32_out;
assign read_data_mux_I[0] = IOCoreReadyValid_inst0_read_config_data;
MuxWithDefaultWrapper_6_32_8_0 read_data_mux (
    .I(read_data_mux_I),
    .S(self_config_config_addr_out[23:16]),
    .EN(and_inst0_out),
    .O(read_data_mux_O)
);
mantle_wire__typeBit32 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
assign clk_out = clk;
assign config_out_config_addr = config_config_addr;
assign config_out_config_data = config_config_data;
assign config_out_read = config_read;
assign config_out_write = config_write;
assign f2io_17_ready = CB_f2io_17_ready_out;
assign f2io_1_ready = CB_f2io_1_ready_out;
assign flush_out = flush;
assign glb2io_17_ready = IOCoreReadyValid_inst0_glb2io_17_ready[0];
assign glb2io_1_ready = IOCoreReadyValid_inst0_glb2io_1_ready[0];
assign hi = const_511_9_out;
assign io2f_1 = IOCoreReadyValid_inst0_io2f_1;
assign io2f_17 = IOCoreReadyValid_inst0_io2f_17;
assign io2f_17_valid = IOCoreReadyValid_inst0_io2f_17_valid[0];
assign io2f_1_valid = IOCoreReadyValid_inst0_io2f_1_valid[0];
assign io2glb_1 = IOCoreReadyValid_inst0_io2glb_1;
assign io2glb_17 = IOCoreReadyValid_inst0_io2glb_17;
assign io2glb_17_valid = IOCoreReadyValid_inst0_io2glb_17_valid[0];
assign io2glb_1_valid = IOCoreReadyValid_inst0_io2glb_1_valid[0];
assign lo = const_0_8_out;
assign read_config_data = PowerDomainOR_O;
assign reset_out = reset;
assign stall_out = stall;
endmodule

module CB_PondTop_input_width_17_num_1 (
    input [16:0] I [20:0],
    output [16:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output enable,
    output [31:0] out_sel,
    output [31:0] read_config_data,
    input ready_in,
    output ready_out,
    input reset,
    input [20:0] valid_in,
    output valid_out
);
wire [16:0] CB_PondTop_input_width_17_num_1_O;
wire CB_PondTop_input_width_17_num_1_ready_out;
wire CB_PondTop_input_width_17_num_1_valid_out;
wire [31:0] CB_PondTop_input_width_17_num_1_out_sel;
wire [0:0] CB_PondTop_input_width_17_num_1_enable_value_O;
wire [4:0] CB_PondTop_input_width_17_num_1_sel_value_O;
wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
wire [5:0] config_reg_0_O;
wire [16:0] CB_PondTop_input_width_17_num_1_I [20:0];
assign CB_PondTop_input_width_17_num_1_I[20] = I[20];
assign CB_PondTop_input_width_17_num_1_I[19] = I[19];
assign CB_PondTop_input_width_17_num_1_I[18] = I[18];
assign CB_PondTop_input_width_17_num_1_I[17] = I[17];
assign CB_PondTop_input_width_17_num_1_I[16] = I[16];
assign CB_PondTop_input_width_17_num_1_I[15] = I[15];
assign CB_PondTop_input_width_17_num_1_I[14] = I[14];
assign CB_PondTop_input_width_17_num_1_I[13] = I[13];
assign CB_PondTop_input_width_17_num_1_I[12] = I[12];
assign CB_PondTop_input_width_17_num_1_I[11] = I[11];
assign CB_PondTop_input_width_17_num_1_I[10] = I[10];
assign CB_PondTop_input_width_17_num_1_I[9] = I[9];
assign CB_PondTop_input_width_17_num_1_I[8] = I[8];
assign CB_PondTop_input_width_17_num_1_I[7] = I[7];
assign CB_PondTop_input_width_17_num_1_I[6] = I[6];
assign CB_PondTop_input_width_17_num_1_I[5] = I[5];
assign CB_PondTop_input_width_17_num_1_I[4] = I[4];
assign CB_PondTop_input_width_17_num_1_I[3] = I[3];
assign CB_PondTop_input_width_17_num_1_I[2] = I[2];
assign CB_PondTop_input_width_17_num_1_I[1] = I[1];
assign CB_PondTop_input_width_17_num_1_I[0] = I[0];
mux_aoi_ready_valid_const_21_17 CB_PondTop_input_width_17_num_1 (
    .I(CB_PondTop_input_width_17_num_1_I),
    .O(CB_PondTop_input_width_17_num_1_O),
    .ready_in(ready_in),
    .ready_out(CB_PondTop_input_width_17_num_1_ready_out),
    .valid_in(valid_in),
    .valid_out(CB_PondTop_input_width_17_num_1_valid_out),
    .S(CB_PondTop_input_width_17_num_1_sel_value_O),
    .out_sel(CB_PondTop_input_width_17_num_1_out_sel)
);
SliceWrapper_6_0_1 CB_PondTop_input_width_17_num_1_enable_value (
    .I(config_reg_0_O),
    .O(CB_PondTop_input_width_17_num_1_enable_value_O)
);
SliceWrapper_6_1_6 CB_PondTop_input_width_17_num_1_sel_value (
    .I(config_reg_0_O),
    .O(CB_PondTop_input_width_17_num_1_sel_value_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_6_32_inst0$bit_const_0_None (
    .out(ZextWrapper_6_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O (
    .in(ZextWrapper_6_32_inst0$self_O_in),
    .out(ZextWrapper_6_32_inst0$self_O_out)
);
ConfigRegister_6_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_PondTop_input_width_17_num_1_O;
assign enable = CB_PondTop_input_width_17_num_1_enable_value_O[0];
assign out_sel = CB_PondTop_input_width_17_num_1_out_sel;
assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
assign ready_out = CB_PondTop_input_width_17_num_1_ready_out;
assign valid_out = CB_PondTop_input_width_17_num_1_valid_out;
endmodule

module CB_PondTop_input_width_17_num_0 (
    input [16:0] I [20:0],
    output [16:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output enable,
    output [31:0] out_sel,
    output [31:0] read_config_data,
    input ready_in,
    output ready_out,
    input reset,
    input [20:0] valid_in,
    output valid_out
);
wire [16:0] CB_PondTop_input_width_17_num_0_O;
wire CB_PondTop_input_width_17_num_0_ready_out;
wire CB_PondTop_input_width_17_num_0_valid_out;
wire [31:0] CB_PondTop_input_width_17_num_0_out_sel;
wire [0:0] CB_PondTop_input_width_17_num_0_enable_value_O;
wire [4:0] CB_PondTop_input_width_17_num_0_sel_value_O;
wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
wire [5:0] config_reg_0_O;
wire [16:0] CB_PondTop_input_width_17_num_0_I [20:0];
assign CB_PondTop_input_width_17_num_0_I[20] = I[20];
assign CB_PondTop_input_width_17_num_0_I[19] = I[19];
assign CB_PondTop_input_width_17_num_0_I[18] = I[18];
assign CB_PondTop_input_width_17_num_0_I[17] = I[17];
assign CB_PondTop_input_width_17_num_0_I[16] = I[16];
assign CB_PondTop_input_width_17_num_0_I[15] = I[15];
assign CB_PondTop_input_width_17_num_0_I[14] = I[14];
assign CB_PondTop_input_width_17_num_0_I[13] = I[13];
assign CB_PondTop_input_width_17_num_0_I[12] = I[12];
assign CB_PondTop_input_width_17_num_0_I[11] = I[11];
assign CB_PondTop_input_width_17_num_0_I[10] = I[10];
assign CB_PondTop_input_width_17_num_0_I[9] = I[9];
assign CB_PondTop_input_width_17_num_0_I[8] = I[8];
assign CB_PondTop_input_width_17_num_0_I[7] = I[7];
assign CB_PondTop_input_width_17_num_0_I[6] = I[6];
assign CB_PondTop_input_width_17_num_0_I[5] = I[5];
assign CB_PondTop_input_width_17_num_0_I[4] = I[4];
assign CB_PondTop_input_width_17_num_0_I[3] = I[3];
assign CB_PondTop_input_width_17_num_0_I[2] = I[2];
assign CB_PondTop_input_width_17_num_0_I[1] = I[1];
assign CB_PondTop_input_width_17_num_0_I[0] = I[0];
mux_aoi_ready_valid_const_21_17 CB_PondTop_input_width_17_num_0 (
    .I(CB_PondTop_input_width_17_num_0_I),
    .O(CB_PondTop_input_width_17_num_0_O),
    .ready_in(ready_in),
    .ready_out(CB_PondTop_input_width_17_num_0_ready_out),
    .valid_in(valid_in),
    .valid_out(CB_PondTop_input_width_17_num_0_valid_out),
    .S(CB_PondTop_input_width_17_num_0_sel_value_O),
    .out_sel(CB_PondTop_input_width_17_num_0_out_sel)
);
SliceWrapper_6_0_1 CB_PondTop_input_width_17_num_0_enable_value (
    .I(config_reg_0_O),
    .O(CB_PondTop_input_width_17_num_0_enable_value_O)
);
SliceWrapper_6_1_6 CB_PondTop_input_width_17_num_0_sel_value (
    .I(config_reg_0_O),
    .O(CB_PondTop_input_width_17_num_0_sel_value_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_6_32_inst0$bit_const_0_None (
    .out(ZextWrapper_6_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O (
    .in(ZextWrapper_6_32_inst0$self_O_in),
    .out(ZextWrapper_6_32_inst0$self_O_out)
);
ConfigRegister_6_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_PondTop_input_width_17_num_0_O;
assign enable = CB_PondTop_input_width_17_num_0_enable_value_O[0];
assign out_sel = CB_PondTop_input_width_17_num_0_out_sel;
assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
assign ready_out = CB_PondTop_input_width_17_num_0_ready_out;
assign valid_out = CB_PondTop_input_width_17_num_0_valid_out;
endmodule

module CB_PE_input_width_1_num_2 (
    input [0:0] I [19:0],
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output enable,
    output [31:0] out_sel,
    output [31:0] read_config_data,
    input ready_in,
    output ready_out,
    input reset,
    input [19:0] valid_in,
    output valid_out
);
wire [0:0] CB_PE_input_width_1_num_2_O;
wire CB_PE_input_width_1_num_2_ready_out;
wire CB_PE_input_width_1_num_2_valid_out;
wire [31:0] CB_PE_input_width_1_num_2_out_sel;
wire [0:0] CB_PE_input_width_1_num_2_enable_value_O;
wire [4:0] CB_PE_input_width_1_num_2_sel_value_O;
wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
wire [5:0] config_reg_0_O;
wire [0:0] CB_PE_input_width_1_num_2_I [19:0];
assign CB_PE_input_width_1_num_2_I[19] = I[19];
assign CB_PE_input_width_1_num_2_I[18] = I[18];
assign CB_PE_input_width_1_num_2_I[17] = I[17];
assign CB_PE_input_width_1_num_2_I[16] = I[16];
assign CB_PE_input_width_1_num_2_I[15] = I[15];
assign CB_PE_input_width_1_num_2_I[14] = I[14];
assign CB_PE_input_width_1_num_2_I[13] = I[13];
assign CB_PE_input_width_1_num_2_I[12] = I[12];
assign CB_PE_input_width_1_num_2_I[11] = I[11];
assign CB_PE_input_width_1_num_2_I[10] = I[10];
assign CB_PE_input_width_1_num_2_I[9] = I[9];
assign CB_PE_input_width_1_num_2_I[8] = I[8];
assign CB_PE_input_width_1_num_2_I[7] = I[7];
assign CB_PE_input_width_1_num_2_I[6] = I[6];
assign CB_PE_input_width_1_num_2_I[5] = I[5];
assign CB_PE_input_width_1_num_2_I[4] = I[4];
assign CB_PE_input_width_1_num_2_I[3] = I[3];
assign CB_PE_input_width_1_num_2_I[2] = I[2];
assign CB_PE_input_width_1_num_2_I[1] = I[1];
assign CB_PE_input_width_1_num_2_I[0] = I[0];
mux_aoi_ready_valid_const_20_1 CB_PE_input_width_1_num_2 (
    .I(CB_PE_input_width_1_num_2_I),
    .O(CB_PE_input_width_1_num_2_O),
    .ready_in(ready_in),
    .ready_out(CB_PE_input_width_1_num_2_ready_out),
    .valid_in(valid_in),
    .valid_out(CB_PE_input_width_1_num_2_valid_out),
    .S(CB_PE_input_width_1_num_2_sel_value_O),
    .out_sel(CB_PE_input_width_1_num_2_out_sel)
);
SliceWrapper_6_0_1 CB_PE_input_width_1_num_2_enable_value (
    .I(config_reg_0_O),
    .O(CB_PE_input_width_1_num_2_enable_value_O)
);
SliceWrapper_6_1_6 CB_PE_input_width_1_num_2_sel_value (
    .I(config_reg_0_O),
    .O(CB_PE_input_width_1_num_2_sel_value_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_6_32_inst0$bit_const_0_None (
    .out(ZextWrapper_6_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O (
    .in(ZextWrapper_6_32_inst0$self_O_in),
    .out(ZextWrapper_6_32_inst0$self_O_out)
);
ConfigRegister_6_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_PE_input_width_1_num_2_O;
assign enable = CB_PE_input_width_1_num_2_enable_value_O[0];
assign out_sel = CB_PE_input_width_1_num_2_out_sel;
assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
assign ready_out = CB_PE_input_width_1_num_2_ready_out;
assign valid_out = CB_PE_input_width_1_num_2_valid_out;
endmodule

module CB_PE_input_width_1_num_1 (
    input [0:0] I [19:0],
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output enable,
    output [31:0] out_sel,
    output [31:0] read_config_data,
    input ready_in,
    output ready_out,
    input reset,
    input [19:0] valid_in,
    output valid_out
);
wire [0:0] CB_PE_input_width_1_num_1_O;
wire CB_PE_input_width_1_num_1_ready_out;
wire CB_PE_input_width_1_num_1_valid_out;
wire [31:0] CB_PE_input_width_1_num_1_out_sel;
wire [0:0] CB_PE_input_width_1_num_1_enable_value_O;
wire [4:0] CB_PE_input_width_1_num_1_sel_value_O;
wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
wire [5:0] config_reg_0_O;
wire [0:0] CB_PE_input_width_1_num_1_I [19:0];
assign CB_PE_input_width_1_num_1_I[19] = I[19];
assign CB_PE_input_width_1_num_1_I[18] = I[18];
assign CB_PE_input_width_1_num_1_I[17] = I[17];
assign CB_PE_input_width_1_num_1_I[16] = I[16];
assign CB_PE_input_width_1_num_1_I[15] = I[15];
assign CB_PE_input_width_1_num_1_I[14] = I[14];
assign CB_PE_input_width_1_num_1_I[13] = I[13];
assign CB_PE_input_width_1_num_1_I[12] = I[12];
assign CB_PE_input_width_1_num_1_I[11] = I[11];
assign CB_PE_input_width_1_num_1_I[10] = I[10];
assign CB_PE_input_width_1_num_1_I[9] = I[9];
assign CB_PE_input_width_1_num_1_I[8] = I[8];
assign CB_PE_input_width_1_num_1_I[7] = I[7];
assign CB_PE_input_width_1_num_1_I[6] = I[6];
assign CB_PE_input_width_1_num_1_I[5] = I[5];
assign CB_PE_input_width_1_num_1_I[4] = I[4];
assign CB_PE_input_width_1_num_1_I[3] = I[3];
assign CB_PE_input_width_1_num_1_I[2] = I[2];
assign CB_PE_input_width_1_num_1_I[1] = I[1];
assign CB_PE_input_width_1_num_1_I[0] = I[0];
mux_aoi_ready_valid_const_20_1 CB_PE_input_width_1_num_1 (
    .I(CB_PE_input_width_1_num_1_I),
    .O(CB_PE_input_width_1_num_1_O),
    .ready_in(ready_in),
    .ready_out(CB_PE_input_width_1_num_1_ready_out),
    .valid_in(valid_in),
    .valid_out(CB_PE_input_width_1_num_1_valid_out),
    .S(CB_PE_input_width_1_num_1_sel_value_O),
    .out_sel(CB_PE_input_width_1_num_1_out_sel)
);
SliceWrapper_6_0_1 CB_PE_input_width_1_num_1_enable_value (
    .I(config_reg_0_O),
    .O(CB_PE_input_width_1_num_1_enable_value_O)
);
SliceWrapper_6_1_6 CB_PE_input_width_1_num_1_sel_value (
    .I(config_reg_0_O),
    .O(CB_PE_input_width_1_num_1_sel_value_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_6_32_inst0$bit_const_0_None (
    .out(ZextWrapper_6_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O (
    .in(ZextWrapper_6_32_inst0$self_O_in),
    .out(ZextWrapper_6_32_inst0$self_O_out)
);
ConfigRegister_6_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_PE_input_width_1_num_1_O;
assign enable = CB_PE_input_width_1_num_1_enable_value_O[0];
assign out_sel = CB_PE_input_width_1_num_1_out_sel;
assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
assign ready_out = CB_PE_input_width_1_num_1_ready_out;
assign valid_out = CB_PE_input_width_1_num_1_valid_out;
endmodule

module CB_PE_input_width_1_num_0 (
    input [0:0] I [20:0],
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output enable,
    output [31:0] out_sel,
    output [31:0] read_config_data,
    input ready_in,
    output ready_out,
    input reset,
    input [20:0] valid_in,
    output valid_out
);
wire [0:0] CB_PE_input_width_1_num_0_O;
wire CB_PE_input_width_1_num_0_ready_out;
wire CB_PE_input_width_1_num_0_valid_out;
wire [31:0] CB_PE_input_width_1_num_0_out_sel;
wire [0:0] CB_PE_input_width_1_num_0_enable_value_O;
wire [4:0] CB_PE_input_width_1_num_0_sel_value_O;
wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
wire [5:0] config_reg_0_O;
wire [0:0] CB_PE_input_width_1_num_0_I [20:0];
assign CB_PE_input_width_1_num_0_I[20] = I[20];
assign CB_PE_input_width_1_num_0_I[19] = I[19];
assign CB_PE_input_width_1_num_0_I[18] = I[18];
assign CB_PE_input_width_1_num_0_I[17] = I[17];
assign CB_PE_input_width_1_num_0_I[16] = I[16];
assign CB_PE_input_width_1_num_0_I[15] = I[15];
assign CB_PE_input_width_1_num_0_I[14] = I[14];
assign CB_PE_input_width_1_num_0_I[13] = I[13];
assign CB_PE_input_width_1_num_0_I[12] = I[12];
assign CB_PE_input_width_1_num_0_I[11] = I[11];
assign CB_PE_input_width_1_num_0_I[10] = I[10];
assign CB_PE_input_width_1_num_0_I[9] = I[9];
assign CB_PE_input_width_1_num_0_I[8] = I[8];
assign CB_PE_input_width_1_num_0_I[7] = I[7];
assign CB_PE_input_width_1_num_0_I[6] = I[6];
assign CB_PE_input_width_1_num_0_I[5] = I[5];
assign CB_PE_input_width_1_num_0_I[4] = I[4];
assign CB_PE_input_width_1_num_0_I[3] = I[3];
assign CB_PE_input_width_1_num_0_I[2] = I[2];
assign CB_PE_input_width_1_num_0_I[1] = I[1];
assign CB_PE_input_width_1_num_0_I[0] = I[0];
mux_aoi_ready_valid_const_21_1 CB_PE_input_width_1_num_0 (
    .I(CB_PE_input_width_1_num_0_I),
    .O(CB_PE_input_width_1_num_0_O),
    .ready_in(ready_in),
    .ready_out(CB_PE_input_width_1_num_0_ready_out),
    .valid_in(valid_in),
    .valid_out(CB_PE_input_width_1_num_0_valid_out),
    .S(CB_PE_input_width_1_num_0_sel_value_O),
    .out_sel(CB_PE_input_width_1_num_0_out_sel)
);
SliceWrapper_6_0_1 CB_PE_input_width_1_num_0_enable_value (
    .I(config_reg_0_O),
    .O(CB_PE_input_width_1_num_0_enable_value_O)
);
SliceWrapper_6_1_6 CB_PE_input_width_1_num_0_sel_value (
    .I(config_reg_0_O),
    .O(CB_PE_input_width_1_num_0_sel_value_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_6_32_inst0$bit_const_0_None (
    .out(ZextWrapper_6_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O (
    .in(ZextWrapper_6_32_inst0$self_O_in),
    .out(ZextWrapper_6_32_inst0$self_O_out)
);
ConfigRegister_6_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_PE_input_width_1_num_0_O;
assign enable = CB_PE_input_width_1_num_0_enable_value_O[0];
assign out_sel = CB_PE_input_width_1_num_0_out_sel;
assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
assign ready_out = CB_PE_input_width_1_num_0_ready_out;
assign valid_out = CB_PE_input_width_1_num_0_valid_out;
endmodule

module CB_PE_input_width_17_num_3 (
    input [16:0] I [19:0],
    output [16:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output enable,
    output [31:0] out_sel,
    output [31:0] read_config_data,
    input ready_in,
    output ready_out,
    input reset,
    input [19:0] valid_in,
    output valid_out
);
wire [16:0] CB_PE_input_width_17_num_3_O;
wire CB_PE_input_width_17_num_3_ready_out;
wire CB_PE_input_width_17_num_3_valid_out;
wire [31:0] CB_PE_input_width_17_num_3_out_sel;
wire [0:0] CB_PE_input_width_17_num_3_enable_value_O;
wire [4:0] CB_PE_input_width_17_num_3_sel_value_O;
wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
wire [5:0] config_reg_0_O;
wire [16:0] CB_PE_input_width_17_num_3_I [19:0];
assign CB_PE_input_width_17_num_3_I[19] = I[19];
assign CB_PE_input_width_17_num_3_I[18] = I[18];
assign CB_PE_input_width_17_num_3_I[17] = I[17];
assign CB_PE_input_width_17_num_3_I[16] = I[16];
assign CB_PE_input_width_17_num_3_I[15] = I[15];
assign CB_PE_input_width_17_num_3_I[14] = I[14];
assign CB_PE_input_width_17_num_3_I[13] = I[13];
assign CB_PE_input_width_17_num_3_I[12] = I[12];
assign CB_PE_input_width_17_num_3_I[11] = I[11];
assign CB_PE_input_width_17_num_3_I[10] = I[10];
assign CB_PE_input_width_17_num_3_I[9] = I[9];
assign CB_PE_input_width_17_num_3_I[8] = I[8];
assign CB_PE_input_width_17_num_3_I[7] = I[7];
assign CB_PE_input_width_17_num_3_I[6] = I[6];
assign CB_PE_input_width_17_num_3_I[5] = I[5];
assign CB_PE_input_width_17_num_3_I[4] = I[4];
assign CB_PE_input_width_17_num_3_I[3] = I[3];
assign CB_PE_input_width_17_num_3_I[2] = I[2];
assign CB_PE_input_width_17_num_3_I[1] = I[1];
assign CB_PE_input_width_17_num_3_I[0] = I[0];
mux_aoi_ready_valid_const_20_17 CB_PE_input_width_17_num_3 (
    .I(CB_PE_input_width_17_num_3_I),
    .O(CB_PE_input_width_17_num_3_O),
    .ready_in(ready_in),
    .ready_out(CB_PE_input_width_17_num_3_ready_out),
    .valid_in(valid_in),
    .valid_out(CB_PE_input_width_17_num_3_valid_out),
    .S(CB_PE_input_width_17_num_3_sel_value_O),
    .out_sel(CB_PE_input_width_17_num_3_out_sel)
);
SliceWrapper_6_0_1 CB_PE_input_width_17_num_3_enable_value (
    .I(config_reg_0_O),
    .O(CB_PE_input_width_17_num_3_enable_value_O)
);
SliceWrapper_6_1_6 CB_PE_input_width_17_num_3_sel_value (
    .I(config_reg_0_O),
    .O(CB_PE_input_width_17_num_3_sel_value_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_6_32_inst0$bit_const_0_None (
    .out(ZextWrapper_6_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O (
    .in(ZextWrapper_6_32_inst0$self_O_in),
    .out(ZextWrapper_6_32_inst0$self_O_out)
);
ConfigRegister_6_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_PE_input_width_17_num_3_O;
assign enable = CB_PE_input_width_17_num_3_enable_value_O[0];
assign out_sel = CB_PE_input_width_17_num_3_out_sel;
assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
assign ready_out = CB_PE_input_width_17_num_3_ready_out;
assign valid_out = CB_PE_input_width_17_num_3_valid_out;
endmodule

module CB_PE_input_width_17_num_2 (
    input [16:0] I [20:0],
    output [16:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output enable,
    output [31:0] out_sel,
    output [31:0] read_config_data,
    input ready_in,
    output ready_out,
    input reset,
    input [20:0] valid_in,
    output valid_out
);
wire [16:0] CB_PE_input_width_17_num_2_O;
wire CB_PE_input_width_17_num_2_ready_out;
wire CB_PE_input_width_17_num_2_valid_out;
wire [31:0] CB_PE_input_width_17_num_2_out_sel;
wire [0:0] CB_PE_input_width_17_num_2_enable_value_O;
wire [4:0] CB_PE_input_width_17_num_2_sel_value_O;
wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
wire [5:0] config_reg_0_O;
wire [16:0] CB_PE_input_width_17_num_2_I [20:0];
assign CB_PE_input_width_17_num_2_I[20] = I[20];
assign CB_PE_input_width_17_num_2_I[19] = I[19];
assign CB_PE_input_width_17_num_2_I[18] = I[18];
assign CB_PE_input_width_17_num_2_I[17] = I[17];
assign CB_PE_input_width_17_num_2_I[16] = I[16];
assign CB_PE_input_width_17_num_2_I[15] = I[15];
assign CB_PE_input_width_17_num_2_I[14] = I[14];
assign CB_PE_input_width_17_num_2_I[13] = I[13];
assign CB_PE_input_width_17_num_2_I[12] = I[12];
assign CB_PE_input_width_17_num_2_I[11] = I[11];
assign CB_PE_input_width_17_num_2_I[10] = I[10];
assign CB_PE_input_width_17_num_2_I[9] = I[9];
assign CB_PE_input_width_17_num_2_I[8] = I[8];
assign CB_PE_input_width_17_num_2_I[7] = I[7];
assign CB_PE_input_width_17_num_2_I[6] = I[6];
assign CB_PE_input_width_17_num_2_I[5] = I[5];
assign CB_PE_input_width_17_num_2_I[4] = I[4];
assign CB_PE_input_width_17_num_2_I[3] = I[3];
assign CB_PE_input_width_17_num_2_I[2] = I[2];
assign CB_PE_input_width_17_num_2_I[1] = I[1];
assign CB_PE_input_width_17_num_2_I[0] = I[0];
mux_aoi_ready_valid_const_21_17 CB_PE_input_width_17_num_2 (
    .I(CB_PE_input_width_17_num_2_I),
    .O(CB_PE_input_width_17_num_2_O),
    .ready_in(ready_in),
    .ready_out(CB_PE_input_width_17_num_2_ready_out),
    .valid_in(valid_in),
    .valid_out(CB_PE_input_width_17_num_2_valid_out),
    .S(CB_PE_input_width_17_num_2_sel_value_O),
    .out_sel(CB_PE_input_width_17_num_2_out_sel)
);
SliceWrapper_6_0_1 CB_PE_input_width_17_num_2_enable_value (
    .I(config_reg_0_O),
    .O(CB_PE_input_width_17_num_2_enable_value_O)
);
SliceWrapper_6_1_6 CB_PE_input_width_17_num_2_sel_value (
    .I(config_reg_0_O),
    .O(CB_PE_input_width_17_num_2_sel_value_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_6_32_inst0$bit_const_0_None (
    .out(ZextWrapper_6_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O (
    .in(ZextWrapper_6_32_inst0$self_O_in),
    .out(ZextWrapper_6_32_inst0$self_O_out)
);
ConfigRegister_6_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_PE_input_width_17_num_2_O;
assign enable = CB_PE_input_width_17_num_2_enable_value_O[0];
assign out_sel = CB_PE_input_width_17_num_2_out_sel;
assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
assign ready_out = CB_PE_input_width_17_num_2_ready_out;
assign valid_out = CB_PE_input_width_17_num_2_valid_out;
endmodule

module CB_PE_input_width_17_num_1 (
    input [16:0] I [20:0],
    output [16:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output enable,
    output [31:0] out_sel,
    output [31:0] read_config_data,
    input ready_in,
    output ready_out,
    input reset,
    input [20:0] valid_in,
    output valid_out
);
wire [16:0] CB_PE_input_width_17_num_1_O;
wire CB_PE_input_width_17_num_1_ready_out;
wire CB_PE_input_width_17_num_1_valid_out;
wire [31:0] CB_PE_input_width_17_num_1_out_sel;
wire [0:0] CB_PE_input_width_17_num_1_enable_value_O;
wire [4:0] CB_PE_input_width_17_num_1_sel_value_O;
wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
wire [5:0] config_reg_0_O;
wire [16:0] CB_PE_input_width_17_num_1_I [20:0];
assign CB_PE_input_width_17_num_1_I[20] = I[20];
assign CB_PE_input_width_17_num_1_I[19] = I[19];
assign CB_PE_input_width_17_num_1_I[18] = I[18];
assign CB_PE_input_width_17_num_1_I[17] = I[17];
assign CB_PE_input_width_17_num_1_I[16] = I[16];
assign CB_PE_input_width_17_num_1_I[15] = I[15];
assign CB_PE_input_width_17_num_1_I[14] = I[14];
assign CB_PE_input_width_17_num_1_I[13] = I[13];
assign CB_PE_input_width_17_num_1_I[12] = I[12];
assign CB_PE_input_width_17_num_1_I[11] = I[11];
assign CB_PE_input_width_17_num_1_I[10] = I[10];
assign CB_PE_input_width_17_num_1_I[9] = I[9];
assign CB_PE_input_width_17_num_1_I[8] = I[8];
assign CB_PE_input_width_17_num_1_I[7] = I[7];
assign CB_PE_input_width_17_num_1_I[6] = I[6];
assign CB_PE_input_width_17_num_1_I[5] = I[5];
assign CB_PE_input_width_17_num_1_I[4] = I[4];
assign CB_PE_input_width_17_num_1_I[3] = I[3];
assign CB_PE_input_width_17_num_1_I[2] = I[2];
assign CB_PE_input_width_17_num_1_I[1] = I[1];
assign CB_PE_input_width_17_num_1_I[0] = I[0];
mux_aoi_ready_valid_const_21_17 CB_PE_input_width_17_num_1 (
    .I(CB_PE_input_width_17_num_1_I),
    .O(CB_PE_input_width_17_num_1_O),
    .ready_in(ready_in),
    .ready_out(CB_PE_input_width_17_num_1_ready_out),
    .valid_in(valid_in),
    .valid_out(CB_PE_input_width_17_num_1_valid_out),
    .S(CB_PE_input_width_17_num_1_sel_value_O),
    .out_sel(CB_PE_input_width_17_num_1_out_sel)
);
SliceWrapper_6_0_1 CB_PE_input_width_17_num_1_enable_value (
    .I(config_reg_0_O),
    .O(CB_PE_input_width_17_num_1_enable_value_O)
);
SliceWrapper_6_1_6 CB_PE_input_width_17_num_1_sel_value (
    .I(config_reg_0_O),
    .O(CB_PE_input_width_17_num_1_sel_value_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_6_32_inst0$bit_const_0_None (
    .out(ZextWrapper_6_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O (
    .in(ZextWrapper_6_32_inst0$self_O_in),
    .out(ZextWrapper_6_32_inst0$self_O_out)
);
ConfigRegister_6_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_PE_input_width_17_num_1_O;
assign enable = CB_PE_input_width_17_num_1_enable_value_O[0];
assign out_sel = CB_PE_input_width_17_num_1_out_sel;
assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
assign ready_out = CB_PE_input_width_17_num_1_ready_out;
assign valid_out = CB_PE_input_width_17_num_1_valid_out;
endmodule

module CB_PE_input_width_17_num_0 (
    input [16:0] I [20:0],
    output [16:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output enable,
    output [31:0] out_sel,
    output [31:0] read_config_data,
    input ready_in,
    output ready_out,
    input reset,
    input [20:0] valid_in,
    output valid_out
);
wire [16:0] CB_PE_input_width_17_num_0_O;
wire CB_PE_input_width_17_num_0_ready_out;
wire CB_PE_input_width_17_num_0_valid_out;
wire [31:0] CB_PE_input_width_17_num_0_out_sel;
wire [0:0] CB_PE_input_width_17_num_0_enable_value_O;
wire [4:0] CB_PE_input_width_17_num_0_sel_value_O;
wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
wire [5:0] config_reg_0_O;
wire [16:0] CB_PE_input_width_17_num_0_I [20:0];
assign CB_PE_input_width_17_num_0_I[20] = I[20];
assign CB_PE_input_width_17_num_0_I[19] = I[19];
assign CB_PE_input_width_17_num_0_I[18] = I[18];
assign CB_PE_input_width_17_num_0_I[17] = I[17];
assign CB_PE_input_width_17_num_0_I[16] = I[16];
assign CB_PE_input_width_17_num_0_I[15] = I[15];
assign CB_PE_input_width_17_num_0_I[14] = I[14];
assign CB_PE_input_width_17_num_0_I[13] = I[13];
assign CB_PE_input_width_17_num_0_I[12] = I[12];
assign CB_PE_input_width_17_num_0_I[11] = I[11];
assign CB_PE_input_width_17_num_0_I[10] = I[10];
assign CB_PE_input_width_17_num_0_I[9] = I[9];
assign CB_PE_input_width_17_num_0_I[8] = I[8];
assign CB_PE_input_width_17_num_0_I[7] = I[7];
assign CB_PE_input_width_17_num_0_I[6] = I[6];
assign CB_PE_input_width_17_num_0_I[5] = I[5];
assign CB_PE_input_width_17_num_0_I[4] = I[4];
assign CB_PE_input_width_17_num_0_I[3] = I[3];
assign CB_PE_input_width_17_num_0_I[2] = I[2];
assign CB_PE_input_width_17_num_0_I[1] = I[1];
assign CB_PE_input_width_17_num_0_I[0] = I[0];
mux_aoi_ready_valid_const_21_17 CB_PE_input_width_17_num_0 (
    .I(CB_PE_input_width_17_num_0_I),
    .O(CB_PE_input_width_17_num_0_O),
    .ready_in(ready_in),
    .ready_out(CB_PE_input_width_17_num_0_ready_out),
    .valid_in(valid_in),
    .valid_out(CB_PE_input_width_17_num_0_valid_out),
    .S(CB_PE_input_width_17_num_0_sel_value_O),
    .out_sel(CB_PE_input_width_17_num_0_out_sel)
);
SliceWrapper_6_0_1 CB_PE_input_width_17_num_0_enable_value (
    .I(config_reg_0_O),
    .O(CB_PE_input_width_17_num_0_enable_value_O)
);
SliceWrapper_6_1_6 CB_PE_input_width_17_num_0_sel_value (
    .I(config_reg_0_O),
    .O(CB_PE_input_width_17_num_0_sel_value_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_6_32_inst0$bit_const_0_None (
    .out(ZextWrapper_6_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O (
    .in(ZextWrapper_6_32_inst0$self_O_in),
    .out(ZextWrapper_6_32_inst0$self_O_out)
);
ConfigRegister_6_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_PE_input_width_17_num_0_O;
assign enable = CB_PE_input_width_17_num_0_enable_value_O[0];
assign out_sel = CB_PE_input_width_17_num_0_out_sel;
assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
assign ready_out = CB_PE_input_width_17_num_0_ready_out;
assign valid_out = CB_PE_input_width_17_num_0_valid_out;
endmodule

module Tile_PE (
    input [0:0] SB_T0_EAST_SB_IN_B1,
    input [16:0] SB_T0_EAST_SB_IN_B17,
    output SB_T0_EAST_SB_IN_B17_ready,
    input SB_T0_EAST_SB_IN_B17_valid,
    output SB_T0_EAST_SB_IN_B1_ready,
    input SB_T0_EAST_SB_IN_B1_valid,
    output [0:0] SB_T0_EAST_SB_OUT_B1,
    output [16:0] SB_T0_EAST_SB_OUT_B17,
    input SB_T0_EAST_SB_OUT_B17_ready,
    output SB_T0_EAST_SB_OUT_B17_valid,
    input SB_T0_EAST_SB_OUT_B1_ready,
    output SB_T0_EAST_SB_OUT_B1_valid,
    input [0:0] SB_T0_NORTH_SB_IN_B1,
    input [16:0] SB_T0_NORTH_SB_IN_B17,
    output SB_T0_NORTH_SB_IN_B17_ready,
    input SB_T0_NORTH_SB_IN_B17_valid,
    output SB_T0_NORTH_SB_IN_B1_ready,
    input SB_T0_NORTH_SB_IN_B1_valid,
    output [0:0] SB_T0_NORTH_SB_OUT_B1,
    output [16:0] SB_T0_NORTH_SB_OUT_B17,
    input SB_T0_NORTH_SB_OUT_B17_ready,
    output SB_T0_NORTH_SB_OUT_B17_valid,
    input SB_T0_NORTH_SB_OUT_B1_ready,
    output SB_T0_NORTH_SB_OUT_B1_valid,
    input [0:0] SB_T0_SOUTH_SB_IN_B1,
    input [16:0] SB_T0_SOUTH_SB_IN_B17,
    output SB_T0_SOUTH_SB_IN_B17_ready,
    input SB_T0_SOUTH_SB_IN_B17_valid,
    output SB_T0_SOUTH_SB_IN_B1_ready,
    input SB_T0_SOUTH_SB_IN_B1_valid,
    output [0:0] SB_T0_SOUTH_SB_OUT_B1,
    output [16:0] SB_T0_SOUTH_SB_OUT_B17,
    input SB_T0_SOUTH_SB_OUT_B17_ready,
    output SB_T0_SOUTH_SB_OUT_B17_valid,
    input SB_T0_SOUTH_SB_OUT_B1_ready,
    output SB_T0_SOUTH_SB_OUT_B1_valid,
    input [0:0] SB_T0_WEST_SB_IN_B1,
    input [16:0] SB_T0_WEST_SB_IN_B17,
    output SB_T0_WEST_SB_IN_B17_ready,
    input SB_T0_WEST_SB_IN_B17_valid,
    output SB_T0_WEST_SB_IN_B1_ready,
    input SB_T0_WEST_SB_IN_B1_valid,
    output [0:0] SB_T0_WEST_SB_OUT_B1,
    output [16:0] SB_T0_WEST_SB_OUT_B17,
    input SB_T0_WEST_SB_OUT_B17_ready,
    output SB_T0_WEST_SB_OUT_B17_valid,
    input SB_T0_WEST_SB_OUT_B1_ready,
    output SB_T0_WEST_SB_OUT_B1_valid,
    input [0:0] SB_T1_EAST_SB_IN_B1,
    input [16:0] SB_T1_EAST_SB_IN_B17,
    output SB_T1_EAST_SB_IN_B17_ready,
    input SB_T1_EAST_SB_IN_B17_valid,
    output SB_T1_EAST_SB_IN_B1_ready,
    input SB_T1_EAST_SB_IN_B1_valid,
    output [0:0] SB_T1_EAST_SB_OUT_B1,
    output [16:0] SB_T1_EAST_SB_OUT_B17,
    input SB_T1_EAST_SB_OUT_B17_ready,
    output SB_T1_EAST_SB_OUT_B17_valid,
    input SB_T1_EAST_SB_OUT_B1_ready,
    output SB_T1_EAST_SB_OUT_B1_valid,
    input [0:0] SB_T1_NORTH_SB_IN_B1,
    input [16:0] SB_T1_NORTH_SB_IN_B17,
    output SB_T1_NORTH_SB_IN_B17_ready,
    input SB_T1_NORTH_SB_IN_B17_valid,
    output SB_T1_NORTH_SB_IN_B1_ready,
    input SB_T1_NORTH_SB_IN_B1_valid,
    output [0:0] SB_T1_NORTH_SB_OUT_B1,
    output [16:0] SB_T1_NORTH_SB_OUT_B17,
    input SB_T1_NORTH_SB_OUT_B17_ready,
    output SB_T1_NORTH_SB_OUT_B17_valid,
    input SB_T1_NORTH_SB_OUT_B1_ready,
    output SB_T1_NORTH_SB_OUT_B1_valid,
    input [0:0] SB_T1_SOUTH_SB_IN_B1,
    input [16:0] SB_T1_SOUTH_SB_IN_B17,
    output SB_T1_SOUTH_SB_IN_B17_ready,
    input SB_T1_SOUTH_SB_IN_B17_valid,
    output SB_T1_SOUTH_SB_IN_B1_ready,
    input SB_T1_SOUTH_SB_IN_B1_valid,
    output [0:0] SB_T1_SOUTH_SB_OUT_B1,
    output [16:0] SB_T1_SOUTH_SB_OUT_B17,
    input SB_T1_SOUTH_SB_OUT_B17_ready,
    output SB_T1_SOUTH_SB_OUT_B17_valid,
    input SB_T1_SOUTH_SB_OUT_B1_ready,
    output SB_T1_SOUTH_SB_OUT_B1_valid,
    input [0:0] SB_T1_WEST_SB_IN_B1,
    input [16:0] SB_T1_WEST_SB_IN_B17,
    output SB_T1_WEST_SB_IN_B17_ready,
    input SB_T1_WEST_SB_IN_B17_valid,
    output SB_T1_WEST_SB_IN_B1_ready,
    input SB_T1_WEST_SB_IN_B1_valid,
    output [0:0] SB_T1_WEST_SB_OUT_B1,
    output [16:0] SB_T1_WEST_SB_OUT_B17,
    input SB_T1_WEST_SB_OUT_B17_ready,
    output SB_T1_WEST_SB_OUT_B17_valid,
    input SB_T1_WEST_SB_OUT_B1_ready,
    output SB_T1_WEST_SB_OUT_B1_valid,
    input [0:0] SB_T2_EAST_SB_IN_B1,
    input [16:0] SB_T2_EAST_SB_IN_B17,
    output SB_T2_EAST_SB_IN_B17_ready,
    input SB_T2_EAST_SB_IN_B17_valid,
    output SB_T2_EAST_SB_IN_B1_ready,
    input SB_T2_EAST_SB_IN_B1_valid,
    output [0:0] SB_T2_EAST_SB_OUT_B1,
    output [16:0] SB_T2_EAST_SB_OUT_B17,
    input SB_T2_EAST_SB_OUT_B17_ready,
    output SB_T2_EAST_SB_OUT_B17_valid,
    input SB_T2_EAST_SB_OUT_B1_ready,
    output SB_T2_EAST_SB_OUT_B1_valid,
    input [0:0] SB_T2_NORTH_SB_IN_B1,
    input [16:0] SB_T2_NORTH_SB_IN_B17,
    output SB_T2_NORTH_SB_IN_B17_ready,
    input SB_T2_NORTH_SB_IN_B17_valid,
    output SB_T2_NORTH_SB_IN_B1_ready,
    input SB_T2_NORTH_SB_IN_B1_valid,
    output [0:0] SB_T2_NORTH_SB_OUT_B1,
    output [16:0] SB_T2_NORTH_SB_OUT_B17,
    input SB_T2_NORTH_SB_OUT_B17_ready,
    output SB_T2_NORTH_SB_OUT_B17_valid,
    input SB_T2_NORTH_SB_OUT_B1_ready,
    output SB_T2_NORTH_SB_OUT_B1_valid,
    input [0:0] SB_T2_SOUTH_SB_IN_B1,
    input [16:0] SB_T2_SOUTH_SB_IN_B17,
    output SB_T2_SOUTH_SB_IN_B17_ready,
    input SB_T2_SOUTH_SB_IN_B17_valid,
    output SB_T2_SOUTH_SB_IN_B1_ready,
    input SB_T2_SOUTH_SB_IN_B1_valid,
    output [0:0] SB_T2_SOUTH_SB_OUT_B1,
    output [16:0] SB_T2_SOUTH_SB_OUT_B17,
    input SB_T2_SOUTH_SB_OUT_B17_ready,
    output SB_T2_SOUTH_SB_OUT_B17_valid,
    input SB_T2_SOUTH_SB_OUT_B1_ready,
    output SB_T2_SOUTH_SB_OUT_B1_valid,
    input [0:0] SB_T2_WEST_SB_IN_B1,
    input [16:0] SB_T2_WEST_SB_IN_B17,
    output SB_T2_WEST_SB_IN_B17_ready,
    input SB_T2_WEST_SB_IN_B17_valid,
    output SB_T2_WEST_SB_IN_B1_ready,
    input SB_T2_WEST_SB_IN_B1_valid,
    output [0:0] SB_T2_WEST_SB_OUT_B1,
    output [16:0] SB_T2_WEST_SB_OUT_B17,
    input SB_T2_WEST_SB_OUT_B17_ready,
    output SB_T2_WEST_SB_OUT_B17_valid,
    input SB_T2_WEST_SB_OUT_B1_ready,
    output SB_T2_WEST_SB_OUT_B1_valid,
    input [0:0] SB_T3_EAST_SB_IN_B1,
    input [16:0] SB_T3_EAST_SB_IN_B17,
    output SB_T3_EAST_SB_IN_B17_ready,
    input SB_T3_EAST_SB_IN_B17_valid,
    output SB_T3_EAST_SB_IN_B1_ready,
    input SB_T3_EAST_SB_IN_B1_valid,
    output [0:0] SB_T3_EAST_SB_OUT_B1,
    output [16:0] SB_T3_EAST_SB_OUT_B17,
    input SB_T3_EAST_SB_OUT_B17_ready,
    output SB_T3_EAST_SB_OUT_B17_valid,
    input SB_T3_EAST_SB_OUT_B1_ready,
    output SB_T3_EAST_SB_OUT_B1_valid,
    input [0:0] SB_T3_NORTH_SB_IN_B1,
    input [16:0] SB_T3_NORTH_SB_IN_B17,
    output SB_T3_NORTH_SB_IN_B17_ready,
    input SB_T3_NORTH_SB_IN_B17_valid,
    output SB_T3_NORTH_SB_IN_B1_ready,
    input SB_T3_NORTH_SB_IN_B1_valid,
    output [0:0] SB_T3_NORTH_SB_OUT_B1,
    output [16:0] SB_T3_NORTH_SB_OUT_B17,
    input SB_T3_NORTH_SB_OUT_B17_ready,
    output SB_T3_NORTH_SB_OUT_B17_valid,
    input SB_T3_NORTH_SB_OUT_B1_ready,
    output SB_T3_NORTH_SB_OUT_B1_valid,
    input [0:0] SB_T3_SOUTH_SB_IN_B1,
    input [16:0] SB_T3_SOUTH_SB_IN_B17,
    output SB_T3_SOUTH_SB_IN_B17_ready,
    input SB_T3_SOUTH_SB_IN_B17_valid,
    output SB_T3_SOUTH_SB_IN_B1_ready,
    input SB_T3_SOUTH_SB_IN_B1_valid,
    output [0:0] SB_T3_SOUTH_SB_OUT_B1,
    output [16:0] SB_T3_SOUTH_SB_OUT_B17,
    input SB_T3_SOUTH_SB_OUT_B17_ready,
    output SB_T3_SOUTH_SB_OUT_B17_valid,
    input SB_T3_SOUTH_SB_OUT_B1_ready,
    output SB_T3_SOUTH_SB_OUT_B1_valid,
    input [0:0] SB_T3_WEST_SB_IN_B1,
    input [16:0] SB_T3_WEST_SB_IN_B17,
    output SB_T3_WEST_SB_IN_B17_ready,
    input SB_T3_WEST_SB_IN_B17_valid,
    output SB_T3_WEST_SB_IN_B1_ready,
    input SB_T3_WEST_SB_IN_B1_valid,
    output [0:0] SB_T3_WEST_SB_OUT_B1,
    output [16:0] SB_T3_WEST_SB_OUT_B17,
    input SB_T3_WEST_SB_OUT_B17_ready,
    output SB_T3_WEST_SB_OUT_B17_valid,
    input SB_T3_WEST_SB_OUT_B1_ready,
    output SB_T3_WEST_SB_OUT_B1_valid,
    input [0:0] SB_T4_EAST_SB_IN_B1,
    input [16:0] SB_T4_EAST_SB_IN_B17,
    output SB_T4_EAST_SB_IN_B17_ready,
    input SB_T4_EAST_SB_IN_B17_valid,
    output SB_T4_EAST_SB_IN_B1_ready,
    input SB_T4_EAST_SB_IN_B1_valid,
    output [0:0] SB_T4_EAST_SB_OUT_B1,
    output [16:0] SB_T4_EAST_SB_OUT_B17,
    input SB_T4_EAST_SB_OUT_B17_ready,
    output SB_T4_EAST_SB_OUT_B17_valid,
    input SB_T4_EAST_SB_OUT_B1_ready,
    output SB_T4_EAST_SB_OUT_B1_valid,
    input [0:0] SB_T4_NORTH_SB_IN_B1,
    input [16:0] SB_T4_NORTH_SB_IN_B17,
    output SB_T4_NORTH_SB_IN_B17_ready,
    input SB_T4_NORTH_SB_IN_B17_valid,
    output SB_T4_NORTH_SB_IN_B1_ready,
    input SB_T4_NORTH_SB_IN_B1_valid,
    output [0:0] SB_T4_NORTH_SB_OUT_B1,
    output [16:0] SB_T4_NORTH_SB_OUT_B17,
    input SB_T4_NORTH_SB_OUT_B17_ready,
    output SB_T4_NORTH_SB_OUT_B17_valid,
    input SB_T4_NORTH_SB_OUT_B1_ready,
    output SB_T4_NORTH_SB_OUT_B1_valid,
    input [0:0] SB_T4_SOUTH_SB_IN_B1,
    input [16:0] SB_T4_SOUTH_SB_IN_B17,
    output SB_T4_SOUTH_SB_IN_B17_ready,
    input SB_T4_SOUTH_SB_IN_B17_valid,
    output SB_T4_SOUTH_SB_IN_B1_ready,
    input SB_T4_SOUTH_SB_IN_B1_valid,
    output [0:0] SB_T4_SOUTH_SB_OUT_B1,
    output [16:0] SB_T4_SOUTH_SB_OUT_B17,
    input SB_T4_SOUTH_SB_OUT_B17_ready,
    output SB_T4_SOUTH_SB_OUT_B17_valid,
    input SB_T4_SOUTH_SB_OUT_B1_ready,
    output SB_T4_SOUTH_SB_OUT_B1_valid,
    input [0:0] SB_T4_WEST_SB_IN_B1,
    input [16:0] SB_T4_WEST_SB_IN_B17,
    output SB_T4_WEST_SB_IN_B17_ready,
    input SB_T4_WEST_SB_IN_B17_valid,
    output SB_T4_WEST_SB_IN_B1_ready,
    input SB_T4_WEST_SB_IN_B1_valid,
    output [0:0] SB_T4_WEST_SB_OUT_B1,
    output [16:0] SB_T4_WEST_SB_OUT_B17,
    input SB_T4_WEST_SB_OUT_B17_ready,
    output SB_T4_WEST_SB_OUT_B17_valid,
    input SB_T4_WEST_SB_OUT_B1_ready,
    output SB_T4_WEST_SB_OUT_B1_valid,
    input clk,
    output clk_out,
    input clk_pass_through,
    output clk_pass_through_out_bot,
    output clk_pass_through_out_right,
    input [31:0] config_config_addr,
    input [31:0] config_config_data,
    output [31:0] config_out_config_addr,
    output [31:0] config_out_config_data,
    output [0:0] config_out_read,
    output [0:0] config_out_write,
    input [0:0] config_read,
    input [0:0] config_write,
    input [0:0] flush,
    output [0:0] flush_out,
    output [8:0] hi,
    output [7:0] lo,
    output [31:0] read_config_data,
    input [31:0] read_config_data_in,
    input reset,
    output reset_out,
    input [0:0] stall,
    output [0:0] stall_out,
    input [15:0] tile_id
);
wire [16:0] CB_PE_input_width_17_num_0_O;
wire CB_PE_input_width_17_num_0_enable;
wire [31:0] CB_PE_input_width_17_num_0_out_sel;
wire [31:0] CB_PE_input_width_17_num_0_read_config_data;
wire CB_PE_input_width_17_num_0_ready_out;
wire CB_PE_input_width_17_num_0_valid_out;
wire [16:0] CB_PE_input_width_17_num_1_O;
wire CB_PE_input_width_17_num_1_enable;
wire [31:0] CB_PE_input_width_17_num_1_out_sel;
wire [31:0] CB_PE_input_width_17_num_1_read_config_data;
wire CB_PE_input_width_17_num_1_ready_out;
wire CB_PE_input_width_17_num_1_valid_out;
wire [16:0] CB_PE_input_width_17_num_2_O;
wire CB_PE_input_width_17_num_2_enable;
wire [31:0] CB_PE_input_width_17_num_2_out_sel;
wire [31:0] CB_PE_input_width_17_num_2_read_config_data;
wire CB_PE_input_width_17_num_2_ready_out;
wire CB_PE_input_width_17_num_2_valid_out;
wire [16:0] CB_PE_input_width_17_num_3_O;
wire CB_PE_input_width_17_num_3_enable;
wire [31:0] CB_PE_input_width_17_num_3_out_sel;
wire [31:0] CB_PE_input_width_17_num_3_read_config_data;
wire CB_PE_input_width_17_num_3_ready_out;
wire CB_PE_input_width_17_num_3_valid_out;
wire [0:0] CB_PE_input_width_1_num_0_O;
wire CB_PE_input_width_1_num_0_enable;
wire [31:0] CB_PE_input_width_1_num_0_out_sel;
wire [31:0] CB_PE_input_width_1_num_0_read_config_data;
wire CB_PE_input_width_1_num_0_ready_out;
wire CB_PE_input_width_1_num_0_valid_out;
wire [0:0] CB_PE_input_width_1_num_1_O;
wire CB_PE_input_width_1_num_1_enable;
wire [31:0] CB_PE_input_width_1_num_1_out_sel;
wire [31:0] CB_PE_input_width_1_num_1_read_config_data;
wire CB_PE_input_width_1_num_1_ready_out;
wire CB_PE_input_width_1_num_1_valid_out;
wire [0:0] CB_PE_input_width_1_num_2_O;
wire CB_PE_input_width_1_num_2_enable;
wire [31:0] CB_PE_input_width_1_num_2_out_sel;
wire [31:0] CB_PE_input_width_1_num_2_read_config_data;
wire CB_PE_input_width_1_num_2_ready_out;
wire CB_PE_input_width_1_num_2_valid_out;
wire [16:0] CB_PondTop_input_width_17_num_0_O;
wire CB_PondTop_input_width_17_num_0_enable;
wire [31:0] CB_PondTop_input_width_17_num_0_out_sel;
wire [31:0] CB_PondTop_input_width_17_num_0_read_config_data;
wire CB_PondTop_input_width_17_num_0_ready_out;
wire CB_PondTop_input_width_17_num_0_valid_out;
wire [16:0] CB_PondTop_input_width_17_num_1_O;
wire CB_PondTop_input_width_17_num_1_enable;
wire [31:0] CB_PondTop_input_width_17_num_1_out_sel;
wire [31:0] CB_PondTop_input_width_17_num_1_read_config_data;
wire CB_PondTop_input_width_17_num_1_ready_out;
wire CB_PondTop_input_width_17_num_1_valid_out;
wire [0:0] CB_flush_O;
wire CB_flush_enable;
wire [31:0] CB_flush_out_sel;
wire [31:0] CB_flush_read_config_data;
wire CB_flush_ready_out;
wire CB_flush_valid_out;
wire DECODE_FEATURE_0_O;
wire DECODE_FEATURE_1_O;
wire DECODE_FEATURE_10_O;
wire DECODE_FEATURE_11_O;
wire DECODE_FEATURE_12_O;
wire DECODE_FEATURE_13_O;
wire DECODE_FEATURE_14_O;
wire DECODE_FEATURE_15_O;
wire DECODE_FEATURE_2_O;
wire DECODE_FEATURE_3_O;
wire DECODE_FEATURE_4_O;
wire DECODE_FEATURE_5_O;
wire DECODE_FEATURE_6_O;
wire DECODE_FEATURE_7_O;
wire DECODE_FEATURE_8_O;
wire DECODE_FEATURE_9_O;
wire FEATURE_AND_0_out;
wire FEATURE_AND_1_out;
wire FEATURE_AND_10_out;
wire FEATURE_AND_11_out;
wire FEATURE_AND_12_out;
wire FEATURE_AND_13_out;
wire FEATURE_AND_14_out;
wire FEATURE_AND_15_out;
wire FEATURE_AND_2_out;
wire FEATURE_AND_3_out;
wire FEATURE_AND_4_out;
wire FEATURE_AND_5_out;
wire FEATURE_AND_6_out;
wire FEATURE_AND_7_out;
wire FEATURE_AND_8_out;
wire FEATURE_AND_9_out;
wire [0:0] PE_inst0_PE_input_width_17_num_0_ready;
wire [0:0] PE_inst0_PE_input_width_17_num_1_ready;
wire [0:0] PE_inst0_PE_input_width_17_num_2_ready;
wire [0:0] PE_inst0_PE_input_width_17_num_3_ready;
wire PE_inst0_PE_input_width_1_num_0_ready;
wire PE_inst0_PE_input_width_1_num_1_ready;
wire PE_inst0_PE_input_width_1_num_2_ready;
wire [16:0] PE_inst0_PE_output_width_17_num_0;
wire [0:0] PE_inst0_PE_output_width_17_num_0_valid;
wire [16:0] PE_inst0_PE_output_width_17_num_1;
wire [0:0] PE_inst0_PE_output_width_17_num_1_valid;
wire [16:0] PE_inst0_PE_output_width_17_num_2;
wire [0:0] PE_inst0_PE_output_width_17_num_2_valid;
wire [0:0] PE_inst0_PE_output_width_1_num_0;
wire PE_inst0_PE_output_width_1_num_0_valid;
wire [31:0] PE_inst0_read_config_data;
wire [0:0] PE_output_width_17_num_0_loopback_valid_out;
wire [0:0] PE_output_width_17_num_1_loopback_valid_out;
wire [0:0] PE_output_width_17_num_2_loopback_valid_out;
wire [0:0] PE_output_width_1_num_0_loopback_valid_out;
wire PondCore_inst0_PondTop_input_width_17_num_0_ready;
wire PondCore_inst0_PondTop_input_width_17_num_1_ready;
wire [16:0] PondCore_inst0_PondTop_output_width_17_num_0;
wire PondCore_inst0_PondTop_output_width_17_num_0_valid;
wire [16:0] PondCore_inst0_PondTop_output_width_17_num_1;
wire PondCore_inst0_PondTop_output_width_17_num_1_valid;
wire [0:0] PondCore_inst0_PondTop_output_width_1_num_0;
wire PondCore_inst0_PondTop_output_width_1_num_0_valid;
wire [0:0] PondCore_inst0_PondTop_output_width_1_num_1;
wire PondCore_inst0_PondTop_output_width_1_num_1_valid;
wire [31:0] PondCore_inst0_read_config_data;
wire [31:0] PondCore_inst0_read_config_data_1;
wire [0:0] PondTop_output_width_17_num_0_loopback_valid_out;
wire [0:0] PondTop_output_width_17_num_1_loopback_valid_out;
wire [0:0] PondTop_output_width_1_num_0_loopback_valid_out;
wire [0:0] PondTop_output_width_1_num_1_loopback_valid_out;
wire [0:0] PowerDomainConfigReg_inst0_ps_en_out;
wire [31:0] PowerDomainConfigReg_inst0_read_config_data;
wire [31:0] PowerDomainOR_O;
wire SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_0_ready_out;
wire SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_1_ready_out;
wire SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_2_ready_out;
wire SB_ID0_5TRACKS_B17_PE_PondTop_output_width_17_num_0_ready_out;
wire SB_ID0_5TRACKS_B17_PE_PondTop_output_width_17_num_1_ready_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_OUT_B17_valid_out;
wire [31:0] SB_ID0_5TRACKS_B17_PE_read_config_data;
wire SB_ID0_5TRACKS_B1_PE_PE_output_width_1_num_0_ready_out;
wire SB_ID0_5TRACKS_B1_PE_PondTop_output_width_1_num_0_ready_out;
wire SB_ID0_5TRACKS_B1_PE_PondTop_output_width_1_num_1_ready_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1_valid_out;
wire [31:0] SB_ID0_5TRACKS_B1_PE_read_config_data;
wire SB_T0_EAST_SB_OUT_B17_ready_and_Z;
wire SB_T0_EAST_SB_OUT_B1_ready_and_Z;
wire SB_T0_NORTH_SB_OUT_B17_ready_and_Z;
wire SB_T0_NORTH_SB_OUT_B1_ready_and_Z;
wire SB_T0_SOUTH_SB_OUT_B17_ready_and_Z;
wire SB_T0_SOUTH_SB_OUT_B1_ready_and_Z;
wire SB_T0_WEST_SB_OUT_B17_ready_and_Z;
wire SB_T0_WEST_SB_OUT_B1_ready_and_Z;
wire SB_T1_EAST_SB_OUT_B17_ready_and_Z;
wire SB_T1_EAST_SB_OUT_B1_ready_and_Z;
wire SB_T1_NORTH_SB_OUT_B17_ready_and_Z;
wire SB_T1_NORTH_SB_OUT_B1_ready_and_Z;
wire SB_T1_SOUTH_SB_OUT_B17_ready_and_Z;
wire SB_T1_SOUTH_SB_OUT_B1_ready_and_Z;
wire SB_T1_WEST_SB_OUT_B17_ready_and_Z;
wire SB_T1_WEST_SB_OUT_B1_ready_and_Z;
wire SB_T2_EAST_SB_OUT_B17_ready_and_Z;
wire SB_T2_EAST_SB_OUT_B1_ready_and_Z;
wire SB_T2_NORTH_SB_OUT_B17_ready_and_Z;
wire SB_T2_NORTH_SB_OUT_B1_ready_and_Z;
wire SB_T2_SOUTH_SB_OUT_B17_ready_and_Z;
wire SB_T2_SOUTH_SB_OUT_B1_ready_and_Z;
wire SB_T2_WEST_SB_OUT_B17_ready_and_Z;
wire SB_T2_WEST_SB_OUT_B1_ready_and_Z;
wire SB_T3_EAST_SB_OUT_B17_ready_and_Z;
wire SB_T3_EAST_SB_OUT_B1_ready_and_Z;
wire SB_T3_NORTH_SB_OUT_B17_ready_and_Z;
wire SB_T3_NORTH_SB_OUT_B1_ready_and_Z;
wire SB_T3_SOUTH_SB_OUT_B17_ready_and_Z;
wire SB_T3_SOUTH_SB_OUT_B1_ready_and_Z;
wire SB_T3_WEST_SB_OUT_B17_ready_and_Z;
wire SB_T3_WEST_SB_OUT_B1_ready_and_Z;
wire SB_T4_EAST_SB_OUT_B17_ready_and_Z;
wire SB_T4_EAST_SB_OUT_B1_ready_and_Z;
wire SB_T4_NORTH_SB_OUT_B17_ready_and_Z;
wire SB_T4_NORTH_SB_OUT_B1_ready_and_Z;
wire SB_T4_SOUTH_SB_OUT_B17_ready_and_Z;
wire SB_T4_SOUTH_SB_OUT_B1_ready_and_Z;
wire SB_T4_WEST_SB_OUT_B17_ready_and_Z;
wire SB_T4_WEST_SB_OUT_B1_ready_and_Z;
wire and_inst0_out;
wire and_inst1_out;
wire bit_const_1_None_out;
wire [7:0] const_0_8_out;
wire [8:0] const_511_9_out;
wire coreir_eq_16_inst0_out;
wire coreir_wrapOutClock_inst0_out;
wire coreir_wrapOutClock_inst1_out;
wire [31:0] read_data_mux_O;
wire [31:0] self_config_config_addr_out;
wire [16:0] CB_PE_input_width_17_num_0_I [20:0];
assign CB_PE_input_width_17_num_0_I[20] = PondCore_inst0_PondTop_output_width_17_num_0;
assign CB_PE_input_width_17_num_0_I[19] = SB_T4_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[18] = SB_T4_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[17] = SB_T4_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[16] = SB_T4_NORTH_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[15] = SB_T3_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[14] = SB_T3_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[13] = SB_T3_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[12] = SB_T3_NORTH_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[11] = SB_T2_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[10] = SB_T2_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[9] = SB_T2_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[8] = SB_T2_NORTH_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[7] = SB_T1_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[6] = SB_T1_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[5] = SB_T1_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[4] = SB_T1_NORTH_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[3] = SB_T0_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[2] = SB_T0_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[1] = SB_T0_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_0_I[0] = SB_T0_NORTH_SB_IN_B17;
wire [20:0] CB_PE_input_width_17_num_0_valid_in;
assign CB_PE_input_width_17_num_0_valid_in = {PondCore_inst0_PondTop_output_width_17_num_0_valid,SB_T4_WEST_SB_IN_B17_valid,SB_T4_EAST_SB_IN_B17_valid,SB_T4_SOUTH_SB_IN_B17_valid,SB_T4_NORTH_SB_IN_B17_valid,SB_T3_WEST_SB_IN_B17_valid,SB_T3_EAST_SB_IN_B17_valid,SB_T3_SOUTH_SB_IN_B17_valid,SB_T3_NORTH_SB_IN_B17_valid,SB_T2_WEST_SB_IN_B17_valid,SB_T2_EAST_SB_IN_B17_valid,SB_T2_SOUTH_SB_IN_B17_valid,SB_T2_NORTH_SB_IN_B17_valid,SB_T1_WEST_SB_IN_B17_valid,SB_T1_EAST_SB_IN_B17_valid,SB_T1_SOUTH_SB_IN_B17_valid,SB_T1_NORTH_SB_IN_B17_valid,SB_T0_WEST_SB_IN_B17_valid,SB_T0_EAST_SB_IN_B17_valid,SB_T0_SOUTH_SB_IN_B17_valid,SB_T0_NORTH_SB_IN_B17_valid};
CB_PE_input_width_17_num_0 CB_PE_input_width_17_num_0 (
    .I(CB_PE_input_width_17_num_0_I),
    .O(CB_PE_input_width_17_num_0_O),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_3_out),
    .enable(CB_PE_input_width_17_num_0_enable),
    .out_sel(CB_PE_input_width_17_num_0_out_sel),
    .read_config_data(CB_PE_input_width_17_num_0_read_config_data),
    .ready_in(PE_inst0_PE_input_width_17_num_0_ready[0]),
    .ready_out(CB_PE_input_width_17_num_0_ready_out),
    .reset(reset),
    .valid_in(CB_PE_input_width_17_num_0_valid_in),
    .valid_out(CB_PE_input_width_17_num_0_valid_out)
);
wire [16:0] CB_PE_input_width_17_num_1_I [20:0];
assign CB_PE_input_width_17_num_1_I[20] = PondCore_inst0_PondTop_output_width_17_num_0;
assign CB_PE_input_width_17_num_1_I[19] = SB_T4_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[18] = SB_T4_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[17] = SB_T4_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[16] = SB_T4_NORTH_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[15] = SB_T3_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[14] = SB_T3_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[13] = SB_T3_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[12] = SB_T3_NORTH_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[11] = SB_T2_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[10] = SB_T2_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[9] = SB_T2_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[8] = SB_T2_NORTH_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[7] = SB_T1_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[6] = SB_T1_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[5] = SB_T1_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[4] = SB_T1_NORTH_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[3] = SB_T0_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[2] = SB_T0_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[1] = SB_T0_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_1_I[0] = SB_T0_NORTH_SB_IN_B17;
wire [20:0] CB_PE_input_width_17_num_1_valid_in;
assign CB_PE_input_width_17_num_1_valid_in = {PondCore_inst0_PondTop_output_width_17_num_0_valid,SB_T4_WEST_SB_IN_B17_valid,SB_T4_EAST_SB_IN_B17_valid,SB_T4_SOUTH_SB_IN_B17_valid,SB_T4_NORTH_SB_IN_B17_valid,SB_T3_WEST_SB_IN_B17_valid,SB_T3_EAST_SB_IN_B17_valid,SB_T3_SOUTH_SB_IN_B17_valid,SB_T3_NORTH_SB_IN_B17_valid,SB_T2_WEST_SB_IN_B17_valid,SB_T2_EAST_SB_IN_B17_valid,SB_T2_SOUTH_SB_IN_B17_valid,SB_T2_NORTH_SB_IN_B17_valid,SB_T1_WEST_SB_IN_B17_valid,SB_T1_EAST_SB_IN_B17_valid,SB_T1_SOUTH_SB_IN_B17_valid,SB_T1_NORTH_SB_IN_B17_valid,SB_T0_WEST_SB_IN_B17_valid,SB_T0_EAST_SB_IN_B17_valid,SB_T0_SOUTH_SB_IN_B17_valid,SB_T0_NORTH_SB_IN_B17_valid};
CB_PE_input_width_17_num_1 CB_PE_input_width_17_num_1 (
    .I(CB_PE_input_width_17_num_1_I),
    .O(CB_PE_input_width_17_num_1_O),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_4_out),
    .enable(CB_PE_input_width_17_num_1_enable),
    .out_sel(CB_PE_input_width_17_num_1_out_sel),
    .read_config_data(CB_PE_input_width_17_num_1_read_config_data),
    .ready_in(PE_inst0_PE_input_width_17_num_1_ready[0]),
    .ready_out(CB_PE_input_width_17_num_1_ready_out),
    .reset(reset),
    .valid_in(CB_PE_input_width_17_num_1_valid_in),
    .valid_out(CB_PE_input_width_17_num_1_valid_out)
);
wire [16:0] CB_PE_input_width_17_num_2_I [20:0];
assign CB_PE_input_width_17_num_2_I[20] = PondCore_inst0_PondTop_output_width_17_num_0;
assign CB_PE_input_width_17_num_2_I[19] = SB_T4_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[18] = SB_T4_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[17] = SB_T4_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[16] = SB_T4_NORTH_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[15] = SB_T3_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[14] = SB_T3_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[13] = SB_T3_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[12] = SB_T3_NORTH_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[11] = SB_T2_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[10] = SB_T2_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[9] = SB_T2_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[8] = SB_T2_NORTH_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[7] = SB_T1_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[6] = SB_T1_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[5] = SB_T1_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[4] = SB_T1_NORTH_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[3] = SB_T0_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[2] = SB_T0_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[1] = SB_T0_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_2_I[0] = SB_T0_NORTH_SB_IN_B17;
wire [20:0] CB_PE_input_width_17_num_2_valid_in;
assign CB_PE_input_width_17_num_2_valid_in = {PondCore_inst0_PondTop_output_width_17_num_0_valid,SB_T4_WEST_SB_IN_B17_valid,SB_T4_EAST_SB_IN_B17_valid,SB_T4_SOUTH_SB_IN_B17_valid,SB_T4_NORTH_SB_IN_B17_valid,SB_T3_WEST_SB_IN_B17_valid,SB_T3_EAST_SB_IN_B17_valid,SB_T3_SOUTH_SB_IN_B17_valid,SB_T3_NORTH_SB_IN_B17_valid,SB_T2_WEST_SB_IN_B17_valid,SB_T2_EAST_SB_IN_B17_valid,SB_T2_SOUTH_SB_IN_B17_valid,SB_T2_NORTH_SB_IN_B17_valid,SB_T1_WEST_SB_IN_B17_valid,SB_T1_EAST_SB_IN_B17_valid,SB_T1_SOUTH_SB_IN_B17_valid,SB_T1_NORTH_SB_IN_B17_valid,SB_T0_WEST_SB_IN_B17_valid,SB_T0_EAST_SB_IN_B17_valid,SB_T0_SOUTH_SB_IN_B17_valid,SB_T0_NORTH_SB_IN_B17_valid};
CB_PE_input_width_17_num_2 CB_PE_input_width_17_num_2 (
    .I(CB_PE_input_width_17_num_2_I),
    .O(CB_PE_input_width_17_num_2_O),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_5_out),
    .enable(CB_PE_input_width_17_num_2_enable),
    .out_sel(CB_PE_input_width_17_num_2_out_sel),
    .read_config_data(CB_PE_input_width_17_num_2_read_config_data),
    .ready_in(PE_inst0_PE_input_width_17_num_2_ready[0]),
    .ready_out(CB_PE_input_width_17_num_2_ready_out),
    .reset(reset),
    .valid_in(CB_PE_input_width_17_num_2_valid_in),
    .valid_out(CB_PE_input_width_17_num_2_valid_out)
);
wire [16:0] CB_PE_input_width_17_num_3_I [19:0];
assign CB_PE_input_width_17_num_3_I[19] = SB_T4_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[18] = SB_T4_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[17] = SB_T4_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[16] = SB_T4_NORTH_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[15] = SB_T3_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[14] = SB_T3_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[13] = SB_T3_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[12] = SB_T3_NORTH_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[11] = SB_T2_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[10] = SB_T2_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[9] = SB_T2_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[8] = SB_T2_NORTH_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[7] = SB_T1_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[6] = SB_T1_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[5] = SB_T1_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[4] = SB_T1_NORTH_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[3] = SB_T0_WEST_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[2] = SB_T0_EAST_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[1] = SB_T0_SOUTH_SB_IN_B17;
assign CB_PE_input_width_17_num_3_I[0] = SB_T0_NORTH_SB_IN_B17;
wire [19:0] CB_PE_input_width_17_num_3_valid_in;
assign CB_PE_input_width_17_num_3_valid_in = {SB_T4_WEST_SB_IN_B17_valid,SB_T4_EAST_SB_IN_B17_valid,SB_T4_SOUTH_SB_IN_B17_valid,SB_T4_NORTH_SB_IN_B17_valid,SB_T3_WEST_SB_IN_B17_valid,SB_T3_EAST_SB_IN_B17_valid,SB_T3_SOUTH_SB_IN_B17_valid,SB_T3_NORTH_SB_IN_B17_valid,SB_T2_WEST_SB_IN_B17_valid,SB_T2_EAST_SB_IN_B17_valid,SB_T2_SOUTH_SB_IN_B17_valid,SB_T2_NORTH_SB_IN_B17_valid,SB_T1_WEST_SB_IN_B17_valid,SB_T1_EAST_SB_IN_B17_valid,SB_T1_SOUTH_SB_IN_B17_valid,SB_T1_NORTH_SB_IN_B17_valid,SB_T0_WEST_SB_IN_B17_valid,SB_T0_EAST_SB_IN_B17_valid,SB_T0_SOUTH_SB_IN_B17_valid,SB_T0_NORTH_SB_IN_B17_valid};
CB_PE_input_width_17_num_3 CB_PE_input_width_17_num_3 (
    .I(CB_PE_input_width_17_num_3_I),
    .O(CB_PE_input_width_17_num_3_O),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_6_out),
    .enable(CB_PE_input_width_17_num_3_enable),
    .out_sel(CB_PE_input_width_17_num_3_out_sel),
    .read_config_data(CB_PE_input_width_17_num_3_read_config_data),
    .ready_in(PE_inst0_PE_input_width_17_num_3_ready[0]),
    .ready_out(CB_PE_input_width_17_num_3_ready_out),
    .reset(reset),
    .valid_in(CB_PE_input_width_17_num_3_valid_in),
    .valid_out(CB_PE_input_width_17_num_3_valid_out)
);
wire [0:0] CB_PE_input_width_1_num_0_I [20:0];
assign CB_PE_input_width_1_num_0_I[20] = PondCore_inst0_PondTop_output_width_1_num_0;
assign CB_PE_input_width_1_num_0_I[19] = SB_T4_WEST_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[18] = SB_T4_EAST_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[17] = SB_T4_SOUTH_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[16] = SB_T4_NORTH_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[15] = SB_T3_WEST_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[14] = SB_T3_EAST_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[13] = SB_T3_SOUTH_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[12] = SB_T3_NORTH_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[11] = SB_T2_WEST_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[10] = SB_T2_EAST_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[9] = SB_T2_SOUTH_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[8] = SB_T2_NORTH_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[7] = SB_T1_WEST_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[6] = SB_T1_EAST_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[5] = SB_T1_SOUTH_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[4] = SB_T1_NORTH_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[3] = SB_T0_WEST_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[2] = SB_T0_EAST_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[1] = SB_T0_SOUTH_SB_IN_B1;
assign CB_PE_input_width_1_num_0_I[0] = SB_T0_NORTH_SB_IN_B1;
wire [20:0] CB_PE_input_width_1_num_0_valid_in;
assign CB_PE_input_width_1_num_0_valid_in = {PondCore_inst0_PondTop_output_width_1_num_0_valid,SB_T4_WEST_SB_IN_B1_valid,SB_T4_EAST_SB_IN_B1_valid,SB_T4_SOUTH_SB_IN_B1_valid,SB_T4_NORTH_SB_IN_B1_valid,SB_T3_WEST_SB_IN_B1_valid,SB_T3_EAST_SB_IN_B1_valid,SB_T3_SOUTH_SB_IN_B1_valid,SB_T3_NORTH_SB_IN_B1_valid,SB_T2_WEST_SB_IN_B1_valid,SB_T2_EAST_SB_IN_B1_valid,SB_T2_SOUTH_SB_IN_B1_valid,SB_T2_NORTH_SB_IN_B1_valid,SB_T1_WEST_SB_IN_B1_valid,SB_T1_EAST_SB_IN_B1_valid,SB_T1_SOUTH_SB_IN_B1_valid,SB_T1_NORTH_SB_IN_B1_valid,SB_T0_WEST_SB_IN_B1_valid,SB_T0_EAST_SB_IN_B1_valid,SB_T0_SOUTH_SB_IN_B1_valid,SB_T0_NORTH_SB_IN_B1_valid};
CB_PE_input_width_1_num_0 CB_PE_input_width_1_num_0 (
    .I(CB_PE_input_width_1_num_0_I),
    .O(CB_PE_input_width_1_num_0_O),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_7_out),
    .enable(CB_PE_input_width_1_num_0_enable),
    .out_sel(CB_PE_input_width_1_num_0_out_sel),
    .read_config_data(CB_PE_input_width_1_num_0_read_config_data),
    .ready_in(PE_inst0_PE_input_width_1_num_0_ready),
    .ready_out(CB_PE_input_width_1_num_0_ready_out),
    .reset(reset),
    .valid_in(CB_PE_input_width_1_num_0_valid_in),
    .valid_out(CB_PE_input_width_1_num_0_valid_out)
);
wire [0:0] CB_PE_input_width_1_num_1_I [19:0];
assign CB_PE_input_width_1_num_1_I[19] = SB_T4_WEST_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[18] = SB_T4_EAST_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[17] = SB_T4_SOUTH_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[16] = SB_T4_NORTH_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[15] = SB_T3_WEST_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[14] = SB_T3_EAST_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[13] = SB_T3_SOUTH_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[12] = SB_T3_NORTH_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[11] = SB_T2_WEST_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[10] = SB_T2_EAST_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[9] = SB_T2_SOUTH_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[8] = SB_T2_NORTH_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[7] = SB_T1_WEST_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[6] = SB_T1_EAST_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[5] = SB_T1_SOUTH_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[4] = SB_T1_NORTH_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[3] = SB_T0_WEST_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[2] = SB_T0_EAST_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[1] = SB_T0_SOUTH_SB_IN_B1;
assign CB_PE_input_width_1_num_1_I[0] = SB_T0_NORTH_SB_IN_B1;
wire [19:0] CB_PE_input_width_1_num_1_valid_in;
assign CB_PE_input_width_1_num_1_valid_in = {SB_T4_WEST_SB_IN_B1_valid,SB_T4_EAST_SB_IN_B1_valid,SB_T4_SOUTH_SB_IN_B1_valid,SB_T4_NORTH_SB_IN_B1_valid,SB_T3_WEST_SB_IN_B1_valid,SB_T3_EAST_SB_IN_B1_valid,SB_T3_SOUTH_SB_IN_B1_valid,SB_T3_NORTH_SB_IN_B1_valid,SB_T2_WEST_SB_IN_B1_valid,SB_T2_EAST_SB_IN_B1_valid,SB_T2_SOUTH_SB_IN_B1_valid,SB_T2_NORTH_SB_IN_B1_valid,SB_T1_WEST_SB_IN_B1_valid,SB_T1_EAST_SB_IN_B1_valid,SB_T1_SOUTH_SB_IN_B1_valid,SB_T1_NORTH_SB_IN_B1_valid,SB_T0_WEST_SB_IN_B1_valid,SB_T0_EAST_SB_IN_B1_valid,SB_T0_SOUTH_SB_IN_B1_valid,SB_T0_NORTH_SB_IN_B1_valid};
CB_PE_input_width_1_num_1 CB_PE_input_width_1_num_1 (
    .I(CB_PE_input_width_1_num_1_I),
    .O(CB_PE_input_width_1_num_1_O),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_8_out),
    .enable(CB_PE_input_width_1_num_1_enable),
    .out_sel(CB_PE_input_width_1_num_1_out_sel),
    .read_config_data(CB_PE_input_width_1_num_1_read_config_data),
    .ready_in(PE_inst0_PE_input_width_1_num_1_ready),
    .ready_out(CB_PE_input_width_1_num_1_ready_out),
    .reset(reset),
    .valid_in(CB_PE_input_width_1_num_1_valid_in),
    .valid_out(CB_PE_input_width_1_num_1_valid_out)
);
wire [0:0] CB_PE_input_width_1_num_2_I [19:0];
assign CB_PE_input_width_1_num_2_I[19] = SB_T4_WEST_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[18] = SB_T4_EAST_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[17] = SB_T4_SOUTH_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[16] = SB_T4_NORTH_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[15] = SB_T3_WEST_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[14] = SB_T3_EAST_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[13] = SB_T3_SOUTH_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[12] = SB_T3_NORTH_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[11] = SB_T2_WEST_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[10] = SB_T2_EAST_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[9] = SB_T2_SOUTH_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[8] = SB_T2_NORTH_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[7] = SB_T1_WEST_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[6] = SB_T1_EAST_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[5] = SB_T1_SOUTH_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[4] = SB_T1_NORTH_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[3] = SB_T0_WEST_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[2] = SB_T0_EAST_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[1] = SB_T0_SOUTH_SB_IN_B1;
assign CB_PE_input_width_1_num_2_I[0] = SB_T0_NORTH_SB_IN_B1;
wire [19:0] CB_PE_input_width_1_num_2_valid_in;
assign CB_PE_input_width_1_num_2_valid_in = {SB_T4_WEST_SB_IN_B1_valid,SB_T4_EAST_SB_IN_B1_valid,SB_T4_SOUTH_SB_IN_B1_valid,SB_T4_NORTH_SB_IN_B1_valid,SB_T3_WEST_SB_IN_B1_valid,SB_T3_EAST_SB_IN_B1_valid,SB_T3_SOUTH_SB_IN_B1_valid,SB_T3_NORTH_SB_IN_B1_valid,SB_T2_WEST_SB_IN_B1_valid,SB_T2_EAST_SB_IN_B1_valid,SB_T2_SOUTH_SB_IN_B1_valid,SB_T2_NORTH_SB_IN_B1_valid,SB_T1_WEST_SB_IN_B1_valid,SB_T1_EAST_SB_IN_B1_valid,SB_T1_SOUTH_SB_IN_B1_valid,SB_T1_NORTH_SB_IN_B1_valid,SB_T0_WEST_SB_IN_B1_valid,SB_T0_EAST_SB_IN_B1_valid,SB_T0_SOUTH_SB_IN_B1_valid,SB_T0_NORTH_SB_IN_B1_valid};
CB_PE_input_width_1_num_2 CB_PE_input_width_1_num_2 (
    .I(CB_PE_input_width_1_num_2_I),
    .O(CB_PE_input_width_1_num_2_O),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_9_out),
    .enable(CB_PE_input_width_1_num_2_enable),
    .out_sel(CB_PE_input_width_1_num_2_out_sel),
    .read_config_data(CB_PE_input_width_1_num_2_read_config_data),
    .ready_in(PE_inst0_PE_input_width_1_num_2_ready),
    .ready_out(CB_PE_input_width_1_num_2_ready_out),
    .reset(reset),
    .valid_in(CB_PE_input_width_1_num_2_valid_in),
    .valid_out(CB_PE_input_width_1_num_2_valid_out)
);
wire [16:0] CB_PondTop_input_width_17_num_0_I [20:0];
assign CB_PondTop_input_width_17_num_0_I[20] = PE_inst0_PE_output_width_17_num_0;
assign CB_PondTop_input_width_17_num_0_I[19] = SB_T4_WEST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[18] = SB_T4_EAST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[17] = SB_T4_SOUTH_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[16] = SB_T4_NORTH_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[15] = SB_T3_WEST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[14] = SB_T3_EAST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[13] = SB_T3_SOUTH_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[12] = SB_T3_NORTH_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[11] = SB_T2_WEST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[10] = SB_T2_EAST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[9] = SB_T2_SOUTH_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[8] = SB_T2_NORTH_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[7] = SB_T1_WEST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[6] = SB_T1_EAST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[5] = SB_T1_SOUTH_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[4] = SB_T1_NORTH_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[3] = SB_T0_WEST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[2] = SB_T0_EAST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[1] = SB_T0_SOUTH_SB_IN_B17;
assign CB_PondTop_input_width_17_num_0_I[0] = SB_T0_NORTH_SB_IN_B17;
wire [20:0] CB_PondTop_input_width_17_num_0_valid_in;
assign CB_PondTop_input_width_17_num_0_valid_in = {PE_inst0_PE_output_width_17_num_0_valid[0],SB_T4_WEST_SB_IN_B17_valid,SB_T4_EAST_SB_IN_B17_valid,SB_T4_SOUTH_SB_IN_B17_valid,SB_T4_NORTH_SB_IN_B17_valid,SB_T3_WEST_SB_IN_B17_valid,SB_T3_EAST_SB_IN_B17_valid,SB_T3_SOUTH_SB_IN_B17_valid,SB_T3_NORTH_SB_IN_B17_valid,SB_T2_WEST_SB_IN_B17_valid,SB_T2_EAST_SB_IN_B17_valid,SB_T2_SOUTH_SB_IN_B17_valid,SB_T2_NORTH_SB_IN_B17_valid,SB_T1_WEST_SB_IN_B17_valid,SB_T1_EAST_SB_IN_B17_valid,SB_T1_SOUTH_SB_IN_B17_valid,SB_T1_NORTH_SB_IN_B17_valid,SB_T0_WEST_SB_IN_B17_valid,SB_T0_EAST_SB_IN_B17_valid,SB_T0_SOUTH_SB_IN_B17_valid,SB_T0_NORTH_SB_IN_B17_valid};
CB_PondTop_input_width_17_num_0 CB_PondTop_input_width_17_num_0 (
    .I(CB_PondTop_input_width_17_num_0_I),
    .O(CB_PondTop_input_width_17_num_0_O),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_10_out),
    .enable(CB_PondTop_input_width_17_num_0_enable),
    .out_sel(CB_PondTop_input_width_17_num_0_out_sel),
    .read_config_data(CB_PondTop_input_width_17_num_0_read_config_data),
    .ready_in(PondCore_inst0_PondTop_input_width_17_num_0_ready),
    .ready_out(CB_PondTop_input_width_17_num_0_ready_out),
    .reset(reset),
    .valid_in(CB_PondTop_input_width_17_num_0_valid_in),
    .valid_out(CB_PondTop_input_width_17_num_0_valid_out)
);
wire [16:0] CB_PondTop_input_width_17_num_1_I [20:0];
assign CB_PondTop_input_width_17_num_1_I[20] = PE_inst0_PE_output_width_17_num_0;
assign CB_PondTop_input_width_17_num_1_I[19] = SB_T4_WEST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[18] = SB_T4_EAST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[17] = SB_T4_SOUTH_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[16] = SB_T4_NORTH_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[15] = SB_T3_WEST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[14] = SB_T3_EAST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[13] = SB_T3_SOUTH_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[12] = SB_T3_NORTH_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[11] = SB_T2_WEST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[10] = SB_T2_EAST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[9] = SB_T2_SOUTH_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[8] = SB_T2_NORTH_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[7] = SB_T1_WEST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[6] = SB_T1_EAST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[5] = SB_T1_SOUTH_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[4] = SB_T1_NORTH_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[3] = SB_T0_WEST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[2] = SB_T0_EAST_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[1] = SB_T0_SOUTH_SB_IN_B17;
assign CB_PondTop_input_width_17_num_1_I[0] = SB_T0_NORTH_SB_IN_B17;
wire [20:0] CB_PondTop_input_width_17_num_1_valid_in;
assign CB_PondTop_input_width_17_num_1_valid_in = {PE_inst0_PE_output_width_17_num_0_valid[0],SB_T4_WEST_SB_IN_B17_valid,SB_T4_EAST_SB_IN_B17_valid,SB_T4_SOUTH_SB_IN_B17_valid,SB_T4_NORTH_SB_IN_B17_valid,SB_T3_WEST_SB_IN_B17_valid,SB_T3_EAST_SB_IN_B17_valid,SB_T3_SOUTH_SB_IN_B17_valid,SB_T3_NORTH_SB_IN_B17_valid,SB_T2_WEST_SB_IN_B17_valid,SB_T2_EAST_SB_IN_B17_valid,SB_T2_SOUTH_SB_IN_B17_valid,SB_T2_NORTH_SB_IN_B17_valid,SB_T1_WEST_SB_IN_B17_valid,SB_T1_EAST_SB_IN_B17_valid,SB_T1_SOUTH_SB_IN_B17_valid,SB_T1_NORTH_SB_IN_B17_valid,SB_T0_WEST_SB_IN_B17_valid,SB_T0_EAST_SB_IN_B17_valid,SB_T0_SOUTH_SB_IN_B17_valid,SB_T0_NORTH_SB_IN_B17_valid};
CB_PondTop_input_width_17_num_1 CB_PondTop_input_width_17_num_1 (
    .I(CB_PondTop_input_width_17_num_1_I),
    .O(CB_PondTop_input_width_17_num_1_O),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_11_out),
    .enable(CB_PondTop_input_width_17_num_1_enable),
    .out_sel(CB_PondTop_input_width_17_num_1_out_sel),
    .read_config_data(CB_PondTop_input_width_17_num_1_read_config_data),
    .ready_in(PondCore_inst0_PondTop_input_width_17_num_1_ready),
    .ready_out(CB_PondTop_input_width_17_num_1_ready_out),
    .reset(reset),
    .valid_in(CB_PondTop_input_width_17_num_1_valid_in),
    .valid_out(CB_PondTop_input_width_17_num_1_valid_out)
);
wire [0:0] CB_flush_I [19:0];
assign CB_flush_I[19] = SB_T4_WEST_SB_IN_B1;
assign CB_flush_I[18] = SB_T4_EAST_SB_IN_B1;
assign CB_flush_I[17] = SB_T4_SOUTH_SB_IN_B1;
assign CB_flush_I[16] = SB_T4_NORTH_SB_IN_B1;
assign CB_flush_I[15] = SB_T3_WEST_SB_IN_B1;
assign CB_flush_I[14] = SB_T3_EAST_SB_IN_B1;
assign CB_flush_I[13] = SB_T3_SOUTH_SB_IN_B1;
assign CB_flush_I[12] = SB_T3_NORTH_SB_IN_B1;
assign CB_flush_I[11] = SB_T2_WEST_SB_IN_B1;
assign CB_flush_I[10] = SB_T2_EAST_SB_IN_B1;
assign CB_flush_I[9] = SB_T2_SOUTH_SB_IN_B1;
assign CB_flush_I[8] = SB_T2_NORTH_SB_IN_B1;
assign CB_flush_I[7] = SB_T1_WEST_SB_IN_B1;
assign CB_flush_I[6] = SB_T1_EAST_SB_IN_B1;
assign CB_flush_I[5] = SB_T1_SOUTH_SB_IN_B1;
assign CB_flush_I[4] = SB_T1_NORTH_SB_IN_B1;
assign CB_flush_I[3] = SB_T0_WEST_SB_IN_B1;
assign CB_flush_I[2] = SB_T0_EAST_SB_IN_B1;
assign CB_flush_I[1] = SB_T0_SOUTH_SB_IN_B1;
assign CB_flush_I[0] = SB_T0_NORTH_SB_IN_B1;
wire [19:0] CB_flush_valid_in;
assign CB_flush_valid_in = {SB_T4_WEST_SB_IN_B1_valid,SB_T4_EAST_SB_IN_B1_valid,SB_T4_SOUTH_SB_IN_B1_valid,SB_T4_NORTH_SB_IN_B1_valid,SB_T3_WEST_SB_IN_B1_valid,SB_T3_EAST_SB_IN_B1_valid,SB_T3_SOUTH_SB_IN_B1_valid,SB_T3_NORTH_SB_IN_B1_valid,SB_T2_WEST_SB_IN_B1_valid,SB_T2_EAST_SB_IN_B1_valid,SB_T2_SOUTH_SB_IN_B1_valid,SB_T2_NORTH_SB_IN_B1_valid,SB_T1_WEST_SB_IN_B1_valid,SB_T1_EAST_SB_IN_B1_valid,SB_T1_SOUTH_SB_IN_B1_valid,SB_T1_NORTH_SB_IN_B1_valid,SB_T0_WEST_SB_IN_B1_valid,SB_T0_EAST_SB_IN_B1_valid,SB_T0_SOUTH_SB_IN_B1_valid,SB_T0_NORTH_SB_IN_B1_valid};
CB_flush CB_flush (
    .I(CB_flush_I),
    .O(CB_flush_O),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_12_out),
    .enable(CB_flush_enable),
    .out_sel(CB_flush_out_sel),
    .read_config_data(CB_flush_read_config_data),
    .ready_in(bit_const_1_None_out),
    .ready_out(CB_flush_ready_out),
    .reset(reset),
    .valid_in(CB_flush_valid_in),
    .valid_out(CB_flush_valid_out)
);
Decode08 DECODE_FEATURE_0 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_0_O)
);
Decode18 DECODE_FEATURE_1 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_1_O)
);
Decode108 DECODE_FEATURE_10 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_10_O)
);
Decode118 DECODE_FEATURE_11 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_11_O)
);
Decode128 DECODE_FEATURE_12 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_12_O)
);
Decode138 DECODE_FEATURE_13 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_13_O)
);
Decode148 DECODE_FEATURE_14 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_14_O)
);
Decode158 DECODE_FEATURE_15 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_15_O)
);
Decode28 DECODE_FEATURE_2 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_2_O)
);
Decode38 DECODE_FEATURE_3 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_3_O)
);
Decode48 DECODE_FEATURE_4 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_4_O)
);
Decode58 DECODE_FEATURE_5 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_5_O)
);
Decode68 DECODE_FEATURE_6 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_6_O)
);
Decode78 DECODE_FEATURE_7 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_7_O)
);
Decode88 DECODE_FEATURE_8 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_8_O)
);
Decode98 DECODE_FEATURE_9 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_9_O)
);
corebit_and FEATURE_AND_0 (
    .in0(DECODE_FEATURE_0_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_0_out)
);
corebit_and FEATURE_AND_1 (
    .in0(DECODE_FEATURE_1_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_1_out)
);
corebit_and FEATURE_AND_10 (
    .in0(DECODE_FEATURE_10_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_10_out)
);
corebit_and FEATURE_AND_11 (
    .in0(DECODE_FEATURE_11_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_11_out)
);
corebit_and FEATURE_AND_12 (
    .in0(DECODE_FEATURE_12_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_12_out)
);
corebit_and FEATURE_AND_13 (
    .in0(DECODE_FEATURE_13_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_13_out)
);
corebit_and FEATURE_AND_14 (
    .in0(DECODE_FEATURE_14_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_14_out)
);
corebit_and FEATURE_AND_15 (
    .in0(DECODE_FEATURE_15_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_15_out)
);
corebit_and FEATURE_AND_2 (
    .in0(DECODE_FEATURE_2_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_2_out)
);
corebit_and FEATURE_AND_3 (
    .in0(DECODE_FEATURE_3_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_3_out)
);
corebit_and FEATURE_AND_4 (
    .in0(DECODE_FEATURE_4_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_4_out)
);
corebit_and FEATURE_AND_5 (
    .in0(DECODE_FEATURE_5_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_5_out)
);
corebit_and FEATURE_AND_6 (
    .in0(DECODE_FEATURE_6_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_6_out)
);
corebit_and FEATURE_AND_7 (
    .in0(DECODE_FEATURE_7_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_7_out)
);
corebit_and FEATURE_AND_8 (
    .in0(DECODE_FEATURE_8_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_8_out)
);
corebit_and FEATURE_AND_9 (
    .in0(DECODE_FEATURE_9_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_9_out)
);
PE PE_inst0 (
    .PE_input_width_17_num_0(CB_PE_input_width_17_num_0_O),
    .PE_input_width_17_num_0_ready(PE_inst0_PE_input_width_17_num_0_ready),
    .PE_input_width_17_num_0_valid(CB_PE_input_width_17_num_0_valid_out),
    .PE_input_width_17_num_1(CB_PE_input_width_17_num_1_O),
    .PE_input_width_17_num_1_ready(PE_inst0_PE_input_width_17_num_1_ready),
    .PE_input_width_17_num_1_valid(CB_PE_input_width_17_num_1_valid_out),
    .PE_input_width_17_num_2(CB_PE_input_width_17_num_2_O),
    .PE_input_width_17_num_2_ready(PE_inst0_PE_input_width_17_num_2_ready),
    .PE_input_width_17_num_2_valid(CB_PE_input_width_17_num_2_valid_out),
    .PE_input_width_17_num_3(CB_PE_input_width_17_num_3_O),
    .PE_input_width_17_num_3_ready(PE_inst0_PE_input_width_17_num_3_ready),
    .PE_input_width_17_num_3_valid(CB_PE_input_width_17_num_3_valid_out),
    .PE_input_width_1_num_0(CB_PE_input_width_1_num_0_O),
    .PE_input_width_1_num_0_ready(PE_inst0_PE_input_width_1_num_0_ready),
    .PE_input_width_1_num_0_valid(CB_PE_input_width_1_num_0_valid_out),
    .PE_input_width_1_num_1(CB_PE_input_width_1_num_1_O),
    .PE_input_width_1_num_1_ready(PE_inst0_PE_input_width_1_num_1_ready),
    .PE_input_width_1_num_1_valid(CB_PE_input_width_1_num_1_valid_out),
    .PE_input_width_1_num_2(CB_PE_input_width_1_num_2_O),
    .PE_input_width_1_num_2_ready(PE_inst0_PE_input_width_1_num_2_ready),
    .PE_input_width_1_num_2_valid(CB_PE_input_width_1_num_2_valid_out),
    .PE_output_width_17_num_0(PE_inst0_PE_output_width_17_num_0),
    .PE_output_width_17_num_0_ready(SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_0_ready_out),
    .PE_output_width_17_num_0_valid(PE_inst0_PE_output_width_17_num_0_valid),
    .PE_output_width_17_num_1(PE_inst0_PE_output_width_17_num_1),
    .PE_output_width_17_num_1_ready(SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_1_ready_out),
    .PE_output_width_17_num_1_valid(PE_inst0_PE_output_width_17_num_1_valid),
    .PE_output_width_17_num_2(PE_inst0_PE_output_width_17_num_2),
    .PE_output_width_17_num_2_ready(SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_2_ready_out),
    .PE_output_width_17_num_2_valid(PE_inst0_PE_output_width_17_num_2_valid),
    .PE_output_width_1_num_0(PE_inst0_PE_output_width_1_num_0),
    .PE_output_width_1_num_0_ready(SB_ID0_5TRACKS_B1_PE_PE_output_width_1_num_0_ready_out),
    .PE_output_width_1_num_0_valid(PE_inst0_PE_output_width_1_num_0_valid),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_0_out),
    .flush(CB_flush_O),
    .flush_core(flush),
    .read_config_data(PE_inst0_read_config_data),
    .reset(reset),
    .stall(stall)
);
ReadyValidLoopBack PE_output_width_17_num_0_loopback (
    .ready_in(SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_0_ready_out),
    .valid_in(PE_inst0_PE_output_width_17_num_0_valid),
    .valid_out(PE_output_width_17_num_0_loopback_valid_out)
);
ReadyValidLoopBack PE_output_width_17_num_1_loopback (
    .ready_in(SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_1_ready_out),
    .valid_in(PE_inst0_PE_output_width_17_num_1_valid),
    .valid_out(PE_output_width_17_num_1_loopback_valid_out)
);
ReadyValidLoopBack PE_output_width_17_num_2_loopback (
    .ready_in(SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_2_ready_out),
    .valid_in(PE_inst0_PE_output_width_17_num_2_valid),
    .valid_out(PE_output_width_17_num_2_loopback_valid_out)
);
ReadyValidLoopBack PE_output_width_1_num_0_loopback (
    .ready_in(SB_ID0_5TRACKS_B1_PE_PE_output_width_1_num_0_ready_out),
    .valid_in(PE_inst0_PE_output_width_1_num_0_valid),
    .valid_out(PE_output_width_1_num_0_loopback_valid_out)
);
PondCore PondCore_inst0 (
    .PondTop_input_width_17_num_0(CB_PondTop_input_width_17_num_0_O),
    .PondTop_input_width_17_num_0_ready(PondCore_inst0_PondTop_input_width_17_num_0_ready),
    .PondTop_input_width_17_num_0_valid(CB_PondTop_input_width_17_num_0_valid_out),
    .PondTop_input_width_17_num_1(CB_PondTop_input_width_17_num_1_O),
    .PondTop_input_width_17_num_1_ready(PondCore_inst0_PondTop_input_width_17_num_1_ready),
    .PondTop_input_width_17_num_1_valid(CB_PondTop_input_width_17_num_1_valid_out),
    .PondTop_output_width_17_num_0(PondCore_inst0_PondTop_output_width_17_num_0),
    .PondTop_output_width_17_num_0_ready(SB_ID0_5TRACKS_B17_PE_PondTop_output_width_17_num_0_ready_out),
    .PondTop_output_width_17_num_0_valid(PondCore_inst0_PondTop_output_width_17_num_0_valid),
    .PondTop_output_width_17_num_1(PondCore_inst0_PondTop_output_width_17_num_1),
    .PondTop_output_width_17_num_1_ready(SB_ID0_5TRACKS_B17_PE_PondTop_output_width_17_num_1_ready_out),
    .PondTop_output_width_17_num_1_valid(PondCore_inst0_PondTop_output_width_17_num_1_valid),
    .PondTop_output_width_1_num_0(PondCore_inst0_PondTop_output_width_1_num_0),
    .PondTop_output_width_1_num_0_ready(SB_ID0_5TRACKS_B1_PE_PondTop_output_width_1_num_0_ready_out),
    .PondTop_output_width_1_num_0_valid(PondCore_inst0_PondTop_output_width_1_num_0_valid),
    .PondTop_output_width_1_num_1(PondCore_inst0_PondTop_output_width_1_num_1),
    .PondTop_output_width_1_num_1_ready(SB_ID0_5TRACKS_B1_PE_PondTop_output_width_1_num_1_ready_out),
    .PondTop_output_width_1_num_1_valid(PondCore_inst0_PondTop_output_width_1_num_1_valid),
    .clk(clk),
    .config_1_config_addr(self_config_config_addr_out[31:24]),
    .config_1_config_data(config_config_data),
    .config_1_read(config_read),
    .config_1_write(FEATURE_AND_2_out),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_en_0(DECODE_FEATURE_2_O),
    .config_read(config_read),
    .config_write(FEATURE_AND_1_out),
    .flush(CB_flush_O),
    .flush_core(flush),
    .read_config_data(PondCore_inst0_read_config_data),
    .read_config_data_1(PondCore_inst0_read_config_data_1),
    .reset(reset),
    .stall(stall)
);
ReadyValidLoopBack PondTop_output_width_17_num_0_loopback (
    .ready_in(SB_ID0_5TRACKS_B17_PE_PondTop_output_width_17_num_0_ready_out),
    .valid_in(PondCore_inst0_PondTop_output_width_17_num_0_valid),
    .valid_out(PondTop_output_width_17_num_0_loopback_valid_out)
);
ReadyValidLoopBack PondTop_output_width_17_num_1_loopback (
    .ready_in(SB_ID0_5TRACKS_B17_PE_PondTop_output_width_17_num_1_ready_out),
    .valid_in(PondCore_inst0_PondTop_output_width_17_num_1_valid),
    .valid_out(PondTop_output_width_17_num_1_loopback_valid_out)
);
ReadyValidLoopBack PondTop_output_width_1_num_0_loopback (
    .ready_in(SB_ID0_5TRACKS_B1_PE_PondTop_output_width_1_num_0_ready_out),
    .valid_in(PondCore_inst0_PondTop_output_width_1_num_0_valid),
    .valid_out(PondTop_output_width_1_num_0_loopback_valid_out)
);
ReadyValidLoopBack PondTop_output_width_1_num_1_loopback (
    .ready_in(SB_ID0_5TRACKS_B1_PE_PondTop_output_width_1_num_1_ready_out),
    .valid_in(PondCore_inst0_PondTop_output_width_1_num_1_valid),
    .valid_out(PondTop_output_width_1_num_1_loopback_valid_out)
);
PowerDomainConfigReg PowerDomainConfigReg_inst0 (
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_15_out),
    .ps_en_out(PowerDomainConfigReg_inst0_ps_en_out),
    .read_config_data(PowerDomainConfigReg_inst0_read_config_data),
    .reset(reset)
);
PowerDomainOR PowerDomainOR (
    .I0(read_data_mux_O),
    .I1(read_config_data_in),
    .O(PowerDomainOR_O),
    .I_not(PowerDomainConfigReg_inst0_ps_en_out)
);
SB_ID0_5TRACKS_B17_PE SB_ID0_5TRACKS_B17_PE (
    .PE_input_width_17_num_0_enable(CB_PE_input_width_17_num_0_enable),
    .PE_input_width_17_num_0_out_sel(CB_PE_input_width_17_num_0_out_sel),
    .PE_input_width_17_num_0_ready(CB_PE_input_width_17_num_0_ready_out),
    .PE_input_width_17_num_1_enable(CB_PE_input_width_17_num_1_enable),
    .PE_input_width_17_num_1_out_sel(CB_PE_input_width_17_num_1_out_sel),
    .PE_input_width_17_num_1_ready(CB_PE_input_width_17_num_1_ready_out),
    .PE_input_width_17_num_2_enable(CB_PE_input_width_17_num_2_enable),
    .PE_input_width_17_num_2_out_sel(CB_PE_input_width_17_num_2_out_sel),
    .PE_input_width_17_num_2_ready(CB_PE_input_width_17_num_2_ready_out),
    .PE_input_width_17_num_3_enable(CB_PE_input_width_17_num_3_enable),
    .PE_input_width_17_num_3_out_sel(CB_PE_input_width_17_num_3_out_sel),
    .PE_input_width_17_num_3_ready(CB_PE_input_width_17_num_3_ready_out),
    .PE_output_width_17_num_0(PE_inst0_PE_output_width_17_num_0),
    .PE_output_width_17_num_0_ready_out(SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_0_ready_out),
    .PE_output_width_17_num_0_valid(PE_output_width_17_num_0_loopback_valid_out[0]),
    .PE_output_width_17_num_1(PE_inst0_PE_output_width_17_num_1),
    .PE_output_width_17_num_1_ready_out(SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_1_ready_out),
    .PE_output_width_17_num_1_valid(PE_output_width_17_num_1_loopback_valid_out[0]),
    .PE_output_width_17_num_2(PE_inst0_PE_output_width_17_num_2),
    .PE_output_width_17_num_2_ready_out(SB_ID0_5TRACKS_B17_PE_PE_output_width_17_num_2_ready_out),
    .PE_output_width_17_num_2_valid(PE_output_width_17_num_2_loopback_valid_out[0]),
    .PondTop_input_width_17_num_0_enable(CB_PondTop_input_width_17_num_0_enable),
    .PondTop_input_width_17_num_0_out_sel(CB_PondTop_input_width_17_num_0_out_sel),
    .PondTop_input_width_17_num_0_ready(CB_PondTop_input_width_17_num_0_ready_out),
    .PondTop_input_width_17_num_1_enable(CB_PondTop_input_width_17_num_1_enable),
    .PondTop_input_width_17_num_1_out_sel(CB_PondTop_input_width_17_num_1_out_sel),
    .PondTop_input_width_17_num_1_ready(CB_PondTop_input_width_17_num_1_ready_out),
    .PondTop_output_width_17_num_0_ready_out(SB_ID0_5TRACKS_B17_PE_PondTop_output_width_17_num_0_ready_out),
    .PondTop_output_width_17_num_0_valid(PondTop_output_width_17_num_0_loopback_valid_out[0]),
    .PondTop_output_width_17_num_1(PondCore_inst0_PondTop_output_width_17_num_1),
    .PondTop_output_width_17_num_1_ready_out(SB_ID0_5TRACKS_B17_PE_PondTop_output_width_17_num_1_ready_out),
    .PondTop_output_width_17_num_1_valid(PondTop_output_width_17_num_1_loopback_valid_out[0]),
    .SB_T0_EAST_SB_IN_B17(SB_T0_EAST_SB_IN_B17),
    .SB_T0_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_IN_B17_enable),
    .SB_T0_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_IN_B17_ready_out),
    .SB_T0_EAST_SB_IN_B17_valid_in(SB_T0_EAST_SB_IN_B17_valid),
    .SB_T0_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_OUT_B17_enable),
    .SB_T0_EAST_SB_OUT_B17_ready_in(SB_T0_EAST_SB_OUT_B17_ready_and_Z),
    .SB_T0_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_OUT_B17_valid_out),
    .SB_T0_NORTH_SB_IN_B17(SB_T0_NORTH_SB_IN_B17),
    .SB_T0_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_IN_B17_enable),
    .SB_T0_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_IN_B17_ready_out),
    .SB_T0_NORTH_SB_IN_B17_valid_in(SB_T0_NORTH_SB_IN_B17_valid),
    .SB_T0_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_OUT_B17_enable),
    .SB_T0_NORTH_SB_OUT_B17_ready_in(SB_T0_NORTH_SB_OUT_B17_ready_and_Z),
    .SB_T0_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_OUT_B17_valid_out),
    .SB_T0_SOUTH_SB_IN_B17(SB_T0_SOUTH_SB_IN_B17),
    .SB_T0_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_IN_B17_enable),
    .SB_T0_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_IN_B17_ready_out),
    .SB_T0_SOUTH_SB_IN_B17_valid_in(SB_T0_SOUTH_SB_IN_B17_valid),
    .SB_T0_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_OUT_B17_enable),
    .SB_T0_SOUTH_SB_OUT_B17_ready_in(SB_T0_SOUTH_SB_OUT_B17_ready_and_Z),
    .SB_T0_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_OUT_B17_valid_out),
    .SB_T0_WEST_SB_IN_B17(SB_T0_WEST_SB_IN_B17),
    .SB_T0_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_IN_B17_enable),
    .SB_T0_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_IN_B17_ready_out),
    .SB_T0_WEST_SB_IN_B17_valid_in(SB_T0_WEST_SB_IN_B17_valid),
    .SB_T0_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_OUT_B17_enable),
    .SB_T0_WEST_SB_OUT_B17_ready_in(SB_T0_WEST_SB_OUT_B17_ready_and_Z),
    .SB_T0_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_OUT_B17_valid_out),
    .SB_T1_EAST_SB_IN_B17(SB_T1_EAST_SB_IN_B17),
    .SB_T1_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_IN_B17_enable),
    .SB_T1_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_IN_B17_ready_out),
    .SB_T1_EAST_SB_IN_B17_valid_in(SB_T1_EAST_SB_IN_B17_valid),
    .SB_T1_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_OUT_B17_enable),
    .SB_T1_EAST_SB_OUT_B17_ready_in(SB_T1_EAST_SB_OUT_B17_ready_and_Z),
    .SB_T1_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_OUT_B17_valid_out),
    .SB_T1_NORTH_SB_IN_B17(SB_T1_NORTH_SB_IN_B17),
    .SB_T1_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_IN_B17_enable),
    .SB_T1_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_IN_B17_ready_out),
    .SB_T1_NORTH_SB_IN_B17_valid_in(SB_T1_NORTH_SB_IN_B17_valid),
    .SB_T1_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_OUT_B17_enable),
    .SB_T1_NORTH_SB_OUT_B17_ready_in(SB_T1_NORTH_SB_OUT_B17_ready_and_Z),
    .SB_T1_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_OUT_B17_valid_out),
    .SB_T1_SOUTH_SB_IN_B17(SB_T1_SOUTH_SB_IN_B17),
    .SB_T1_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_IN_B17_enable),
    .SB_T1_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_IN_B17_ready_out),
    .SB_T1_SOUTH_SB_IN_B17_valid_in(SB_T1_SOUTH_SB_IN_B17_valid),
    .SB_T1_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_OUT_B17_enable),
    .SB_T1_SOUTH_SB_OUT_B17_ready_in(SB_T1_SOUTH_SB_OUT_B17_ready_and_Z),
    .SB_T1_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_OUT_B17_valid_out),
    .SB_T1_WEST_SB_IN_B17(SB_T1_WEST_SB_IN_B17),
    .SB_T1_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_IN_B17_enable),
    .SB_T1_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_IN_B17_ready_out),
    .SB_T1_WEST_SB_IN_B17_valid_in(SB_T1_WEST_SB_IN_B17_valid),
    .SB_T1_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_OUT_B17_enable),
    .SB_T1_WEST_SB_OUT_B17_ready_in(SB_T1_WEST_SB_OUT_B17_ready_and_Z),
    .SB_T1_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_OUT_B17_valid_out),
    .SB_T2_EAST_SB_IN_B17(SB_T2_EAST_SB_IN_B17),
    .SB_T2_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_IN_B17_enable),
    .SB_T2_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_IN_B17_ready_out),
    .SB_T2_EAST_SB_IN_B17_valid_in(SB_T2_EAST_SB_IN_B17_valid),
    .SB_T2_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_OUT_B17_enable),
    .SB_T2_EAST_SB_OUT_B17_ready_in(SB_T2_EAST_SB_OUT_B17_ready_and_Z),
    .SB_T2_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_OUT_B17_valid_out),
    .SB_T2_NORTH_SB_IN_B17(SB_T2_NORTH_SB_IN_B17),
    .SB_T2_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_IN_B17_enable),
    .SB_T2_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_IN_B17_ready_out),
    .SB_T2_NORTH_SB_IN_B17_valid_in(SB_T2_NORTH_SB_IN_B17_valid),
    .SB_T2_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_OUT_B17_enable),
    .SB_T2_NORTH_SB_OUT_B17_ready_in(SB_T2_NORTH_SB_OUT_B17_ready_and_Z),
    .SB_T2_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_OUT_B17_valid_out),
    .SB_T2_SOUTH_SB_IN_B17(SB_T2_SOUTH_SB_IN_B17),
    .SB_T2_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_IN_B17_enable),
    .SB_T2_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_IN_B17_ready_out),
    .SB_T2_SOUTH_SB_IN_B17_valid_in(SB_T2_SOUTH_SB_IN_B17_valid),
    .SB_T2_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_OUT_B17_enable),
    .SB_T2_SOUTH_SB_OUT_B17_ready_in(SB_T2_SOUTH_SB_OUT_B17_ready_and_Z),
    .SB_T2_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_OUT_B17_valid_out),
    .SB_T2_WEST_SB_IN_B17(SB_T2_WEST_SB_IN_B17),
    .SB_T2_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_IN_B17_enable),
    .SB_T2_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_IN_B17_ready_out),
    .SB_T2_WEST_SB_IN_B17_valid_in(SB_T2_WEST_SB_IN_B17_valid),
    .SB_T2_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_OUT_B17_enable),
    .SB_T2_WEST_SB_OUT_B17_ready_in(SB_T2_WEST_SB_OUT_B17_ready_and_Z),
    .SB_T2_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_OUT_B17_valid_out),
    .SB_T3_EAST_SB_IN_B17(SB_T3_EAST_SB_IN_B17),
    .SB_T3_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_IN_B17_enable),
    .SB_T3_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_IN_B17_ready_out),
    .SB_T3_EAST_SB_IN_B17_valid_in(SB_T3_EAST_SB_IN_B17_valid),
    .SB_T3_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_OUT_B17_enable),
    .SB_T3_EAST_SB_OUT_B17_ready_in(SB_T3_EAST_SB_OUT_B17_ready_and_Z),
    .SB_T3_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_OUT_B17_valid_out),
    .SB_T3_NORTH_SB_IN_B17(SB_T3_NORTH_SB_IN_B17),
    .SB_T3_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_IN_B17_enable),
    .SB_T3_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_IN_B17_ready_out),
    .SB_T3_NORTH_SB_IN_B17_valid_in(SB_T3_NORTH_SB_IN_B17_valid),
    .SB_T3_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_OUT_B17_enable),
    .SB_T3_NORTH_SB_OUT_B17_ready_in(SB_T3_NORTH_SB_OUT_B17_ready_and_Z),
    .SB_T3_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_OUT_B17_valid_out),
    .SB_T3_SOUTH_SB_IN_B17(SB_T3_SOUTH_SB_IN_B17),
    .SB_T3_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_IN_B17_enable),
    .SB_T3_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_IN_B17_ready_out),
    .SB_T3_SOUTH_SB_IN_B17_valid_in(SB_T3_SOUTH_SB_IN_B17_valid),
    .SB_T3_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_OUT_B17_enable),
    .SB_T3_SOUTH_SB_OUT_B17_ready_in(SB_T3_SOUTH_SB_OUT_B17_ready_and_Z),
    .SB_T3_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_OUT_B17_valid_out),
    .SB_T3_WEST_SB_IN_B17(SB_T3_WEST_SB_IN_B17),
    .SB_T3_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_IN_B17_enable),
    .SB_T3_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_IN_B17_ready_out),
    .SB_T3_WEST_SB_IN_B17_valid_in(SB_T3_WEST_SB_IN_B17_valid),
    .SB_T3_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_OUT_B17_enable),
    .SB_T3_WEST_SB_OUT_B17_ready_in(SB_T3_WEST_SB_OUT_B17_ready_and_Z),
    .SB_T3_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_OUT_B17_valid_out),
    .SB_T4_EAST_SB_IN_B17(SB_T4_EAST_SB_IN_B17),
    .SB_T4_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_IN_B17_enable),
    .SB_T4_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_IN_B17_ready_out),
    .SB_T4_EAST_SB_IN_B17_valid_in(SB_T4_EAST_SB_IN_B17_valid),
    .SB_T4_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_OUT_B17_enable),
    .SB_T4_EAST_SB_OUT_B17_ready_in(SB_T4_EAST_SB_OUT_B17_ready_and_Z),
    .SB_T4_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_OUT_B17_valid_out),
    .SB_T4_NORTH_SB_IN_B17(SB_T4_NORTH_SB_IN_B17),
    .SB_T4_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_IN_B17_enable),
    .SB_T4_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_IN_B17_ready_out),
    .SB_T4_NORTH_SB_IN_B17_valid_in(SB_T4_NORTH_SB_IN_B17_valid),
    .SB_T4_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_OUT_B17_enable),
    .SB_T4_NORTH_SB_OUT_B17_ready_in(SB_T4_NORTH_SB_OUT_B17_ready_and_Z),
    .SB_T4_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_OUT_B17_valid_out),
    .SB_T4_SOUTH_SB_IN_B17(SB_T4_SOUTH_SB_IN_B17),
    .SB_T4_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_IN_B17_enable),
    .SB_T4_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_IN_B17_ready_out),
    .SB_T4_SOUTH_SB_IN_B17_valid_in(SB_T4_SOUTH_SB_IN_B17_valid),
    .SB_T4_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_OUT_B17_enable),
    .SB_T4_SOUTH_SB_OUT_B17_ready_in(SB_T4_SOUTH_SB_OUT_B17_ready_and_Z),
    .SB_T4_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_OUT_B17_valid_out),
    .SB_T4_WEST_SB_IN_B17(SB_T4_WEST_SB_IN_B17),
    .SB_T4_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_IN_B17_enable),
    .SB_T4_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_IN_B17_ready_out),
    .SB_T4_WEST_SB_IN_B17_valid_in(SB_T4_WEST_SB_IN_B17_valid),
    .SB_T4_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_OUT_B17_enable),
    .SB_T4_WEST_SB_OUT_B17_ready_in(SB_T4_WEST_SB_OUT_B17_ready_and_Z),
    .SB_T4_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_OUT_B17_valid_out),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_14_out),
    .read_config_data(SB_ID0_5TRACKS_B17_PE_read_config_data),
    .reset(reset),
    .stall(stall)
);
SB_ID0_5TRACKS_B1_PE SB_ID0_5TRACKS_B1_PE (
    .PE_input_width_1_num_0_enable(CB_PE_input_width_1_num_0_enable),
    .PE_input_width_1_num_0_out_sel(CB_PE_input_width_1_num_0_out_sel),
    .PE_input_width_1_num_0_ready(CB_PE_input_width_1_num_0_ready_out),
    .PE_input_width_1_num_1_enable(CB_PE_input_width_1_num_1_enable),
    .PE_input_width_1_num_1_out_sel(CB_PE_input_width_1_num_1_out_sel),
    .PE_input_width_1_num_1_ready(CB_PE_input_width_1_num_1_ready_out),
    .PE_input_width_1_num_2_enable(CB_PE_input_width_1_num_2_enable),
    .PE_input_width_1_num_2_out_sel(CB_PE_input_width_1_num_2_out_sel),
    .PE_input_width_1_num_2_ready(CB_PE_input_width_1_num_2_ready_out),
    .PE_output_width_1_num_0(PE_inst0_PE_output_width_1_num_0),
    .PE_output_width_1_num_0_ready_out(SB_ID0_5TRACKS_B1_PE_PE_output_width_1_num_0_ready_out),
    .PE_output_width_1_num_0_valid(PE_output_width_1_num_0_loopback_valid_out[0]),
    .PondTop_output_width_1_num_0(PondCore_inst0_PondTop_output_width_1_num_0),
    .PondTop_output_width_1_num_0_ready_out(SB_ID0_5TRACKS_B1_PE_PondTop_output_width_1_num_0_ready_out),
    .PondTop_output_width_1_num_0_valid(PondTop_output_width_1_num_0_loopback_valid_out[0]),
    .PondTop_output_width_1_num_1(PondCore_inst0_PondTop_output_width_1_num_1),
    .PondTop_output_width_1_num_1_ready_out(SB_ID0_5TRACKS_B1_PE_PondTop_output_width_1_num_1_ready_out),
    .PondTop_output_width_1_num_1_valid(PondTop_output_width_1_num_1_loopback_valid_out[0]),
    .SB_T0_EAST_SB_IN_B1(SB_T0_EAST_SB_IN_B1),
    .SB_T0_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_IN_B1_enable),
    .SB_T0_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_IN_B1_ready_out),
    .SB_T0_EAST_SB_IN_B1_valid_in(SB_T0_EAST_SB_IN_B1_valid),
    .SB_T0_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1_enable),
    .SB_T0_EAST_SB_OUT_B1_ready_in(SB_T0_EAST_SB_OUT_B1_ready_and_Z),
    .SB_T0_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1_valid_out),
    .SB_T0_NORTH_SB_IN_B1(SB_T0_NORTH_SB_IN_B1),
    .SB_T0_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_IN_B1_enable),
    .SB_T0_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_IN_B1_ready_out),
    .SB_T0_NORTH_SB_IN_B1_valid_in(SB_T0_NORTH_SB_IN_B1_valid),
    .SB_T0_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1_enable),
    .SB_T0_NORTH_SB_OUT_B1_ready_in(SB_T0_NORTH_SB_OUT_B1_ready_and_Z),
    .SB_T0_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1_valid_out),
    .SB_T0_SOUTH_SB_IN_B1(SB_T0_SOUTH_SB_IN_B1),
    .SB_T0_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_IN_B1_enable),
    .SB_T0_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_IN_B1_ready_out),
    .SB_T0_SOUTH_SB_IN_B1_valid_in(SB_T0_SOUTH_SB_IN_B1_valid),
    .SB_T0_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1_enable),
    .SB_T0_SOUTH_SB_OUT_B1_ready_in(SB_T0_SOUTH_SB_OUT_B1_ready_and_Z),
    .SB_T0_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1_valid_out),
    .SB_T0_WEST_SB_IN_B1(SB_T0_WEST_SB_IN_B1),
    .SB_T0_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_IN_B1_enable),
    .SB_T0_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_IN_B1_ready_out),
    .SB_T0_WEST_SB_IN_B1_valid_in(SB_T0_WEST_SB_IN_B1_valid),
    .SB_T0_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1_enable),
    .SB_T0_WEST_SB_OUT_B1_ready_in(SB_T0_WEST_SB_OUT_B1_ready_and_Z),
    .SB_T0_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1_valid_out),
    .SB_T1_EAST_SB_IN_B1(SB_T1_EAST_SB_IN_B1),
    .SB_T1_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_IN_B1_enable),
    .SB_T1_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_IN_B1_ready_out),
    .SB_T1_EAST_SB_IN_B1_valid_in(SB_T1_EAST_SB_IN_B1_valid),
    .SB_T1_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1_enable),
    .SB_T1_EAST_SB_OUT_B1_ready_in(SB_T1_EAST_SB_OUT_B1_ready_and_Z),
    .SB_T1_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1_valid_out),
    .SB_T1_NORTH_SB_IN_B1(SB_T1_NORTH_SB_IN_B1),
    .SB_T1_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_IN_B1_enable),
    .SB_T1_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_IN_B1_ready_out),
    .SB_T1_NORTH_SB_IN_B1_valid_in(SB_T1_NORTH_SB_IN_B1_valid),
    .SB_T1_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1_enable),
    .SB_T1_NORTH_SB_OUT_B1_ready_in(SB_T1_NORTH_SB_OUT_B1_ready_and_Z),
    .SB_T1_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1_valid_out),
    .SB_T1_SOUTH_SB_IN_B1(SB_T1_SOUTH_SB_IN_B1),
    .SB_T1_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_IN_B1_enable),
    .SB_T1_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_IN_B1_ready_out),
    .SB_T1_SOUTH_SB_IN_B1_valid_in(SB_T1_SOUTH_SB_IN_B1_valid),
    .SB_T1_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1_enable),
    .SB_T1_SOUTH_SB_OUT_B1_ready_in(SB_T1_SOUTH_SB_OUT_B1_ready_and_Z),
    .SB_T1_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1_valid_out),
    .SB_T1_WEST_SB_IN_B1(SB_T1_WEST_SB_IN_B1),
    .SB_T1_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_IN_B1_enable),
    .SB_T1_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_IN_B1_ready_out),
    .SB_T1_WEST_SB_IN_B1_valid_in(SB_T1_WEST_SB_IN_B1_valid),
    .SB_T1_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1_enable),
    .SB_T1_WEST_SB_OUT_B1_ready_in(SB_T1_WEST_SB_OUT_B1_ready_and_Z),
    .SB_T1_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1_valid_out),
    .SB_T2_EAST_SB_IN_B1(SB_T2_EAST_SB_IN_B1),
    .SB_T2_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_IN_B1_enable),
    .SB_T2_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_IN_B1_ready_out),
    .SB_T2_EAST_SB_IN_B1_valid_in(SB_T2_EAST_SB_IN_B1_valid),
    .SB_T2_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1_enable),
    .SB_T2_EAST_SB_OUT_B1_ready_in(SB_T2_EAST_SB_OUT_B1_ready_and_Z),
    .SB_T2_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1_valid_out),
    .SB_T2_NORTH_SB_IN_B1(SB_T2_NORTH_SB_IN_B1),
    .SB_T2_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_IN_B1_enable),
    .SB_T2_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_IN_B1_ready_out),
    .SB_T2_NORTH_SB_IN_B1_valid_in(SB_T2_NORTH_SB_IN_B1_valid),
    .SB_T2_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1_enable),
    .SB_T2_NORTH_SB_OUT_B1_ready_in(SB_T2_NORTH_SB_OUT_B1_ready_and_Z),
    .SB_T2_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1_valid_out),
    .SB_T2_SOUTH_SB_IN_B1(SB_T2_SOUTH_SB_IN_B1),
    .SB_T2_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_IN_B1_enable),
    .SB_T2_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_IN_B1_ready_out),
    .SB_T2_SOUTH_SB_IN_B1_valid_in(SB_T2_SOUTH_SB_IN_B1_valid),
    .SB_T2_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1_enable),
    .SB_T2_SOUTH_SB_OUT_B1_ready_in(SB_T2_SOUTH_SB_OUT_B1_ready_and_Z),
    .SB_T2_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1_valid_out),
    .SB_T2_WEST_SB_IN_B1(SB_T2_WEST_SB_IN_B1),
    .SB_T2_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_IN_B1_enable),
    .SB_T2_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_IN_B1_ready_out),
    .SB_T2_WEST_SB_IN_B1_valid_in(SB_T2_WEST_SB_IN_B1_valid),
    .SB_T2_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1_enable),
    .SB_T2_WEST_SB_OUT_B1_ready_in(SB_T2_WEST_SB_OUT_B1_ready_and_Z),
    .SB_T2_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1_valid_out),
    .SB_T3_EAST_SB_IN_B1(SB_T3_EAST_SB_IN_B1),
    .SB_T3_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_IN_B1_enable),
    .SB_T3_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_IN_B1_ready_out),
    .SB_T3_EAST_SB_IN_B1_valid_in(SB_T3_EAST_SB_IN_B1_valid),
    .SB_T3_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1_enable),
    .SB_T3_EAST_SB_OUT_B1_ready_in(SB_T3_EAST_SB_OUT_B1_ready_and_Z),
    .SB_T3_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1_valid_out),
    .SB_T3_NORTH_SB_IN_B1(SB_T3_NORTH_SB_IN_B1),
    .SB_T3_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_IN_B1_enable),
    .SB_T3_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_IN_B1_ready_out),
    .SB_T3_NORTH_SB_IN_B1_valid_in(SB_T3_NORTH_SB_IN_B1_valid),
    .SB_T3_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1_enable),
    .SB_T3_NORTH_SB_OUT_B1_ready_in(SB_T3_NORTH_SB_OUT_B1_ready_and_Z),
    .SB_T3_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1_valid_out),
    .SB_T3_SOUTH_SB_IN_B1(SB_T3_SOUTH_SB_IN_B1),
    .SB_T3_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_IN_B1_enable),
    .SB_T3_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_IN_B1_ready_out),
    .SB_T3_SOUTH_SB_IN_B1_valid_in(SB_T3_SOUTH_SB_IN_B1_valid),
    .SB_T3_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1_enable),
    .SB_T3_SOUTH_SB_OUT_B1_ready_in(SB_T3_SOUTH_SB_OUT_B1_ready_and_Z),
    .SB_T3_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1_valid_out),
    .SB_T3_WEST_SB_IN_B1(SB_T3_WEST_SB_IN_B1),
    .SB_T3_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_IN_B1_enable),
    .SB_T3_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_IN_B1_ready_out),
    .SB_T3_WEST_SB_IN_B1_valid_in(SB_T3_WEST_SB_IN_B1_valid),
    .SB_T3_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1_enable),
    .SB_T3_WEST_SB_OUT_B1_ready_in(SB_T3_WEST_SB_OUT_B1_ready_and_Z),
    .SB_T3_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1_valid_out),
    .SB_T4_EAST_SB_IN_B1(SB_T4_EAST_SB_IN_B1),
    .SB_T4_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_IN_B1_enable),
    .SB_T4_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_IN_B1_ready_out),
    .SB_T4_EAST_SB_IN_B1_valid_in(SB_T4_EAST_SB_IN_B1_valid),
    .SB_T4_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1_enable),
    .SB_T4_EAST_SB_OUT_B1_ready_in(SB_T4_EAST_SB_OUT_B1_ready_and_Z),
    .SB_T4_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1_valid_out),
    .SB_T4_NORTH_SB_IN_B1(SB_T4_NORTH_SB_IN_B1),
    .SB_T4_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_IN_B1_enable),
    .SB_T4_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_IN_B1_ready_out),
    .SB_T4_NORTH_SB_IN_B1_valid_in(SB_T4_NORTH_SB_IN_B1_valid),
    .SB_T4_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1_enable),
    .SB_T4_NORTH_SB_OUT_B1_ready_in(SB_T4_NORTH_SB_OUT_B1_ready_and_Z),
    .SB_T4_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1_valid_out),
    .SB_T4_SOUTH_SB_IN_B1(SB_T4_SOUTH_SB_IN_B1),
    .SB_T4_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_IN_B1_enable),
    .SB_T4_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_IN_B1_ready_out),
    .SB_T4_SOUTH_SB_IN_B1_valid_in(SB_T4_SOUTH_SB_IN_B1_valid),
    .SB_T4_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1_enable),
    .SB_T4_SOUTH_SB_OUT_B1_ready_in(SB_T4_SOUTH_SB_OUT_B1_ready_and_Z),
    .SB_T4_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1_valid_out),
    .SB_T4_WEST_SB_IN_B1(SB_T4_WEST_SB_IN_B1),
    .SB_T4_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_IN_B1_enable),
    .SB_T4_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_IN_B1_ready_out),
    .SB_T4_WEST_SB_IN_B1_valid_in(SB_T4_WEST_SB_IN_B1_valid),
    .SB_T4_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1_enable),
    .SB_T4_WEST_SB_OUT_B1_ready_in(SB_T4_WEST_SB_OUT_B1_ready_and_Z),
    .SB_T4_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1_valid_out),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_13_out),
    .read_config_data(SB_ID0_5TRACKS_B1_PE_read_config_data),
    .reset(reset),
    .stall(stall)
);
and_cell SB_T0_EAST_SB_OUT_B17_ready_and (
    .A(SB_T0_EAST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_OUT_B17_enable),
    .Z(SB_T0_EAST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T0_EAST_SB_OUT_B1_ready_and (
    .A(SB_T0_EAST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1_enable),
    .Z(SB_T0_EAST_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T0_NORTH_SB_OUT_B17_ready_and (
    .A(SB_T0_NORTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_OUT_B17_enable),
    .Z(SB_T0_NORTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T0_NORTH_SB_OUT_B1_ready_and (
    .A(SB_T0_NORTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1_enable),
    .Z(SB_T0_NORTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T0_SOUTH_SB_OUT_B17_ready_and (
    .A(SB_T0_SOUTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_OUT_B17_enable),
    .Z(SB_T0_SOUTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T0_SOUTH_SB_OUT_B1_ready_and (
    .A(SB_T0_SOUTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1_enable),
    .Z(SB_T0_SOUTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T0_WEST_SB_OUT_B17_ready_and (
    .A(SB_T0_WEST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_OUT_B17_enable),
    .Z(SB_T0_WEST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T0_WEST_SB_OUT_B1_ready_and (
    .A(SB_T0_WEST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1_enable),
    .Z(SB_T0_WEST_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T1_EAST_SB_OUT_B17_ready_and (
    .A(SB_T1_EAST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_OUT_B17_enable),
    .Z(SB_T1_EAST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T1_EAST_SB_OUT_B1_ready_and (
    .A(SB_T1_EAST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1_enable),
    .Z(SB_T1_EAST_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T1_NORTH_SB_OUT_B17_ready_and (
    .A(SB_T1_NORTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_OUT_B17_enable),
    .Z(SB_T1_NORTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T1_NORTH_SB_OUT_B1_ready_and (
    .A(SB_T1_NORTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1_enable),
    .Z(SB_T1_NORTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T1_SOUTH_SB_OUT_B17_ready_and (
    .A(SB_T1_SOUTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_OUT_B17_enable),
    .Z(SB_T1_SOUTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T1_SOUTH_SB_OUT_B1_ready_and (
    .A(SB_T1_SOUTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1_enable),
    .Z(SB_T1_SOUTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T1_WEST_SB_OUT_B17_ready_and (
    .A(SB_T1_WEST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_OUT_B17_enable),
    .Z(SB_T1_WEST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T1_WEST_SB_OUT_B1_ready_and (
    .A(SB_T1_WEST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1_enable),
    .Z(SB_T1_WEST_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T2_EAST_SB_OUT_B17_ready_and (
    .A(SB_T2_EAST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_OUT_B17_enable),
    .Z(SB_T2_EAST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T2_EAST_SB_OUT_B1_ready_and (
    .A(SB_T2_EAST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1_enable),
    .Z(SB_T2_EAST_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T2_NORTH_SB_OUT_B17_ready_and (
    .A(SB_T2_NORTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_OUT_B17_enable),
    .Z(SB_T2_NORTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T2_NORTH_SB_OUT_B1_ready_and (
    .A(SB_T2_NORTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1_enable),
    .Z(SB_T2_NORTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T2_SOUTH_SB_OUT_B17_ready_and (
    .A(SB_T2_SOUTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_OUT_B17_enable),
    .Z(SB_T2_SOUTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T2_SOUTH_SB_OUT_B1_ready_and (
    .A(SB_T2_SOUTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1_enable),
    .Z(SB_T2_SOUTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T2_WEST_SB_OUT_B17_ready_and (
    .A(SB_T2_WEST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_OUT_B17_enable),
    .Z(SB_T2_WEST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T2_WEST_SB_OUT_B1_ready_and (
    .A(SB_T2_WEST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1_enable),
    .Z(SB_T2_WEST_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T3_EAST_SB_OUT_B17_ready_and (
    .A(SB_T3_EAST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_OUT_B17_enable),
    .Z(SB_T3_EAST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T3_EAST_SB_OUT_B1_ready_and (
    .A(SB_T3_EAST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1_enable),
    .Z(SB_T3_EAST_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T3_NORTH_SB_OUT_B17_ready_and (
    .A(SB_T3_NORTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_OUT_B17_enable),
    .Z(SB_T3_NORTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T3_NORTH_SB_OUT_B1_ready_and (
    .A(SB_T3_NORTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1_enable),
    .Z(SB_T3_NORTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T3_SOUTH_SB_OUT_B17_ready_and (
    .A(SB_T3_SOUTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_OUT_B17_enable),
    .Z(SB_T3_SOUTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T3_SOUTH_SB_OUT_B1_ready_and (
    .A(SB_T3_SOUTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1_enable),
    .Z(SB_T3_SOUTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T3_WEST_SB_OUT_B17_ready_and (
    .A(SB_T3_WEST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_OUT_B17_enable),
    .Z(SB_T3_WEST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T3_WEST_SB_OUT_B1_ready_and (
    .A(SB_T3_WEST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1_enable),
    .Z(SB_T3_WEST_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T4_EAST_SB_OUT_B17_ready_and (
    .A(SB_T4_EAST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_OUT_B17_enable),
    .Z(SB_T4_EAST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T4_EAST_SB_OUT_B1_ready_and (
    .A(SB_T4_EAST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1_enable),
    .Z(SB_T4_EAST_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T4_NORTH_SB_OUT_B17_ready_and (
    .A(SB_T4_NORTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_OUT_B17_enable),
    .Z(SB_T4_NORTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T4_NORTH_SB_OUT_B1_ready_and (
    .A(SB_T4_NORTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1_enable),
    .Z(SB_T4_NORTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T4_SOUTH_SB_OUT_B17_ready_and (
    .A(SB_T4_SOUTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_OUT_B17_enable),
    .Z(SB_T4_SOUTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T4_SOUTH_SB_OUT_B1_ready_and (
    .A(SB_T4_SOUTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1_enable),
    .Z(SB_T4_SOUTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T4_WEST_SB_OUT_B17_ready_and (
    .A(SB_T4_WEST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_OUT_B17_enable),
    .Z(SB_T4_WEST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T4_WEST_SB_OUT_B1_ready_and (
    .A(SB_T4_WEST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1_enable),
    .Z(SB_T4_WEST_SB_OUT_B1_ready_and_Z)
);
corebit_and and_inst0 (
    .in0(coreir_eq_16_inst0_out),
    .in1(config_read[0]),
    .out(and_inst0_out)
);
corebit_and and_inst1 (
    .in0(coreir_eq_16_inst0_out),
    .in1(config_write[0]),
    .out(and_inst1_out)
);
corebit_const #(
    .value(1'b1)
) bit_const_1_None (
    .out(bit_const_1_None_out)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
coreir_const #(
    .value(9'h1ff),
    .width(9)
) const_511_9 (
    .out(const_511_9_out)
);
coreir_eq #(
    .width(16)
) coreir_eq_16_inst0 (
    .in0(tile_id),
    .in1(self_config_config_addr_out[15:0]),
    .out(coreir_eq_16_inst0_out)
);
coreir_wrap coreir_wrapOutClock_inst0 (
    .in(clk_pass_through),
    .out(coreir_wrapOutClock_inst0_out)
);
coreir_wrap coreir_wrapOutClock_inst1 (
    .in(clk_pass_through),
    .out(coreir_wrapOutClock_inst1_out)
);
wire [31:0] read_data_mux_I [15:0];
assign read_data_mux_I[15] = PowerDomainConfigReg_inst0_read_config_data;
assign read_data_mux_I[14] = SB_ID0_5TRACKS_B17_PE_read_config_data;
assign read_data_mux_I[13] = SB_ID0_5TRACKS_B1_PE_read_config_data;
assign read_data_mux_I[12] = CB_flush_read_config_data;
assign read_data_mux_I[11] = CB_PondTop_input_width_17_num_1_read_config_data;
assign read_data_mux_I[10] = CB_PondTop_input_width_17_num_0_read_config_data;
assign read_data_mux_I[9] = CB_PE_input_width_1_num_2_read_config_data;
assign read_data_mux_I[8] = CB_PE_input_width_1_num_1_read_config_data;
assign read_data_mux_I[7] = CB_PE_input_width_1_num_0_read_config_data;
assign read_data_mux_I[6] = CB_PE_input_width_17_num_3_read_config_data;
assign read_data_mux_I[5] = CB_PE_input_width_17_num_2_read_config_data;
assign read_data_mux_I[4] = CB_PE_input_width_17_num_1_read_config_data;
assign read_data_mux_I[3] = CB_PE_input_width_17_num_0_read_config_data;
assign read_data_mux_I[2] = PondCore_inst0_read_config_data_1;
assign read_data_mux_I[1] = PondCore_inst0_read_config_data;
assign read_data_mux_I[0] = PE_inst0_read_config_data;
MuxWithDefaultWrapper_16_32_8_0 read_data_mux (
    .I(read_data_mux_I),
    .S(self_config_config_addr_out[23:16]),
    .EN(and_inst0_out),
    .O(read_data_mux_O)
);
mantle_wire__typeBit32 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
assign SB_T0_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_IN_B17_ready_out;
assign SB_T0_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_IN_B1_ready_out;
assign SB_T0_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1;
assign SB_T0_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_OUT_B17;
assign SB_T0_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T0_EAST_SB_OUT_B17_valid_out;
assign SB_T0_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1_valid_out;
assign SB_T0_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_IN_B17_ready_out;
assign SB_T0_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_IN_B1_ready_out;
assign SB_T0_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1;
assign SB_T0_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_OUT_B17;
assign SB_T0_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T0_NORTH_SB_OUT_B17_valid_out;
assign SB_T0_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1_valid_out;
assign SB_T0_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_IN_B17_ready_out;
assign SB_T0_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_IN_B1_ready_out;
assign SB_T0_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1;
assign SB_T0_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_OUT_B17;
assign SB_T0_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T0_SOUTH_SB_OUT_B17_valid_out;
assign SB_T0_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1_valid_out;
assign SB_T0_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_IN_B17_ready_out;
assign SB_T0_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_IN_B1_ready_out;
assign SB_T0_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1;
assign SB_T0_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_OUT_B17;
assign SB_T0_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T0_WEST_SB_OUT_B17_valid_out;
assign SB_T0_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1_valid_out;
assign SB_T1_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_IN_B17_ready_out;
assign SB_T1_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_IN_B1_ready_out;
assign SB_T1_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1;
assign SB_T1_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_OUT_B17;
assign SB_T1_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T1_EAST_SB_OUT_B17_valid_out;
assign SB_T1_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1_valid_out;
assign SB_T1_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_IN_B17_ready_out;
assign SB_T1_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_IN_B1_ready_out;
assign SB_T1_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1;
assign SB_T1_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_OUT_B17;
assign SB_T1_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T1_NORTH_SB_OUT_B17_valid_out;
assign SB_T1_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1_valid_out;
assign SB_T1_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_IN_B17_ready_out;
assign SB_T1_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_IN_B1_ready_out;
assign SB_T1_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1;
assign SB_T1_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_OUT_B17;
assign SB_T1_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T1_SOUTH_SB_OUT_B17_valid_out;
assign SB_T1_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1_valid_out;
assign SB_T1_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_IN_B17_ready_out;
assign SB_T1_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_IN_B1_ready_out;
assign SB_T1_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1;
assign SB_T1_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_OUT_B17;
assign SB_T1_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T1_WEST_SB_OUT_B17_valid_out;
assign SB_T1_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1_valid_out;
assign SB_T2_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_IN_B17_ready_out;
assign SB_T2_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_IN_B1_ready_out;
assign SB_T2_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1;
assign SB_T2_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_OUT_B17;
assign SB_T2_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T2_EAST_SB_OUT_B17_valid_out;
assign SB_T2_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1_valid_out;
assign SB_T2_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_IN_B17_ready_out;
assign SB_T2_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_IN_B1_ready_out;
assign SB_T2_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1;
assign SB_T2_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_OUT_B17;
assign SB_T2_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T2_NORTH_SB_OUT_B17_valid_out;
assign SB_T2_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1_valid_out;
assign SB_T2_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_IN_B17_ready_out;
assign SB_T2_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_IN_B1_ready_out;
assign SB_T2_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1;
assign SB_T2_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_OUT_B17;
assign SB_T2_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T2_SOUTH_SB_OUT_B17_valid_out;
assign SB_T2_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1_valid_out;
assign SB_T2_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_IN_B17_ready_out;
assign SB_T2_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_IN_B1_ready_out;
assign SB_T2_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1;
assign SB_T2_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_OUT_B17;
assign SB_T2_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T2_WEST_SB_OUT_B17_valid_out;
assign SB_T2_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1_valid_out;
assign SB_T3_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_IN_B17_ready_out;
assign SB_T3_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_IN_B1_ready_out;
assign SB_T3_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1;
assign SB_T3_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_OUT_B17;
assign SB_T3_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T3_EAST_SB_OUT_B17_valid_out;
assign SB_T3_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1_valid_out;
assign SB_T3_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_IN_B17_ready_out;
assign SB_T3_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_IN_B1_ready_out;
assign SB_T3_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1;
assign SB_T3_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_OUT_B17;
assign SB_T3_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T3_NORTH_SB_OUT_B17_valid_out;
assign SB_T3_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1_valid_out;
assign SB_T3_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_IN_B17_ready_out;
assign SB_T3_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_IN_B1_ready_out;
assign SB_T3_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1;
assign SB_T3_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_OUT_B17;
assign SB_T3_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T3_SOUTH_SB_OUT_B17_valid_out;
assign SB_T3_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1_valid_out;
assign SB_T3_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_IN_B17_ready_out;
assign SB_T3_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_IN_B1_ready_out;
assign SB_T3_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1;
assign SB_T3_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_OUT_B17;
assign SB_T3_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T3_WEST_SB_OUT_B17_valid_out;
assign SB_T3_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1_valid_out;
assign SB_T4_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_IN_B17_ready_out;
assign SB_T4_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_IN_B1_ready_out;
assign SB_T4_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1;
assign SB_T4_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_OUT_B17;
assign SB_T4_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T4_EAST_SB_OUT_B17_valid_out;
assign SB_T4_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1_valid_out;
assign SB_T4_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_IN_B17_ready_out;
assign SB_T4_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_IN_B1_ready_out;
assign SB_T4_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1;
assign SB_T4_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_OUT_B17;
assign SB_T4_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T4_NORTH_SB_OUT_B17_valid_out;
assign SB_T4_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1_valid_out;
assign SB_T4_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_IN_B17_ready_out;
assign SB_T4_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_IN_B1_ready_out;
assign SB_T4_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1;
assign SB_T4_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_OUT_B17;
assign SB_T4_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T4_SOUTH_SB_OUT_B17_valid_out;
assign SB_T4_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1_valid_out;
assign SB_T4_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_IN_B17_ready_out;
assign SB_T4_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_IN_B1_ready_out;
assign SB_T4_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1;
assign SB_T4_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_OUT_B17;
assign SB_T4_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_PE_SB_T4_WEST_SB_OUT_B17_valid_out;
assign SB_T4_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1_valid_out;
assign clk_out = coreir_wrapOutClock_inst0_out;
assign clk_pass_through_out_bot = clk_pass_through;
assign clk_pass_through_out_right = coreir_wrapOutClock_inst1_out;
assign config_out_config_addr = config_config_addr;
assign config_out_config_data = config_config_data;
assign config_out_read = config_read;
assign config_out_write = config_write;
assign flush_out = flush;
assign hi = const_511_9_out;
assign lo = const_0_8_out;
assign read_config_data = PowerDomainOR_O;
assign reset_out = reset;
assign stall_out = stall;
endmodule

module CB_MEM_input_width_1_num_1 (
    input [0:0] I [19:0],
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output enable,
    output [31:0] out_sel,
    output [31:0] read_config_data,
    input ready_in,
    output ready_out,
    input reset,
    input [19:0] valid_in,
    output valid_out
);
wire [0:0] CB_MEM_input_width_1_num_1_O;
wire CB_MEM_input_width_1_num_1_ready_out;
wire CB_MEM_input_width_1_num_1_valid_out;
wire [31:0] CB_MEM_input_width_1_num_1_out_sel;
wire [0:0] CB_MEM_input_width_1_num_1_enable_value_O;
wire [4:0] CB_MEM_input_width_1_num_1_sel_value_O;
wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
wire [5:0] config_reg_0_O;
wire [0:0] CB_MEM_input_width_1_num_1_I [19:0];
assign CB_MEM_input_width_1_num_1_I[19] = I[19];
assign CB_MEM_input_width_1_num_1_I[18] = I[18];
assign CB_MEM_input_width_1_num_1_I[17] = I[17];
assign CB_MEM_input_width_1_num_1_I[16] = I[16];
assign CB_MEM_input_width_1_num_1_I[15] = I[15];
assign CB_MEM_input_width_1_num_1_I[14] = I[14];
assign CB_MEM_input_width_1_num_1_I[13] = I[13];
assign CB_MEM_input_width_1_num_1_I[12] = I[12];
assign CB_MEM_input_width_1_num_1_I[11] = I[11];
assign CB_MEM_input_width_1_num_1_I[10] = I[10];
assign CB_MEM_input_width_1_num_1_I[9] = I[9];
assign CB_MEM_input_width_1_num_1_I[8] = I[8];
assign CB_MEM_input_width_1_num_1_I[7] = I[7];
assign CB_MEM_input_width_1_num_1_I[6] = I[6];
assign CB_MEM_input_width_1_num_1_I[5] = I[5];
assign CB_MEM_input_width_1_num_1_I[4] = I[4];
assign CB_MEM_input_width_1_num_1_I[3] = I[3];
assign CB_MEM_input_width_1_num_1_I[2] = I[2];
assign CB_MEM_input_width_1_num_1_I[1] = I[1];
assign CB_MEM_input_width_1_num_1_I[0] = I[0];
mux_aoi_ready_valid_const_20_1 CB_MEM_input_width_1_num_1 (
    .I(CB_MEM_input_width_1_num_1_I),
    .O(CB_MEM_input_width_1_num_1_O),
    .ready_in(ready_in),
    .ready_out(CB_MEM_input_width_1_num_1_ready_out),
    .valid_in(valid_in),
    .valid_out(CB_MEM_input_width_1_num_1_valid_out),
    .S(CB_MEM_input_width_1_num_1_sel_value_O),
    .out_sel(CB_MEM_input_width_1_num_1_out_sel)
);
SliceWrapper_6_0_1 CB_MEM_input_width_1_num_1_enable_value (
    .I(config_reg_0_O),
    .O(CB_MEM_input_width_1_num_1_enable_value_O)
);
SliceWrapper_6_1_6 CB_MEM_input_width_1_num_1_sel_value (
    .I(config_reg_0_O),
    .O(CB_MEM_input_width_1_num_1_sel_value_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_6_32_inst0$bit_const_0_None (
    .out(ZextWrapper_6_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O (
    .in(ZextWrapper_6_32_inst0$self_O_in),
    .out(ZextWrapper_6_32_inst0$self_O_out)
);
ConfigRegister_6_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_MEM_input_width_1_num_1_O;
assign enable = CB_MEM_input_width_1_num_1_enable_value_O[0];
assign out_sel = CB_MEM_input_width_1_num_1_out_sel;
assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
assign ready_out = CB_MEM_input_width_1_num_1_ready_out;
assign valid_out = CB_MEM_input_width_1_num_1_valid_out;
endmodule

module CB_MEM_input_width_1_num_0 (
    input [0:0] I [19:0],
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output enable,
    output [31:0] out_sel,
    output [31:0] read_config_data,
    input ready_in,
    output ready_out,
    input reset,
    input [19:0] valid_in,
    output valid_out
);
wire [0:0] CB_MEM_input_width_1_num_0_O;
wire CB_MEM_input_width_1_num_0_ready_out;
wire CB_MEM_input_width_1_num_0_valid_out;
wire [31:0] CB_MEM_input_width_1_num_0_out_sel;
wire [0:0] CB_MEM_input_width_1_num_0_enable_value_O;
wire [4:0] CB_MEM_input_width_1_num_0_sel_value_O;
wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
wire [5:0] config_reg_0_O;
wire [0:0] CB_MEM_input_width_1_num_0_I [19:0];
assign CB_MEM_input_width_1_num_0_I[19] = I[19];
assign CB_MEM_input_width_1_num_0_I[18] = I[18];
assign CB_MEM_input_width_1_num_0_I[17] = I[17];
assign CB_MEM_input_width_1_num_0_I[16] = I[16];
assign CB_MEM_input_width_1_num_0_I[15] = I[15];
assign CB_MEM_input_width_1_num_0_I[14] = I[14];
assign CB_MEM_input_width_1_num_0_I[13] = I[13];
assign CB_MEM_input_width_1_num_0_I[12] = I[12];
assign CB_MEM_input_width_1_num_0_I[11] = I[11];
assign CB_MEM_input_width_1_num_0_I[10] = I[10];
assign CB_MEM_input_width_1_num_0_I[9] = I[9];
assign CB_MEM_input_width_1_num_0_I[8] = I[8];
assign CB_MEM_input_width_1_num_0_I[7] = I[7];
assign CB_MEM_input_width_1_num_0_I[6] = I[6];
assign CB_MEM_input_width_1_num_0_I[5] = I[5];
assign CB_MEM_input_width_1_num_0_I[4] = I[4];
assign CB_MEM_input_width_1_num_0_I[3] = I[3];
assign CB_MEM_input_width_1_num_0_I[2] = I[2];
assign CB_MEM_input_width_1_num_0_I[1] = I[1];
assign CB_MEM_input_width_1_num_0_I[0] = I[0];
mux_aoi_ready_valid_const_20_1 CB_MEM_input_width_1_num_0 (
    .I(CB_MEM_input_width_1_num_0_I),
    .O(CB_MEM_input_width_1_num_0_O),
    .ready_in(ready_in),
    .ready_out(CB_MEM_input_width_1_num_0_ready_out),
    .valid_in(valid_in),
    .valid_out(CB_MEM_input_width_1_num_0_valid_out),
    .S(CB_MEM_input_width_1_num_0_sel_value_O),
    .out_sel(CB_MEM_input_width_1_num_0_out_sel)
);
SliceWrapper_6_0_1 CB_MEM_input_width_1_num_0_enable_value (
    .I(config_reg_0_O),
    .O(CB_MEM_input_width_1_num_0_enable_value_O)
);
SliceWrapper_6_1_6 CB_MEM_input_width_1_num_0_sel_value (
    .I(config_reg_0_O),
    .O(CB_MEM_input_width_1_num_0_sel_value_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_6_32_inst0$bit_const_0_None (
    .out(ZextWrapper_6_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O (
    .in(ZextWrapper_6_32_inst0$self_O_in),
    .out(ZextWrapper_6_32_inst0$self_O_out)
);
ConfigRegister_6_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_MEM_input_width_1_num_0_O;
assign enable = CB_MEM_input_width_1_num_0_enable_value_O[0];
assign out_sel = CB_MEM_input_width_1_num_0_out_sel;
assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
assign ready_out = CB_MEM_input_width_1_num_0_ready_out;
assign valid_out = CB_MEM_input_width_1_num_0_valid_out;
endmodule

module CB_MEM_input_width_17_num_3 (
    input [16:0] I [19:0],
    output [16:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output enable,
    output [31:0] out_sel,
    output [31:0] read_config_data,
    input ready_in,
    output ready_out,
    input reset,
    input [19:0] valid_in,
    output valid_out
);
wire [16:0] CB_MEM_input_width_17_num_3_O;
wire CB_MEM_input_width_17_num_3_ready_out;
wire CB_MEM_input_width_17_num_3_valid_out;
wire [31:0] CB_MEM_input_width_17_num_3_out_sel;
wire [0:0] CB_MEM_input_width_17_num_3_enable_value_O;
wire [4:0] CB_MEM_input_width_17_num_3_sel_value_O;
wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
wire [5:0] config_reg_0_O;
wire [16:0] CB_MEM_input_width_17_num_3_I [19:0];
assign CB_MEM_input_width_17_num_3_I[19] = I[19];
assign CB_MEM_input_width_17_num_3_I[18] = I[18];
assign CB_MEM_input_width_17_num_3_I[17] = I[17];
assign CB_MEM_input_width_17_num_3_I[16] = I[16];
assign CB_MEM_input_width_17_num_3_I[15] = I[15];
assign CB_MEM_input_width_17_num_3_I[14] = I[14];
assign CB_MEM_input_width_17_num_3_I[13] = I[13];
assign CB_MEM_input_width_17_num_3_I[12] = I[12];
assign CB_MEM_input_width_17_num_3_I[11] = I[11];
assign CB_MEM_input_width_17_num_3_I[10] = I[10];
assign CB_MEM_input_width_17_num_3_I[9] = I[9];
assign CB_MEM_input_width_17_num_3_I[8] = I[8];
assign CB_MEM_input_width_17_num_3_I[7] = I[7];
assign CB_MEM_input_width_17_num_3_I[6] = I[6];
assign CB_MEM_input_width_17_num_3_I[5] = I[5];
assign CB_MEM_input_width_17_num_3_I[4] = I[4];
assign CB_MEM_input_width_17_num_3_I[3] = I[3];
assign CB_MEM_input_width_17_num_3_I[2] = I[2];
assign CB_MEM_input_width_17_num_3_I[1] = I[1];
assign CB_MEM_input_width_17_num_3_I[0] = I[0];
mux_aoi_ready_valid_const_20_17 CB_MEM_input_width_17_num_3 (
    .I(CB_MEM_input_width_17_num_3_I),
    .O(CB_MEM_input_width_17_num_3_O),
    .ready_in(ready_in),
    .ready_out(CB_MEM_input_width_17_num_3_ready_out),
    .valid_in(valid_in),
    .valid_out(CB_MEM_input_width_17_num_3_valid_out),
    .S(CB_MEM_input_width_17_num_3_sel_value_O),
    .out_sel(CB_MEM_input_width_17_num_3_out_sel)
);
SliceWrapper_6_0_1 CB_MEM_input_width_17_num_3_enable_value (
    .I(config_reg_0_O),
    .O(CB_MEM_input_width_17_num_3_enable_value_O)
);
SliceWrapper_6_1_6 CB_MEM_input_width_17_num_3_sel_value (
    .I(config_reg_0_O),
    .O(CB_MEM_input_width_17_num_3_sel_value_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_6_32_inst0$bit_const_0_None (
    .out(ZextWrapper_6_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O (
    .in(ZextWrapper_6_32_inst0$self_O_in),
    .out(ZextWrapper_6_32_inst0$self_O_out)
);
ConfigRegister_6_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_MEM_input_width_17_num_3_O;
assign enable = CB_MEM_input_width_17_num_3_enable_value_O[0];
assign out_sel = CB_MEM_input_width_17_num_3_out_sel;
assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
assign ready_out = CB_MEM_input_width_17_num_3_ready_out;
assign valid_out = CB_MEM_input_width_17_num_3_valid_out;
endmodule

module CB_MEM_input_width_17_num_2 (
    input [16:0] I [19:0],
    output [16:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output enable,
    output [31:0] out_sel,
    output [31:0] read_config_data,
    input ready_in,
    output ready_out,
    input reset,
    input [19:0] valid_in,
    output valid_out
);
wire [16:0] CB_MEM_input_width_17_num_2_O;
wire CB_MEM_input_width_17_num_2_ready_out;
wire CB_MEM_input_width_17_num_2_valid_out;
wire [31:0] CB_MEM_input_width_17_num_2_out_sel;
wire [0:0] CB_MEM_input_width_17_num_2_enable_value_O;
wire [4:0] CB_MEM_input_width_17_num_2_sel_value_O;
wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
wire [5:0] config_reg_0_O;
wire [16:0] CB_MEM_input_width_17_num_2_I [19:0];
assign CB_MEM_input_width_17_num_2_I[19] = I[19];
assign CB_MEM_input_width_17_num_2_I[18] = I[18];
assign CB_MEM_input_width_17_num_2_I[17] = I[17];
assign CB_MEM_input_width_17_num_2_I[16] = I[16];
assign CB_MEM_input_width_17_num_2_I[15] = I[15];
assign CB_MEM_input_width_17_num_2_I[14] = I[14];
assign CB_MEM_input_width_17_num_2_I[13] = I[13];
assign CB_MEM_input_width_17_num_2_I[12] = I[12];
assign CB_MEM_input_width_17_num_2_I[11] = I[11];
assign CB_MEM_input_width_17_num_2_I[10] = I[10];
assign CB_MEM_input_width_17_num_2_I[9] = I[9];
assign CB_MEM_input_width_17_num_2_I[8] = I[8];
assign CB_MEM_input_width_17_num_2_I[7] = I[7];
assign CB_MEM_input_width_17_num_2_I[6] = I[6];
assign CB_MEM_input_width_17_num_2_I[5] = I[5];
assign CB_MEM_input_width_17_num_2_I[4] = I[4];
assign CB_MEM_input_width_17_num_2_I[3] = I[3];
assign CB_MEM_input_width_17_num_2_I[2] = I[2];
assign CB_MEM_input_width_17_num_2_I[1] = I[1];
assign CB_MEM_input_width_17_num_2_I[0] = I[0];
mux_aoi_ready_valid_const_20_17 CB_MEM_input_width_17_num_2 (
    .I(CB_MEM_input_width_17_num_2_I),
    .O(CB_MEM_input_width_17_num_2_O),
    .ready_in(ready_in),
    .ready_out(CB_MEM_input_width_17_num_2_ready_out),
    .valid_in(valid_in),
    .valid_out(CB_MEM_input_width_17_num_2_valid_out),
    .S(CB_MEM_input_width_17_num_2_sel_value_O),
    .out_sel(CB_MEM_input_width_17_num_2_out_sel)
);
SliceWrapper_6_0_1 CB_MEM_input_width_17_num_2_enable_value (
    .I(config_reg_0_O),
    .O(CB_MEM_input_width_17_num_2_enable_value_O)
);
SliceWrapper_6_1_6 CB_MEM_input_width_17_num_2_sel_value (
    .I(config_reg_0_O),
    .O(CB_MEM_input_width_17_num_2_sel_value_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_6_32_inst0$bit_const_0_None (
    .out(ZextWrapper_6_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O (
    .in(ZextWrapper_6_32_inst0$self_O_in),
    .out(ZextWrapper_6_32_inst0$self_O_out)
);
ConfigRegister_6_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_MEM_input_width_17_num_2_O;
assign enable = CB_MEM_input_width_17_num_2_enable_value_O[0];
assign out_sel = CB_MEM_input_width_17_num_2_out_sel;
assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
assign ready_out = CB_MEM_input_width_17_num_2_ready_out;
assign valid_out = CB_MEM_input_width_17_num_2_valid_out;
endmodule

module CB_MEM_input_width_17_num_1 (
    input [16:0] I [19:0],
    output [16:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output enable,
    output [31:0] out_sel,
    output [31:0] read_config_data,
    input ready_in,
    output ready_out,
    input reset,
    input [19:0] valid_in,
    output valid_out
);
wire [16:0] CB_MEM_input_width_17_num_1_O;
wire CB_MEM_input_width_17_num_1_ready_out;
wire CB_MEM_input_width_17_num_1_valid_out;
wire [31:0] CB_MEM_input_width_17_num_1_out_sel;
wire [0:0] CB_MEM_input_width_17_num_1_enable_value_O;
wire [4:0] CB_MEM_input_width_17_num_1_sel_value_O;
wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
wire [5:0] config_reg_0_O;
wire [16:0] CB_MEM_input_width_17_num_1_I [19:0];
assign CB_MEM_input_width_17_num_1_I[19] = I[19];
assign CB_MEM_input_width_17_num_1_I[18] = I[18];
assign CB_MEM_input_width_17_num_1_I[17] = I[17];
assign CB_MEM_input_width_17_num_1_I[16] = I[16];
assign CB_MEM_input_width_17_num_1_I[15] = I[15];
assign CB_MEM_input_width_17_num_1_I[14] = I[14];
assign CB_MEM_input_width_17_num_1_I[13] = I[13];
assign CB_MEM_input_width_17_num_1_I[12] = I[12];
assign CB_MEM_input_width_17_num_1_I[11] = I[11];
assign CB_MEM_input_width_17_num_1_I[10] = I[10];
assign CB_MEM_input_width_17_num_1_I[9] = I[9];
assign CB_MEM_input_width_17_num_1_I[8] = I[8];
assign CB_MEM_input_width_17_num_1_I[7] = I[7];
assign CB_MEM_input_width_17_num_1_I[6] = I[6];
assign CB_MEM_input_width_17_num_1_I[5] = I[5];
assign CB_MEM_input_width_17_num_1_I[4] = I[4];
assign CB_MEM_input_width_17_num_1_I[3] = I[3];
assign CB_MEM_input_width_17_num_1_I[2] = I[2];
assign CB_MEM_input_width_17_num_1_I[1] = I[1];
assign CB_MEM_input_width_17_num_1_I[0] = I[0];
mux_aoi_ready_valid_const_20_17 CB_MEM_input_width_17_num_1 (
    .I(CB_MEM_input_width_17_num_1_I),
    .O(CB_MEM_input_width_17_num_1_O),
    .ready_in(ready_in),
    .ready_out(CB_MEM_input_width_17_num_1_ready_out),
    .valid_in(valid_in),
    .valid_out(CB_MEM_input_width_17_num_1_valid_out),
    .S(CB_MEM_input_width_17_num_1_sel_value_O),
    .out_sel(CB_MEM_input_width_17_num_1_out_sel)
);
SliceWrapper_6_0_1 CB_MEM_input_width_17_num_1_enable_value (
    .I(config_reg_0_O),
    .O(CB_MEM_input_width_17_num_1_enable_value_O)
);
SliceWrapper_6_1_6 CB_MEM_input_width_17_num_1_sel_value (
    .I(config_reg_0_O),
    .O(CB_MEM_input_width_17_num_1_sel_value_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_6_32_inst0$bit_const_0_None (
    .out(ZextWrapper_6_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O (
    .in(ZextWrapper_6_32_inst0$self_O_in),
    .out(ZextWrapper_6_32_inst0$self_O_out)
);
ConfigRegister_6_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_MEM_input_width_17_num_1_O;
assign enable = CB_MEM_input_width_17_num_1_enable_value_O[0];
assign out_sel = CB_MEM_input_width_17_num_1_out_sel;
assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
assign ready_out = CB_MEM_input_width_17_num_1_ready_out;
assign valid_out = CB_MEM_input_width_17_num_1_valid_out;
endmodule

module CB_MEM_input_width_17_num_0 (
    input [16:0] I [19:0],
    output [16:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output enable,
    output [31:0] out_sel,
    output [31:0] read_config_data,
    input ready_in,
    output ready_out,
    input reset,
    input [19:0] valid_in,
    output valid_out
);
wire [16:0] CB_MEM_input_width_17_num_0_O;
wire CB_MEM_input_width_17_num_0_ready_out;
wire CB_MEM_input_width_17_num_0_valid_out;
wire [31:0] CB_MEM_input_width_17_num_0_out_sel;
wire [0:0] CB_MEM_input_width_17_num_0_enable_value_O;
wire [4:0] CB_MEM_input_width_17_num_0_sel_value_O;
wire ZextWrapper_6_32_inst0$bit_const_0_None_out;
wire [31:0] ZextWrapper_6_32_inst0$self_O_in;
wire [5:0] config_reg_0_O;
wire [16:0] CB_MEM_input_width_17_num_0_I [19:0];
assign CB_MEM_input_width_17_num_0_I[19] = I[19];
assign CB_MEM_input_width_17_num_0_I[18] = I[18];
assign CB_MEM_input_width_17_num_0_I[17] = I[17];
assign CB_MEM_input_width_17_num_0_I[16] = I[16];
assign CB_MEM_input_width_17_num_0_I[15] = I[15];
assign CB_MEM_input_width_17_num_0_I[14] = I[14];
assign CB_MEM_input_width_17_num_0_I[13] = I[13];
assign CB_MEM_input_width_17_num_0_I[12] = I[12];
assign CB_MEM_input_width_17_num_0_I[11] = I[11];
assign CB_MEM_input_width_17_num_0_I[10] = I[10];
assign CB_MEM_input_width_17_num_0_I[9] = I[9];
assign CB_MEM_input_width_17_num_0_I[8] = I[8];
assign CB_MEM_input_width_17_num_0_I[7] = I[7];
assign CB_MEM_input_width_17_num_0_I[6] = I[6];
assign CB_MEM_input_width_17_num_0_I[5] = I[5];
assign CB_MEM_input_width_17_num_0_I[4] = I[4];
assign CB_MEM_input_width_17_num_0_I[3] = I[3];
assign CB_MEM_input_width_17_num_0_I[2] = I[2];
assign CB_MEM_input_width_17_num_0_I[1] = I[1];
assign CB_MEM_input_width_17_num_0_I[0] = I[0];
mux_aoi_ready_valid_const_20_17 CB_MEM_input_width_17_num_0 (
    .I(CB_MEM_input_width_17_num_0_I),
    .O(CB_MEM_input_width_17_num_0_O),
    .ready_in(ready_in),
    .ready_out(CB_MEM_input_width_17_num_0_ready_out),
    .valid_in(valid_in),
    .valid_out(CB_MEM_input_width_17_num_0_valid_out),
    .S(CB_MEM_input_width_17_num_0_sel_value_O),
    .out_sel(CB_MEM_input_width_17_num_0_out_sel)
);
SliceWrapper_6_0_1 CB_MEM_input_width_17_num_0_enable_value (
    .I(config_reg_0_O),
    .O(CB_MEM_input_width_17_num_0_enable_value_O)
);
SliceWrapper_6_1_6 CB_MEM_input_width_17_num_0_sel_value (
    .I(config_reg_0_O),
    .O(CB_MEM_input_width_17_num_0_sel_value_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_6_32_inst0$bit_const_0_None (
    .out(ZextWrapper_6_32_inst0$bit_const_0_None_out)
);
wire [31:0] ZextWrapper_6_32_inst0$self_O_out;
assign ZextWrapper_6_32_inst0$self_O_out = {ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,ZextWrapper_6_32_inst0$bit_const_0_None_out,config_reg_0_O};
mantle_wire__typeBitIn32 ZextWrapper_6_32_inst0$self_O (
    .in(ZextWrapper_6_32_inst0$self_O_in),
    .out(ZextWrapper_6_32_inst0$self_O_out)
);
ConfigRegister_6_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = CB_MEM_input_width_17_num_0_O;
assign enable = CB_MEM_input_width_17_num_0_enable_value_O[0];
assign out_sel = CB_MEM_input_width_17_num_0_out_sel;
assign read_config_data = ZextWrapper_6_32_inst0$self_O_in;
assign ready_out = CB_MEM_input_width_17_num_0_ready_out;
assign valid_out = CB_MEM_input_width_17_num_0_valid_out;
endmodule

module Tile_MemCore (
    input [0:0] SB_T0_EAST_SB_IN_B1,
    input [16:0] SB_T0_EAST_SB_IN_B17,
    output SB_T0_EAST_SB_IN_B17_ready,
    input SB_T0_EAST_SB_IN_B17_valid,
    output SB_T0_EAST_SB_IN_B1_ready,
    input SB_T0_EAST_SB_IN_B1_valid,
    output [0:0] SB_T0_EAST_SB_OUT_B1,
    output [16:0] SB_T0_EAST_SB_OUT_B17,
    input SB_T0_EAST_SB_OUT_B17_ready,
    output SB_T0_EAST_SB_OUT_B17_valid,
    input SB_T0_EAST_SB_OUT_B1_ready,
    output SB_T0_EAST_SB_OUT_B1_valid,
    input [0:0] SB_T0_NORTH_SB_IN_B1,
    input [16:0] SB_T0_NORTH_SB_IN_B17,
    output SB_T0_NORTH_SB_IN_B17_ready,
    input SB_T0_NORTH_SB_IN_B17_valid,
    output SB_T0_NORTH_SB_IN_B1_ready,
    input SB_T0_NORTH_SB_IN_B1_valid,
    output [0:0] SB_T0_NORTH_SB_OUT_B1,
    output [16:0] SB_T0_NORTH_SB_OUT_B17,
    input SB_T0_NORTH_SB_OUT_B17_ready,
    output SB_T0_NORTH_SB_OUT_B17_valid,
    input SB_T0_NORTH_SB_OUT_B1_ready,
    output SB_T0_NORTH_SB_OUT_B1_valid,
    input [0:0] SB_T0_SOUTH_SB_IN_B1,
    input [16:0] SB_T0_SOUTH_SB_IN_B17,
    output SB_T0_SOUTH_SB_IN_B17_ready,
    input SB_T0_SOUTH_SB_IN_B17_valid,
    output SB_T0_SOUTH_SB_IN_B1_ready,
    input SB_T0_SOUTH_SB_IN_B1_valid,
    output [0:0] SB_T0_SOUTH_SB_OUT_B1,
    output [16:0] SB_T0_SOUTH_SB_OUT_B17,
    input SB_T0_SOUTH_SB_OUT_B17_ready,
    output SB_T0_SOUTH_SB_OUT_B17_valid,
    input SB_T0_SOUTH_SB_OUT_B1_ready,
    output SB_T0_SOUTH_SB_OUT_B1_valid,
    input [0:0] SB_T0_WEST_SB_IN_B1,
    input [16:0] SB_T0_WEST_SB_IN_B17,
    output SB_T0_WEST_SB_IN_B17_ready,
    input SB_T0_WEST_SB_IN_B17_valid,
    output SB_T0_WEST_SB_IN_B1_ready,
    input SB_T0_WEST_SB_IN_B1_valid,
    output [0:0] SB_T0_WEST_SB_OUT_B1,
    output [16:0] SB_T0_WEST_SB_OUT_B17,
    input SB_T0_WEST_SB_OUT_B17_ready,
    output SB_T0_WEST_SB_OUT_B17_valid,
    input SB_T0_WEST_SB_OUT_B1_ready,
    output SB_T0_WEST_SB_OUT_B1_valid,
    input [0:0] SB_T1_EAST_SB_IN_B1,
    input [16:0] SB_T1_EAST_SB_IN_B17,
    output SB_T1_EAST_SB_IN_B17_ready,
    input SB_T1_EAST_SB_IN_B17_valid,
    output SB_T1_EAST_SB_IN_B1_ready,
    input SB_T1_EAST_SB_IN_B1_valid,
    output [0:0] SB_T1_EAST_SB_OUT_B1,
    output [16:0] SB_T1_EAST_SB_OUT_B17,
    input SB_T1_EAST_SB_OUT_B17_ready,
    output SB_T1_EAST_SB_OUT_B17_valid,
    input SB_T1_EAST_SB_OUT_B1_ready,
    output SB_T1_EAST_SB_OUT_B1_valid,
    input [0:0] SB_T1_NORTH_SB_IN_B1,
    input [16:0] SB_T1_NORTH_SB_IN_B17,
    output SB_T1_NORTH_SB_IN_B17_ready,
    input SB_T1_NORTH_SB_IN_B17_valid,
    output SB_T1_NORTH_SB_IN_B1_ready,
    input SB_T1_NORTH_SB_IN_B1_valid,
    output [0:0] SB_T1_NORTH_SB_OUT_B1,
    output [16:0] SB_T1_NORTH_SB_OUT_B17,
    input SB_T1_NORTH_SB_OUT_B17_ready,
    output SB_T1_NORTH_SB_OUT_B17_valid,
    input SB_T1_NORTH_SB_OUT_B1_ready,
    output SB_T1_NORTH_SB_OUT_B1_valid,
    input [0:0] SB_T1_SOUTH_SB_IN_B1,
    input [16:0] SB_T1_SOUTH_SB_IN_B17,
    output SB_T1_SOUTH_SB_IN_B17_ready,
    input SB_T1_SOUTH_SB_IN_B17_valid,
    output SB_T1_SOUTH_SB_IN_B1_ready,
    input SB_T1_SOUTH_SB_IN_B1_valid,
    output [0:0] SB_T1_SOUTH_SB_OUT_B1,
    output [16:0] SB_T1_SOUTH_SB_OUT_B17,
    input SB_T1_SOUTH_SB_OUT_B17_ready,
    output SB_T1_SOUTH_SB_OUT_B17_valid,
    input SB_T1_SOUTH_SB_OUT_B1_ready,
    output SB_T1_SOUTH_SB_OUT_B1_valid,
    input [0:0] SB_T1_WEST_SB_IN_B1,
    input [16:0] SB_T1_WEST_SB_IN_B17,
    output SB_T1_WEST_SB_IN_B17_ready,
    input SB_T1_WEST_SB_IN_B17_valid,
    output SB_T1_WEST_SB_IN_B1_ready,
    input SB_T1_WEST_SB_IN_B1_valid,
    output [0:0] SB_T1_WEST_SB_OUT_B1,
    output [16:0] SB_T1_WEST_SB_OUT_B17,
    input SB_T1_WEST_SB_OUT_B17_ready,
    output SB_T1_WEST_SB_OUT_B17_valid,
    input SB_T1_WEST_SB_OUT_B1_ready,
    output SB_T1_WEST_SB_OUT_B1_valid,
    input [0:0] SB_T2_EAST_SB_IN_B1,
    input [16:0] SB_T2_EAST_SB_IN_B17,
    output SB_T2_EAST_SB_IN_B17_ready,
    input SB_T2_EAST_SB_IN_B17_valid,
    output SB_T2_EAST_SB_IN_B1_ready,
    input SB_T2_EAST_SB_IN_B1_valid,
    output [0:0] SB_T2_EAST_SB_OUT_B1,
    output [16:0] SB_T2_EAST_SB_OUT_B17,
    input SB_T2_EAST_SB_OUT_B17_ready,
    output SB_T2_EAST_SB_OUT_B17_valid,
    input SB_T2_EAST_SB_OUT_B1_ready,
    output SB_T2_EAST_SB_OUT_B1_valid,
    input [0:0] SB_T2_NORTH_SB_IN_B1,
    input [16:0] SB_T2_NORTH_SB_IN_B17,
    output SB_T2_NORTH_SB_IN_B17_ready,
    input SB_T2_NORTH_SB_IN_B17_valid,
    output SB_T2_NORTH_SB_IN_B1_ready,
    input SB_T2_NORTH_SB_IN_B1_valid,
    output [0:0] SB_T2_NORTH_SB_OUT_B1,
    output [16:0] SB_T2_NORTH_SB_OUT_B17,
    input SB_T2_NORTH_SB_OUT_B17_ready,
    output SB_T2_NORTH_SB_OUT_B17_valid,
    input SB_T2_NORTH_SB_OUT_B1_ready,
    output SB_T2_NORTH_SB_OUT_B1_valid,
    input [0:0] SB_T2_SOUTH_SB_IN_B1,
    input [16:0] SB_T2_SOUTH_SB_IN_B17,
    output SB_T2_SOUTH_SB_IN_B17_ready,
    input SB_T2_SOUTH_SB_IN_B17_valid,
    output SB_T2_SOUTH_SB_IN_B1_ready,
    input SB_T2_SOUTH_SB_IN_B1_valid,
    output [0:0] SB_T2_SOUTH_SB_OUT_B1,
    output [16:0] SB_T2_SOUTH_SB_OUT_B17,
    input SB_T2_SOUTH_SB_OUT_B17_ready,
    output SB_T2_SOUTH_SB_OUT_B17_valid,
    input SB_T2_SOUTH_SB_OUT_B1_ready,
    output SB_T2_SOUTH_SB_OUT_B1_valid,
    input [0:0] SB_T2_WEST_SB_IN_B1,
    input [16:0] SB_T2_WEST_SB_IN_B17,
    output SB_T2_WEST_SB_IN_B17_ready,
    input SB_T2_WEST_SB_IN_B17_valid,
    output SB_T2_WEST_SB_IN_B1_ready,
    input SB_T2_WEST_SB_IN_B1_valid,
    output [0:0] SB_T2_WEST_SB_OUT_B1,
    output [16:0] SB_T2_WEST_SB_OUT_B17,
    input SB_T2_WEST_SB_OUT_B17_ready,
    output SB_T2_WEST_SB_OUT_B17_valid,
    input SB_T2_WEST_SB_OUT_B1_ready,
    output SB_T2_WEST_SB_OUT_B1_valid,
    input [0:0] SB_T3_EAST_SB_IN_B1,
    input [16:0] SB_T3_EAST_SB_IN_B17,
    output SB_T3_EAST_SB_IN_B17_ready,
    input SB_T3_EAST_SB_IN_B17_valid,
    output SB_T3_EAST_SB_IN_B1_ready,
    input SB_T3_EAST_SB_IN_B1_valid,
    output [0:0] SB_T3_EAST_SB_OUT_B1,
    output [16:0] SB_T3_EAST_SB_OUT_B17,
    input SB_T3_EAST_SB_OUT_B17_ready,
    output SB_T3_EAST_SB_OUT_B17_valid,
    input SB_T3_EAST_SB_OUT_B1_ready,
    output SB_T3_EAST_SB_OUT_B1_valid,
    input [0:0] SB_T3_NORTH_SB_IN_B1,
    input [16:0] SB_T3_NORTH_SB_IN_B17,
    output SB_T3_NORTH_SB_IN_B17_ready,
    input SB_T3_NORTH_SB_IN_B17_valid,
    output SB_T3_NORTH_SB_IN_B1_ready,
    input SB_T3_NORTH_SB_IN_B1_valid,
    output [0:0] SB_T3_NORTH_SB_OUT_B1,
    output [16:0] SB_T3_NORTH_SB_OUT_B17,
    input SB_T3_NORTH_SB_OUT_B17_ready,
    output SB_T3_NORTH_SB_OUT_B17_valid,
    input SB_T3_NORTH_SB_OUT_B1_ready,
    output SB_T3_NORTH_SB_OUT_B1_valid,
    input [0:0] SB_T3_SOUTH_SB_IN_B1,
    input [16:0] SB_T3_SOUTH_SB_IN_B17,
    output SB_T3_SOUTH_SB_IN_B17_ready,
    input SB_T3_SOUTH_SB_IN_B17_valid,
    output SB_T3_SOUTH_SB_IN_B1_ready,
    input SB_T3_SOUTH_SB_IN_B1_valid,
    output [0:0] SB_T3_SOUTH_SB_OUT_B1,
    output [16:0] SB_T3_SOUTH_SB_OUT_B17,
    input SB_T3_SOUTH_SB_OUT_B17_ready,
    output SB_T3_SOUTH_SB_OUT_B17_valid,
    input SB_T3_SOUTH_SB_OUT_B1_ready,
    output SB_T3_SOUTH_SB_OUT_B1_valid,
    input [0:0] SB_T3_WEST_SB_IN_B1,
    input [16:0] SB_T3_WEST_SB_IN_B17,
    output SB_T3_WEST_SB_IN_B17_ready,
    input SB_T3_WEST_SB_IN_B17_valid,
    output SB_T3_WEST_SB_IN_B1_ready,
    input SB_T3_WEST_SB_IN_B1_valid,
    output [0:0] SB_T3_WEST_SB_OUT_B1,
    output [16:0] SB_T3_WEST_SB_OUT_B17,
    input SB_T3_WEST_SB_OUT_B17_ready,
    output SB_T3_WEST_SB_OUT_B17_valid,
    input SB_T3_WEST_SB_OUT_B1_ready,
    output SB_T3_WEST_SB_OUT_B1_valid,
    input [0:0] SB_T4_EAST_SB_IN_B1,
    input [16:0] SB_T4_EAST_SB_IN_B17,
    output SB_T4_EAST_SB_IN_B17_ready,
    input SB_T4_EAST_SB_IN_B17_valid,
    output SB_T4_EAST_SB_IN_B1_ready,
    input SB_T4_EAST_SB_IN_B1_valid,
    output [0:0] SB_T4_EAST_SB_OUT_B1,
    output [16:0] SB_T4_EAST_SB_OUT_B17,
    input SB_T4_EAST_SB_OUT_B17_ready,
    output SB_T4_EAST_SB_OUT_B17_valid,
    input SB_T4_EAST_SB_OUT_B1_ready,
    output SB_T4_EAST_SB_OUT_B1_valid,
    input [0:0] SB_T4_NORTH_SB_IN_B1,
    input [16:0] SB_T4_NORTH_SB_IN_B17,
    output SB_T4_NORTH_SB_IN_B17_ready,
    input SB_T4_NORTH_SB_IN_B17_valid,
    output SB_T4_NORTH_SB_IN_B1_ready,
    input SB_T4_NORTH_SB_IN_B1_valid,
    output [0:0] SB_T4_NORTH_SB_OUT_B1,
    output [16:0] SB_T4_NORTH_SB_OUT_B17,
    input SB_T4_NORTH_SB_OUT_B17_ready,
    output SB_T4_NORTH_SB_OUT_B17_valid,
    input SB_T4_NORTH_SB_OUT_B1_ready,
    output SB_T4_NORTH_SB_OUT_B1_valid,
    input [0:0] SB_T4_SOUTH_SB_IN_B1,
    input [16:0] SB_T4_SOUTH_SB_IN_B17,
    output SB_T4_SOUTH_SB_IN_B17_ready,
    input SB_T4_SOUTH_SB_IN_B17_valid,
    output SB_T4_SOUTH_SB_IN_B1_ready,
    input SB_T4_SOUTH_SB_IN_B1_valid,
    output [0:0] SB_T4_SOUTH_SB_OUT_B1,
    output [16:0] SB_T4_SOUTH_SB_OUT_B17,
    input SB_T4_SOUTH_SB_OUT_B17_ready,
    output SB_T4_SOUTH_SB_OUT_B17_valid,
    input SB_T4_SOUTH_SB_OUT_B1_ready,
    output SB_T4_SOUTH_SB_OUT_B1_valid,
    input [0:0] SB_T4_WEST_SB_IN_B1,
    input [16:0] SB_T4_WEST_SB_IN_B17,
    output SB_T4_WEST_SB_IN_B17_ready,
    input SB_T4_WEST_SB_IN_B17_valid,
    output SB_T4_WEST_SB_IN_B1_ready,
    input SB_T4_WEST_SB_IN_B1_valid,
    output [0:0] SB_T4_WEST_SB_OUT_B1,
    output [16:0] SB_T4_WEST_SB_OUT_B17,
    input SB_T4_WEST_SB_OUT_B17_ready,
    output SB_T4_WEST_SB_OUT_B17_valid,
    input SB_T4_WEST_SB_OUT_B1_ready,
    output SB_T4_WEST_SB_OUT_B1_valid,
    input clk,
    output clk_out,
    input [31:0] config_config_addr,
    input [31:0] config_config_data,
    output [31:0] config_out_config_addr,
    output [31:0] config_out_config_data,
    output [0:0] config_out_read,
    output [0:0] config_out_write,
    input [0:0] config_read,
    input [0:0] config_write,
    input [0:0] flush,
    output [0:0] flush_out,
    output [8:0] hi,
    output [7:0] lo,
    output [31:0] read_config_data,
    input [31:0] read_config_data_in,
    input reset,
    output reset_out,
    input [0:0] stall,
    output [0:0] stall_out,
    input [15:0] tile_id
);
wire [16:0] CB_MEM_input_width_17_num_0_O;
wire CB_MEM_input_width_17_num_0_enable;
wire [31:0] CB_MEM_input_width_17_num_0_out_sel;
wire [31:0] CB_MEM_input_width_17_num_0_read_config_data;
wire CB_MEM_input_width_17_num_0_ready_out;
wire CB_MEM_input_width_17_num_0_valid_out;
wire [16:0] CB_MEM_input_width_17_num_1_O;
wire CB_MEM_input_width_17_num_1_enable;
wire [31:0] CB_MEM_input_width_17_num_1_out_sel;
wire [31:0] CB_MEM_input_width_17_num_1_read_config_data;
wire CB_MEM_input_width_17_num_1_ready_out;
wire CB_MEM_input_width_17_num_1_valid_out;
wire [16:0] CB_MEM_input_width_17_num_2_O;
wire CB_MEM_input_width_17_num_2_enable;
wire [31:0] CB_MEM_input_width_17_num_2_out_sel;
wire [31:0] CB_MEM_input_width_17_num_2_read_config_data;
wire CB_MEM_input_width_17_num_2_ready_out;
wire CB_MEM_input_width_17_num_2_valid_out;
wire [16:0] CB_MEM_input_width_17_num_3_O;
wire CB_MEM_input_width_17_num_3_enable;
wire [31:0] CB_MEM_input_width_17_num_3_out_sel;
wire [31:0] CB_MEM_input_width_17_num_3_read_config_data;
wire CB_MEM_input_width_17_num_3_ready_out;
wire CB_MEM_input_width_17_num_3_valid_out;
wire [0:0] CB_MEM_input_width_1_num_0_O;
wire CB_MEM_input_width_1_num_0_enable;
wire [31:0] CB_MEM_input_width_1_num_0_out_sel;
wire [31:0] CB_MEM_input_width_1_num_0_read_config_data;
wire CB_MEM_input_width_1_num_0_ready_out;
wire CB_MEM_input_width_1_num_0_valid_out;
wire [0:0] CB_MEM_input_width_1_num_1_O;
wire CB_MEM_input_width_1_num_1_enable;
wire [31:0] CB_MEM_input_width_1_num_1_out_sel;
wire [31:0] CB_MEM_input_width_1_num_1_read_config_data;
wire CB_MEM_input_width_1_num_1_ready_out;
wire CB_MEM_input_width_1_num_1_valid_out;
wire [0:0] CB_flush_O;
wire CB_flush_enable;
wire [31:0] CB_flush_out_sel;
wire [31:0] CB_flush_read_config_data;
wire CB_flush_ready_out;
wire CB_flush_valid_out;
wire DECODE_FEATURE_0_O;
wire DECODE_FEATURE_1_O;
wire DECODE_FEATURE_10_O;
wire DECODE_FEATURE_11_O;
wire DECODE_FEATURE_12_O;
wire DECODE_FEATURE_2_O;
wire DECODE_FEATURE_3_O;
wire DECODE_FEATURE_4_O;
wire DECODE_FEATURE_5_O;
wire DECODE_FEATURE_6_O;
wire DECODE_FEATURE_7_O;
wire DECODE_FEATURE_8_O;
wire DECODE_FEATURE_9_O;
wire FEATURE_AND_0_out;
wire FEATURE_AND_1_out;
wire FEATURE_AND_10_out;
wire FEATURE_AND_11_out;
wire FEATURE_AND_12_out;
wire FEATURE_AND_2_out;
wire FEATURE_AND_3_out;
wire FEATURE_AND_4_out;
wire FEATURE_AND_5_out;
wire FEATURE_AND_6_out;
wire FEATURE_AND_7_out;
wire FEATURE_AND_8_out;
wire FEATURE_AND_9_out;
wire [0:0] MEM_output_width_17_num_0_loopback_valid_out;
wire [0:0] MEM_output_width_17_num_1_loopback_valid_out;
wire [0:0] MEM_output_width_17_num_2_loopback_valid_out;
wire [0:0] MEM_output_width_1_num_0_loopback_valid_out;
wire [0:0] MEM_output_width_1_num_1_loopback_valid_out;
wire [0:0] MEM_output_width_1_num_2_loopback_valid_out;
wire [0:0] MemCore_inst0_MEM_input_width_17_num_0_ready;
wire [0:0] MemCore_inst0_MEM_input_width_17_num_1_ready;
wire [0:0] MemCore_inst0_MEM_input_width_17_num_2_ready;
wire [0:0] MemCore_inst0_MEM_input_width_17_num_3_ready;
wire MemCore_inst0_MEM_input_width_1_num_0_ready;
wire MemCore_inst0_MEM_input_width_1_num_1_ready;
wire [16:0] MemCore_inst0_MEM_output_width_17_num_0;
wire [0:0] MemCore_inst0_MEM_output_width_17_num_0_valid;
wire [16:0] MemCore_inst0_MEM_output_width_17_num_1;
wire [0:0] MemCore_inst0_MEM_output_width_17_num_1_valid;
wire [16:0] MemCore_inst0_MEM_output_width_17_num_2;
wire [0:0] MemCore_inst0_MEM_output_width_17_num_2_valid;
wire [0:0] MemCore_inst0_MEM_output_width_1_num_0;
wire MemCore_inst0_MEM_output_width_1_num_0_valid;
wire [0:0] MemCore_inst0_MEM_output_width_1_num_1;
wire MemCore_inst0_MEM_output_width_1_num_1_valid;
wire [0:0] MemCore_inst0_MEM_output_width_1_num_2;
wire MemCore_inst0_MEM_output_width_1_num_2_valid;
wire [31:0] MemCore_inst0_read_config_data;
wire [31:0] MemCore_inst0_read_config_data_1;
wire [31:0] MemCore_inst0_read_config_data_2;
wire [0:0] PowerDomainConfigReg_inst0_ps_en_out;
wire [31:0] PowerDomainConfigReg_inst0_read_config_data;
wire [31:0] PowerDomainOR_O;
wire SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_0_ready_out;
wire SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_1_ready_out;
wire SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_2_ready_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_OUT_B17_valid_out;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_IN_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_IN_B17_ready_out;
wire [16:0] SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_OUT_B17;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_OUT_B17_enable;
wire SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_OUT_B17_valid_out;
wire [31:0] SB_ID0_5TRACKS_B17_MemCore_read_config_data;
wire SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_0_ready_out;
wire SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_1_ready_out;
wire SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_2_ready_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1_valid_out;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_IN_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_IN_B1_ready_out;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1_enable;
wire SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1_valid_out;
wire [31:0] SB_ID0_5TRACKS_B1_MemCore_read_config_data;
wire SB_T0_EAST_SB_OUT_B17_ready_and_Z;
wire SB_T0_EAST_SB_OUT_B1_ready_and_Z;
wire SB_T0_NORTH_SB_OUT_B17_ready_and_Z;
wire SB_T0_NORTH_SB_OUT_B1_ready_and_Z;
wire SB_T0_SOUTH_SB_OUT_B17_ready_and_Z;
wire SB_T0_SOUTH_SB_OUT_B1_ready_and_Z;
wire SB_T0_WEST_SB_OUT_B17_ready_and_Z;
wire SB_T0_WEST_SB_OUT_B1_ready_and_Z;
wire SB_T1_EAST_SB_OUT_B17_ready_and_Z;
wire SB_T1_EAST_SB_OUT_B1_ready_and_Z;
wire SB_T1_NORTH_SB_OUT_B17_ready_and_Z;
wire SB_T1_NORTH_SB_OUT_B1_ready_and_Z;
wire SB_T1_SOUTH_SB_OUT_B17_ready_and_Z;
wire SB_T1_SOUTH_SB_OUT_B1_ready_and_Z;
wire SB_T1_WEST_SB_OUT_B17_ready_and_Z;
wire SB_T1_WEST_SB_OUT_B1_ready_and_Z;
wire SB_T2_EAST_SB_OUT_B17_ready_and_Z;
wire SB_T2_EAST_SB_OUT_B1_ready_and_Z;
wire SB_T2_NORTH_SB_OUT_B17_ready_and_Z;
wire SB_T2_NORTH_SB_OUT_B1_ready_and_Z;
wire SB_T2_SOUTH_SB_OUT_B17_ready_and_Z;
wire SB_T2_SOUTH_SB_OUT_B1_ready_and_Z;
wire SB_T2_WEST_SB_OUT_B17_ready_and_Z;
wire SB_T2_WEST_SB_OUT_B1_ready_and_Z;
wire SB_T3_EAST_SB_OUT_B17_ready_and_Z;
wire SB_T3_EAST_SB_OUT_B1_ready_and_Z;
wire SB_T3_NORTH_SB_OUT_B17_ready_and_Z;
wire SB_T3_NORTH_SB_OUT_B1_ready_and_Z;
wire SB_T3_SOUTH_SB_OUT_B17_ready_and_Z;
wire SB_T3_SOUTH_SB_OUT_B1_ready_and_Z;
wire SB_T3_WEST_SB_OUT_B17_ready_and_Z;
wire SB_T3_WEST_SB_OUT_B1_ready_and_Z;
wire SB_T4_EAST_SB_OUT_B17_ready_and_Z;
wire SB_T4_EAST_SB_OUT_B1_ready_and_Z;
wire SB_T4_NORTH_SB_OUT_B17_ready_and_Z;
wire SB_T4_NORTH_SB_OUT_B1_ready_and_Z;
wire SB_T4_SOUTH_SB_OUT_B17_ready_and_Z;
wire SB_T4_SOUTH_SB_OUT_B1_ready_and_Z;
wire SB_T4_WEST_SB_OUT_B17_ready_and_Z;
wire SB_T4_WEST_SB_OUT_B1_ready_and_Z;
wire and_inst0_out;
wire and_inst1_out;
wire bit_const_1_None_out;
wire [7:0] const_0_8_out;
wire [8:0] const_511_9_out;
wire coreir_eq_16_inst0_out;
wire [31:0] read_data_mux_O;
wire [31:0] self_config_config_addr_out;
wire [16:0] CB_MEM_input_width_17_num_0_I [19:0];
assign CB_MEM_input_width_17_num_0_I[19] = SB_T4_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[18] = SB_T4_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[17] = SB_T4_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[16] = SB_T4_NORTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[15] = SB_T3_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[14] = SB_T3_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[13] = SB_T3_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[12] = SB_T3_NORTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[11] = SB_T2_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[10] = SB_T2_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[9] = SB_T2_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[8] = SB_T2_NORTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[7] = SB_T1_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[6] = SB_T1_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[5] = SB_T1_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[4] = SB_T1_NORTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[3] = SB_T0_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[2] = SB_T0_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[1] = SB_T0_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_0_I[0] = SB_T0_NORTH_SB_IN_B17;
wire [19:0] CB_MEM_input_width_17_num_0_valid_in;
assign CB_MEM_input_width_17_num_0_valid_in = {SB_T4_WEST_SB_IN_B17_valid,SB_T4_EAST_SB_IN_B17_valid,SB_T4_SOUTH_SB_IN_B17_valid,SB_T4_NORTH_SB_IN_B17_valid,SB_T3_WEST_SB_IN_B17_valid,SB_T3_EAST_SB_IN_B17_valid,SB_T3_SOUTH_SB_IN_B17_valid,SB_T3_NORTH_SB_IN_B17_valid,SB_T2_WEST_SB_IN_B17_valid,SB_T2_EAST_SB_IN_B17_valid,SB_T2_SOUTH_SB_IN_B17_valid,SB_T2_NORTH_SB_IN_B17_valid,SB_T1_WEST_SB_IN_B17_valid,SB_T1_EAST_SB_IN_B17_valid,SB_T1_SOUTH_SB_IN_B17_valid,SB_T1_NORTH_SB_IN_B17_valid,SB_T0_WEST_SB_IN_B17_valid,SB_T0_EAST_SB_IN_B17_valid,SB_T0_SOUTH_SB_IN_B17_valid,SB_T0_NORTH_SB_IN_B17_valid};
CB_MEM_input_width_17_num_0 CB_MEM_input_width_17_num_0 (
    .I(CB_MEM_input_width_17_num_0_I),
    .O(CB_MEM_input_width_17_num_0_O),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_3_out),
    .enable(CB_MEM_input_width_17_num_0_enable),
    .out_sel(CB_MEM_input_width_17_num_0_out_sel),
    .read_config_data(CB_MEM_input_width_17_num_0_read_config_data),
    .ready_in(MemCore_inst0_MEM_input_width_17_num_0_ready[0]),
    .ready_out(CB_MEM_input_width_17_num_0_ready_out),
    .reset(reset),
    .valid_in(CB_MEM_input_width_17_num_0_valid_in),
    .valid_out(CB_MEM_input_width_17_num_0_valid_out)
);
wire [16:0] CB_MEM_input_width_17_num_1_I [19:0];
assign CB_MEM_input_width_17_num_1_I[19] = SB_T4_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[18] = SB_T4_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[17] = SB_T4_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[16] = SB_T4_NORTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[15] = SB_T3_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[14] = SB_T3_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[13] = SB_T3_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[12] = SB_T3_NORTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[11] = SB_T2_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[10] = SB_T2_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[9] = SB_T2_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[8] = SB_T2_NORTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[7] = SB_T1_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[6] = SB_T1_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[5] = SB_T1_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[4] = SB_T1_NORTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[3] = SB_T0_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[2] = SB_T0_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[1] = SB_T0_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_1_I[0] = SB_T0_NORTH_SB_IN_B17;
wire [19:0] CB_MEM_input_width_17_num_1_valid_in;
assign CB_MEM_input_width_17_num_1_valid_in = {SB_T4_WEST_SB_IN_B17_valid,SB_T4_EAST_SB_IN_B17_valid,SB_T4_SOUTH_SB_IN_B17_valid,SB_T4_NORTH_SB_IN_B17_valid,SB_T3_WEST_SB_IN_B17_valid,SB_T3_EAST_SB_IN_B17_valid,SB_T3_SOUTH_SB_IN_B17_valid,SB_T3_NORTH_SB_IN_B17_valid,SB_T2_WEST_SB_IN_B17_valid,SB_T2_EAST_SB_IN_B17_valid,SB_T2_SOUTH_SB_IN_B17_valid,SB_T2_NORTH_SB_IN_B17_valid,SB_T1_WEST_SB_IN_B17_valid,SB_T1_EAST_SB_IN_B17_valid,SB_T1_SOUTH_SB_IN_B17_valid,SB_T1_NORTH_SB_IN_B17_valid,SB_T0_WEST_SB_IN_B17_valid,SB_T0_EAST_SB_IN_B17_valid,SB_T0_SOUTH_SB_IN_B17_valid,SB_T0_NORTH_SB_IN_B17_valid};
CB_MEM_input_width_17_num_1 CB_MEM_input_width_17_num_1 (
    .I(CB_MEM_input_width_17_num_1_I),
    .O(CB_MEM_input_width_17_num_1_O),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_4_out),
    .enable(CB_MEM_input_width_17_num_1_enable),
    .out_sel(CB_MEM_input_width_17_num_1_out_sel),
    .read_config_data(CB_MEM_input_width_17_num_1_read_config_data),
    .ready_in(MemCore_inst0_MEM_input_width_17_num_1_ready[0]),
    .ready_out(CB_MEM_input_width_17_num_1_ready_out),
    .reset(reset),
    .valid_in(CB_MEM_input_width_17_num_1_valid_in),
    .valid_out(CB_MEM_input_width_17_num_1_valid_out)
);
wire [16:0] CB_MEM_input_width_17_num_2_I [19:0];
assign CB_MEM_input_width_17_num_2_I[19] = SB_T4_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[18] = SB_T4_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[17] = SB_T4_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[16] = SB_T4_NORTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[15] = SB_T3_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[14] = SB_T3_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[13] = SB_T3_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[12] = SB_T3_NORTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[11] = SB_T2_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[10] = SB_T2_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[9] = SB_T2_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[8] = SB_T2_NORTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[7] = SB_T1_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[6] = SB_T1_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[5] = SB_T1_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[4] = SB_T1_NORTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[3] = SB_T0_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[2] = SB_T0_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[1] = SB_T0_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_2_I[0] = SB_T0_NORTH_SB_IN_B17;
wire [19:0] CB_MEM_input_width_17_num_2_valid_in;
assign CB_MEM_input_width_17_num_2_valid_in = {SB_T4_WEST_SB_IN_B17_valid,SB_T4_EAST_SB_IN_B17_valid,SB_T4_SOUTH_SB_IN_B17_valid,SB_T4_NORTH_SB_IN_B17_valid,SB_T3_WEST_SB_IN_B17_valid,SB_T3_EAST_SB_IN_B17_valid,SB_T3_SOUTH_SB_IN_B17_valid,SB_T3_NORTH_SB_IN_B17_valid,SB_T2_WEST_SB_IN_B17_valid,SB_T2_EAST_SB_IN_B17_valid,SB_T2_SOUTH_SB_IN_B17_valid,SB_T2_NORTH_SB_IN_B17_valid,SB_T1_WEST_SB_IN_B17_valid,SB_T1_EAST_SB_IN_B17_valid,SB_T1_SOUTH_SB_IN_B17_valid,SB_T1_NORTH_SB_IN_B17_valid,SB_T0_WEST_SB_IN_B17_valid,SB_T0_EAST_SB_IN_B17_valid,SB_T0_SOUTH_SB_IN_B17_valid,SB_T0_NORTH_SB_IN_B17_valid};
CB_MEM_input_width_17_num_2 CB_MEM_input_width_17_num_2 (
    .I(CB_MEM_input_width_17_num_2_I),
    .O(CB_MEM_input_width_17_num_2_O),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_5_out),
    .enable(CB_MEM_input_width_17_num_2_enable),
    .out_sel(CB_MEM_input_width_17_num_2_out_sel),
    .read_config_data(CB_MEM_input_width_17_num_2_read_config_data),
    .ready_in(MemCore_inst0_MEM_input_width_17_num_2_ready[0]),
    .ready_out(CB_MEM_input_width_17_num_2_ready_out),
    .reset(reset),
    .valid_in(CB_MEM_input_width_17_num_2_valid_in),
    .valid_out(CB_MEM_input_width_17_num_2_valid_out)
);
wire [16:0] CB_MEM_input_width_17_num_3_I [19:0];
assign CB_MEM_input_width_17_num_3_I[19] = SB_T4_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[18] = SB_T4_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[17] = SB_T4_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[16] = SB_T4_NORTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[15] = SB_T3_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[14] = SB_T3_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[13] = SB_T3_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[12] = SB_T3_NORTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[11] = SB_T2_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[10] = SB_T2_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[9] = SB_T2_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[8] = SB_T2_NORTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[7] = SB_T1_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[6] = SB_T1_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[5] = SB_T1_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[4] = SB_T1_NORTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[3] = SB_T0_WEST_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[2] = SB_T0_EAST_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[1] = SB_T0_SOUTH_SB_IN_B17;
assign CB_MEM_input_width_17_num_3_I[0] = SB_T0_NORTH_SB_IN_B17;
wire [19:0] CB_MEM_input_width_17_num_3_valid_in;
assign CB_MEM_input_width_17_num_3_valid_in = {SB_T4_WEST_SB_IN_B17_valid,SB_T4_EAST_SB_IN_B17_valid,SB_T4_SOUTH_SB_IN_B17_valid,SB_T4_NORTH_SB_IN_B17_valid,SB_T3_WEST_SB_IN_B17_valid,SB_T3_EAST_SB_IN_B17_valid,SB_T3_SOUTH_SB_IN_B17_valid,SB_T3_NORTH_SB_IN_B17_valid,SB_T2_WEST_SB_IN_B17_valid,SB_T2_EAST_SB_IN_B17_valid,SB_T2_SOUTH_SB_IN_B17_valid,SB_T2_NORTH_SB_IN_B17_valid,SB_T1_WEST_SB_IN_B17_valid,SB_T1_EAST_SB_IN_B17_valid,SB_T1_SOUTH_SB_IN_B17_valid,SB_T1_NORTH_SB_IN_B17_valid,SB_T0_WEST_SB_IN_B17_valid,SB_T0_EAST_SB_IN_B17_valid,SB_T0_SOUTH_SB_IN_B17_valid,SB_T0_NORTH_SB_IN_B17_valid};
CB_MEM_input_width_17_num_3 CB_MEM_input_width_17_num_3 (
    .I(CB_MEM_input_width_17_num_3_I),
    .O(CB_MEM_input_width_17_num_3_O),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_6_out),
    .enable(CB_MEM_input_width_17_num_3_enable),
    .out_sel(CB_MEM_input_width_17_num_3_out_sel),
    .read_config_data(CB_MEM_input_width_17_num_3_read_config_data),
    .ready_in(MemCore_inst0_MEM_input_width_17_num_3_ready[0]),
    .ready_out(CB_MEM_input_width_17_num_3_ready_out),
    .reset(reset),
    .valid_in(CB_MEM_input_width_17_num_3_valid_in),
    .valid_out(CB_MEM_input_width_17_num_3_valid_out)
);
wire [0:0] CB_MEM_input_width_1_num_0_I [19:0];
assign CB_MEM_input_width_1_num_0_I[19] = SB_T4_WEST_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[18] = SB_T4_EAST_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[17] = SB_T4_SOUTH_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[16] = SB_T4_NORTH_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[15] = SB_T3_WEST_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[14] = SB_T3_EAST_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[13] = SB_T3_SOUTH_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[12] = SB_T3_NORTH_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[11] = SB_T2_WEST_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[10] = SB_T2_EAST_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[9] = SB_T2_SOUTH_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[8] = SB_T2_NORTH_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[7] = SB_T1_WEST_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[6] = SB_T1_EAST_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[5] = SB_T1_SOUTH_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[4] = SB_T1_NORTH_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[3] = SB_T0_WEST_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[2] = SB_T0_EAST_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[1] = SB_T0_SOUTH_SB_IN_B1;
assign CB_MEM_input_width_1_num_0_I[0] = SB_T0_NORTH_SB_IN_B1;
wire [19:0] CB_MEM_input_width_1_num_0_valid_in;
assign CB_MEM_input_width_1_num_0_valid_in = {SB_T4_WEST_SB_IN_B1_valid,SB_T4_EAST_SB_IN_B1_valid,SB_T4_SOUTH_SB_IN_B1_valid,SB_T4_NORTH_SB_IN_B1_valid,SB_T3_WEST_SB_IN_B1_valid,SB_T3_EAST_SB_IN_B1_valid,SB_T3_SOUTH_SB_IN_B1_valid,SB_T3_NORTH_SB_IN_B1_valid,SB_T2_WEST_SB_IN_B1_valid,SB_T2_EAST_SB_IN_B1_valid,SB_T2_SOUTH_SB_IN_B1_valid,SB_T2_NORTH_SB_IN_B1_valid,SB_T1_WEST_SB_IN_B1_valid,SB_T1_EAST_SB_IN_B1_valid,SB_T1_SOUTH_SB_IN_B1_valid,SB_T1_NORTH_SB_IN_B1_valid,SB_T0_WEST_SB_IN_B1_valid,SB_T0_EAST_SB_IN_B1_valid,SB_T0_SOUTH_SB_IN_B1_valid,SB_T0_NORTH_SB_IN_B1_valid};
CB_MEM_input_width_1_num_0 CB_MEM_input_width_1_num_0 (
    .I(CB_MEM_input_width_1_num_0_I),
    .O(CB_MEM_input_width_1_num_0_O),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_7_out),
    .enable(CB_MEM_input_width_1_num_0_enable),
    .out_sel(CB_MEM_input_width_1_num_0_out_sel),
    .read_config_data(CB_MEM_input_width_1_num_0_read_config_data),
    .ready_in(MemCore_inst0_MEM_input_width_1_num_0_ready),
    .ready_out(CB_MEM_input_width_1_num_0_ready_out),
    .reset(reset),
    .valid_in(CB_MEM_input_width_1_num_0_valid_in),
    .valid_out(CB_MEM_input_width_1_num_0_valid_out)
);
wire [0:0] CB_MEM_input_width_1_num_1_I [19:0];
assign CB_MEM_input_width_1_num_1_I[19] = SB_T4_WEST_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[18] = SB_T4_EAST_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[17] = SB_T4_SOUTH_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[16] = SB_T4_NORTH_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[15] = SB_T3_WEST_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[14] = SB_T3_EAST_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[13] = SB_T3_SOUTH_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[12] = SB_T3_NORTH_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[11] = SB_T2_WEST_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[10] = SB_T2_EAST_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[9] = SB_T2_SOUTH_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[8] = SB_T2_NORTH_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[7] = SB_T1_WEST_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[6] = SB_T1_EAST_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[5] = SB_T1_SOUTH_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[4] = SB_T1_NORTH_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[3] = SB_T0_WEST_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[2] = SB_T0_EAST_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[1] = SB_T0_SOUTH_SB_IN_B1;
assign CB_MEM_input_width_1_num_1_I[0] = SB_T0_NORTH_SB_IN_B1;
wire [19:0] CB_MEM_input_width_1_num_1_valid_in;
assign CB_MEM_input_width_1_num_1_valid_in = {SB_T4_WEST_SB_IN_B1_valid,SB_T4_EAST_SB_IN_B1_valid,SB_T4_SOUTH_SB_IN_B1_valid,SB_T4_NORTH_SB_IN_B1_valid,SB_T3_WEST_SB_IN_B1_valid,SB_T3_EAST_SB_IN_B1_valid,SB_T3_SOUTH_SB_IN_B1_valid,SB_T3_NORTH_SB_IN_B1_valid,SB_T2_WEST_SB_IN_B1_valid,SB_T2_EAST_SB_IN_B1_valid,SB_T2_SOUTH_SB_IN_B1_valid,SB_T2_NORTH_SB_IN_B1_valid,SB_T1_WEST_SB_IN_B1_valid,SB_T1_EAST_SB_IN_B1_valid,SB_T1_SOUTH_SB_IN_B1_valid,SB_T1_NORTH_SB_IN_B1_valid,SB_T0_WEST_SB_IN_B1_valid,SB_T0_EAST_SB_IN_B1_valid,SB_T0_SOUTH_SB_IN_B1_valid,SB_T0_NORTH_SB_IN_B1_valid};
CB_MEM_input_width_1_num_1 CB_MEM_input_width_1_num_1 (
    .I(CB_MEM_input_width_1_num_1_I),
    .O(CB_MEM_input_width_1_num_1_O),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_8_out),
    .enable(CB_MEM_input_width_1_num_1_enable),
    .out_sel(CB_MEM_input_width_1_num_1_out_sel),
    .read_config_data(CB_MEM_input_width_1_num_1_read_config_data),
    .ready_in(MemCore_inst0_MEM_input_width_1_num_1_ready),
    .ready_out(CB_MEM_input_width_1_num_1_ready_out),
    .reset(reset),
    .valid_in(CB_MEM_input_width_1_num_1_valid_in),
    .valid_out(CB_MEM_input_width_1_num_1_valid_out)
);
wire [0:0] CB_flush_I [19:0];
assign CB_flush_I[19] = SB_T4_WEST_SB_IN_B1;
assign CB_flush_I[18] = SB_T4_EAST_SB_IN_B1;
assign CB_flush_I[17] = SB_T4_SOUTH_SB_IN_B1;
assign CB_flush_I[16] = SB_T4_NORTH_SB_IN_B1;
assign CB_flush_I[15] = SB_T3_WEST_SB_IN_B1;
assign CB_flush_I[14] = SB_T3_EAST_SB_IN_B1;
assign CB_flush_I[13] = SB_T3_SOUTH_SB_IN_B1;
assign CB_flush_I[12] = SB_T3_NORTH_SB_IN_B1;
assign CB_flush_I[11] = SB_T2_WEST_SB_IN_B1;
assign CB_flush_I[10] = SB_T2_EAST_SB_IN_B1;
assign CB_flush_I[9] = SB_T2_SOUTH_SB_IN_B1;
assign CB_flush_I[8] = SB_T2_NORTH_SB_IN_B1;
assign CB_flush_I[7] = SB_T1_WEST_SB_IN_B1;
assign CB_flush_I[6] = SB_T1_EAST_SB_IN_B1;
assign CB_flush_I[5] = SB_T1_SOUTH_SB_IN_B1;
assign CB_flush_I[4] = SB_T1_NORTH_SB_IN_B1;
assign CB_flush_I[3] = SB_T0_WEST_SB_IN_B1;
assign CB_flush_I[2] = SB_T0_EAST_SB_IN_B1;
assign CB_flush_I[1] = SB_T0_SOUTH_SB_IN_B1;
assign CB_flush_I[0] = SB_T0_NORTH_SB_IN_B1;
wire [19:0] CB_flush_valid_in;
assign CB_flush_valid_in = {SB_T4_WEST_SB_IN_B1_valid,SB_T4_EAST_SB_IN_B1_valid,SB_T4_SOUTH_SB_IN_B1_valid,SB_T4_NORTH_SB_IN_B1_valid,SB_T3_WEST_SB_IN_B1_valid,SB_T3_EAST_SB_IN_B1_valid,SB_T3_SOUTH_SB_IN_B1_valid,SB_T3_NORTH_SB_IN_B1_valid,SB_T2_WEST_SB_IN_B1_valid,SB_T2_EAST_SB_IN_B1_valid,SB_T2_SOUTH_SB_IN_B1_valid,SB_T2_NORTH_SB_IN_B1_valid,SB_T1_WEST_SB_IN_B1_valid,SB_T1_EAST_SB_IN_B1_valid,SB_T1_SOUTH_SB_IN_B1_valid,SB_T1_NORTH_SB_IN_B1_valid,SB_T0_WEST_SB_IN_B1_valid,SB_T0_EAST_SB_IN_B1_valid,SB_T0_SOUTH_SB_IN_B1_valid,SB_T0_NORTH_SB_IN_B1_valid};
CB_flush CB_flush (
    .I(CB_flush_I),
    .O(CB_flush_O),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_9_out),
    .enable(CB_flush_enable),
    .out_sel(CB_flush_out_sel),
    .read_config_data(CB_flush_read_config_data),
    .ready_in(bit_const_1_None_out),
    .ready_out(CB_flush_ready_out),
    .reset(reset),
    .valid_in(CB_flush_valid_in),
    .valid_out(CB_flush_valid_out)
);
Decode08 DECODE_FEATURE_0 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_0_O)
);
Decode18 DECODE_FEATURE_1 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_1_O)
);
Decode108 DECODE_FEATURE_10 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_10_O)
);
Decode118 DECODE_FEATURE_11 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_11_O)
);
Decode128 DECODE_FEATURE_12 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_12_O)
);
Decode28 DECODE_FEATURE_2 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_2_O)
);
Decode38 DECODE_FEATURE_3 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_3_O)
);
Decode48 DECODE_FEATURE_4 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_4_O)
);
Decode58 DECODE_FEATURE_5 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_5_O)
);
Decode68 DECODE_FEATURE_6 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_6_O)
);
Decode78 DECODE_FEATURE_7 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_7_O)
);
Decode88 DECODE_FEATURE_8 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_8_O)
);
Decode98 DECODE_FEATURE_9 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_9_O)
);
corebit_and FEATURE_AND_0 (
    .in0(DECODE_FEATURE_0_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_0_out)
);
corebit_and FEATURE_AND_1 (
    .in0(DECODE_FEATURE_1_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_1_out)
);
corebit_and FEATURE_AND_10 (
    .in0(DECODE_FEATURE_10_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_10_out)
);
corebit_and FEATURE_AND_11 (
    .in0(DECODE_FEATURE_11_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_11_out)
);
corebit_and FEATURE_AND_12 (
    .in0(DECODE_FEATURE_12_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_12_out)
);
corebit_and FEATURE_AND_2 (
    .in0(DECODE_FEATURE_2_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_2_out)
);
corebit_and FEATURE_AND_3 (
    .in0(DECODE_FEATURE_3_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_3_out)
);
corebit_and FEATURE_AND_4 (
    .in0(DECODE_FEATURE_4_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_4_out)
);
corebit_and FEATURE_AND_5 (
    .in0(DECODE_FEATURE_5_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_5_out)
);
corebit_and FEATURE_AND_6 (
    .in0(DECODE_FEATURE_6_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_6_out)
);
corebit_and FEATURE_AND_7 (
    .in0(DECODE_FEATURE_7_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_7_out)
);
corebit_and FEATURE_AND_8 (
    .in0(DECODE_FEATURE_8_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_8_out)
);
corebit_and FEATURE_AND_9 (
    .in0(DECODE_FEATURE_9_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_9_out)
);
ReadyValidLoopBack MEM_output_width_17_num_0_loopback (
    .ready_in(SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_0_ready_out),
    .valid_in(MemCore_inst0_MEM_output_width_17_num_0_valid),
    .valid_out(MEM_output_width_17_num_0_loopback_valid_out)
);
ReadyValidLoopBack MEM_output_width_17_num_1_loopback (
    .ready_in(SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_1_ready_out),
    .valid_in(MemCore_inst0_MEM_output_width_17_num_1_valid),
    .valid_out(MEM_output_width_17_num_1_loopback_valid_out)
);
ReadyValidLoopBack MEM_output_width_17_num_2_loopback (
    .ready_in(SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_2_ready_out),
    .valid_in(MemCore_inst0_MEM_output_width_17_num_2_valid),
    .valid_out(MEM_output_width_17_num_2_loopback_valid_out)
);
ReadyValidLoopBack MEM_output_width_1_num_0_loopback (
    .ready_in(SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_0_ready_out),
    .valid_in(MemCore_inst0_MEM_output_width_1_num_0_valid),
    .valid_out(MEM_output_width_1_num_0_loopback_valid_out)
);
ReadyValidLoopBack MEM_output_width_1_num_1_loopback (
    .ready_in(SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_1_ready_out),
    .valid_in(MemCore_inst0_MEM_output_width_1_num_1_valid),
    .valid_out(MEM_output_width_1_num_1_loopback_valid_out)
);
ReadyValidLoopBack MEM_output_width_1_num_2_loopback (
    .ready_in(SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_2_ready_out),
    .valid_in(MemCore_inst0_MEM_output_width_1_num_2_valid),
    .valid_out(MEM_output_width_1_num_2_loopback_valid_out)
);
MemCore MemCore_inst0 (
    .MEM_input_width_17_num_0(CB_MEM_input_width_17_num_0_O),
    .MEM_input_width_17_num_0_ready(MemCore_inst0_MEM_input_width_17_num_0_ready),
    .MEM_input_width_17_num_0_valid(CB_MEM_input_width_17_num_0_valid_out),
    .MEM_input_width_17_num_1(CB_MEM_input_width_17_num_1_O),
    .MEM_input_width_17_num_1_ready(MemCore_inst0_MEM_input_width_17_num_1_ready),
    .MEM_input_width_17_num_1_valid(CB_MEM_input_width_17_num_1_valid_out),
    .MEM_input_width_17_num_2(CB_MEM_input_width_17_num_2_O),
    .MEM_input_width_17_num_2_ready(MemCore_inst0_MEM_input_width_17_num_2_ready),
    .MEM_input_width_17_num_2_valid(CB_MEM_input_width_17_num_2_valid_out),
    .MEM_input_width_17_num_3(CB_MEM_input_width_17_num_3_O),
    .MEM_input_width_17_num_3_ready(MemCore_inst0_MEM_input_width_17_num_3_ready),
    .MEM_input_width_17_num_3_valid(CB_MEM_input_width_17_num_3_valid_out),
    .MEM_input_width_1_num_0(CB_MEM_input_width_1_num_0_O),
    .MEM_input_width_1_num_0_ready(MemCore_inst0_MEM_input_width_1_num_0_ready),
    .MEM_input_width_1_num_0_valid(CB_MEM_input_width_1_num_0_valid_out),
    .MEM_input_width_1_num_1(CB_MEM_input_width_1_num_1_O),
    .MEM_input_width_1_num_1_ready(MemCore_inst0_MEM_input_width_1_num_1_ready),
    .MEM_input_width_1_num_1_valid(CB_MEM_input_width_1_num_1_valid_out),
    .MEM_output_width_17_num_0(MemCore_inst0_MEM_output_width_17_num_0),
    .MEM_output_width_17_num_0_ready(SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_0_ready_out),
    .MEM_output_width_17_num_0_valid(MemCore_inst0_MEM_output_width_17_num_0_valid),
    .MEM_output_width_17_num_1(MemCore_inst0_MEM_output_width_17_num_1),
    .MEM_output_width_17_num_1_ready(SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_1_ready_out),
    .MEM_output_width_17_num_1_valid(MemCore_inst0_MEM_output_width_17_num_1_valid),
    .MEM_output_width_17_num_2(MemCore_inst0_MEM_output_width_17_num_2),
    .MEM_output_width_17_num_2_ready(SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_2_ready_out),
    .MEM_output_width_17_num_2_valid(MemCore_inst0_MEM_output_width_17_num_2_valid),
    .MEM_output_width_1_num_0(MemCore_inst0_MEM_output_width_1_num_0),
    .MEM_output_width_1_num_0_ready(SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_0_ready_out),
    .MEM_output_width_1_num_0_valid(MemCore_inst0_MEM_output_width_1_num_0_valid),
    .MEM_output_width_1_num_1(MemCore_inst0_MEM_output_width_1_num_1),
    .MEM_output_width_1_num_1_ready(SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_1_ready_out),
    .MEM_output_width_1_num_1_valid(MemCore_inst0_MEM_output_width_1_num_1_valid),
    .MEM_output_width_1_num_2(MemCore_inst0_MEM_output_width_1_num_2),
    .MEM_output_width_1_num_2_ready(SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_2_ready_out),
    .MEM_output_width_1_num_2_valid(MemCore_inst0_MEM_output_width_1_num_2_valid),
    .clk(clk),
    .config_1_config_addr(self_config_config_addr_out[31:24]),
    .config_1_config_data(config_config_data),
    .config_1_read(config_read),
    .config_1_write(FEATURE_AND_1_out),
    .config_2_config_addr(self_config_config_addr_out[31:24]),
    .config_2_config_data(config_config_data),
    .config_2_read(config_read),
    .config_2_write(FEATURE_AND_2_out),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_en_0(DECODE_FEATURE_1_O),
    .config_en_1(DECODE_FEATURE_2_O),
    .config_read(config_read),
    .config_write(FEATURE_AND_0_out),
    .flush(CB_flush_O),
    .flush_core(flush),
    .read_config_data(MemCore_inst0_read_config_data),
    .read_config_data_1(MemCore_inst0_read_config_data_1),
    .read_config_data_2(MemCore_inst0_read_config_data_2),
    .reset(reset),
    .stall(stall)
);
PowerDomainConfigReg PowerDomainConfigReg_inst0 (
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_12_out),
    .ps_en_out(PowerDomainConfigReg_inst0_ps_en_out),
    .read_config_data(PowerDomainConfigReg_inst0_read_config_data),
    .reset(reset)
);
PowerDomainOR PowerDomainOR (
    .I0(read_data_mux_O),
    .I1(read_config_data_in),
    .O(PowerDomainOR_O),
    .I_not(PowerDomainConfigReg_inst0_ps_en_out)
);
SB_ID0_5TRACKS_B17_MemCore SB_ID0_5TRACKS_B17_MemCore (
    .MEM_input_width_17_num_0_enable(CB_MEM_input_width_17_num_0_enable),
    .MEM_input_width_17_num_0_out_sel(CB_MEM_input_width_17_num_0_out_sel),
    .MEM_input_width_17_num_0_ready(CB_MEM_input_width_17_num_0_ready_out),
    .MEM_input_width_17_num_1_enable(CB_MEM_input_width_17_num_1_enable),
    .MEM_input_width_17_num_1_out_sel(CB_MEM_input_width_17_num_1_out_sel),
    .MEM_input_width_17_num_1_ready(CB_MEM_input_width_17_num_1_ready_out),
    .MEM_input_width_17_num_2_enable(CB_MEM_input_width_17_num_2_enable),
    .MEM_input_width_17_num_2_out_sel(CB_MEM_input_width_17_num_2_out_sel),
    .MEM_input_width_17_num_2_ready(CB_MEM_input_width_17_num_2_ready_out),
    .MEM_input_width_17_num_3_enable(CB_MEM_input_width_17_num_3_enable),
    .MEM_input_width_17_num_3_out_sel(CB_MEM_input_width_17_num_3_out_sel),
    .MEM_input_width_17_num_3_ready(CB_MEM_input_width_17_num_3_ready_out),
    .MEM_output_width_17_num_0(MemCore_inst0_MEM_output_width_17_num_0),
    .MEM_output_width_17_num_0_ready_out(SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_0_ready_out),
    .MEM_output_width_17_num_0_valid(MEM_output_width_17_num_0_loopback_valid_out[0]),
    .MEM_output_width_17_num_1(MemCore_inst0_MEM_output_width_17_num_1),
    .MEM_output_width_17_num_1_ready_out(SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_1_ready_out),
    .MEM_output_width_17_num_1_valid(MEM_output_width_17_num_1_loopback_valid_out[0]),
    .MEM_output_width_17_num_2(MemCore_inst0_MEM_output_width_17_num_2),
    .MEM_output_width_17_num_2_ready_out(SB_ID0_5TRACKS_B17_MemCore_MEM_output_width_17_num_2_ready_out),
    .MEM_output_width_17_num_2_valid(MEM_output_width_17_num_2_loopback_valid_out[0]),
    .SB_T0_EAST_SB_IN_B17(SB_T0_EAST_SB_IN_B17),
    .SB_T0_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_IN_B17_enable),
    .SB_T0_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_IN_B17_ready_out),
    .SB_T0_EAST_SB_IN_B17_valid_in(SB_T0_EAST_SB_IN_B17_valid),
    .SB_T0_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_OUT_B17_enable),
    .SB_T0_EAST_SB_OUT_B17_ready_in(SB_T0_EAST_SB_OUT_B17_ready_and_Z),
    .SB_T0_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_OUT_B17_valid_out),
    .SB_T0_NORTH_SB_IN_B17(SB_T0_NORTH_SB_IN_B17),
    .SB_T0_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_IN_B17_enable),
    .SB_T0_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_IN_B17_ready_out),
    .SB_T0_NORTH_SB_IN_B17_valid_in(SB_T0_NORTH_SB_IN_B17_valid),
    .SB_T0_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_OUT_B17_enable),
    .SB_T0_NORTH_SB_OUT_B17_ready_in(SB_T0_NORTH_SB_OUT_B17_ready_and_Z),
    .SB_T0_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_OUT_B17_valid_out),
    .SB_T0_SOUTH_SB_IN_B17(SB_T0_SOUTH_SB_IN_B17),
    .SB_T0_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_IN_B17_enable),
    .SB_T0_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_IN_B17_ready_out),
    .SB_T0_SOUTH_SB_IN_B17_valid_in(SB_T0_SOUTH_SB_IN_B17_valid),
    .SB_T0_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_OUT_B17_enable),
    .SB_T0_SOUTH_SB_OUT_B17_ready_in(SB_T0_SOUTH_SB_OUT_B17_ready_and_Z),
    .SB_T0_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_OUT_B17_valid_out),
    .SB_T0_WEST_SB_IN_B17(SB_T0_WEST_SB_IN_B17),
    .SB_T0_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_IN_B17_enable),
    .SB_T0_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_IN_B17_ready_out),
    .SB_T0_WEST_SB_IN_B17_valid_in(SB_T0_WEST_SB_IN_B17_valid),
    .SB_T0_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_OUT_B17_enable),
    .SB_T0_WEST_SB_OUT_B17_ready_in(SB_T0_WEST_SB_OUT_B17_ready_and_Z),
    .SB_T0_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_OUT_B17_valid_out),
    .SB_T1_EAST_SB_IN_B17(SB_T1_EAST_SB_IN_B17),
    .SB_T1_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_IN_B17_enable),
    .SB_T1_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_IN_B17_ready_out),
    .SB_T1_EAST_SB_IN_B17_valid_in(SB_T1_EAST_SB_IN_B17_valid),
    .SB_T1_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_OUT_B17_enable),
    .SB_T1_EAST_SB_OUT_B17_ready_in(SB_T1_EAST_SB_OUT_B17_ready_and_Z),
    .SB_T1_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_OUT_B17_valid_out),
    .SB_T1_NORTH_SB_IN_B17(SB_T1_NORTH_SB_IN_B17),
    .SB_T1_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_IN_B17_enable),
    .SB_T1_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_IN_B17_ready_out),
    .SB_T1_NORTH_SB_IN_B17_valid_in(SB_T1_NORTH_SB_IN_B17_valid),
    .SB_T1_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_OUT_B17_enable),
    .SB_T1_NORTH_SB_OUT_B17_ready_in(SB_T1_NORTH_SB_OUT_B17_ready_and_Z),
    .SB_T1_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_OUT_B17_valid_out),
    .SB_T1_SOUTH_SB_IN_B17(SB_T1_SOUTH_SB_IN_B17),
    .SB_T1_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_IN_B17_enable),
    .SB_T1_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_IN_B17_ready_out),
    .SB_T1_SOUTH_SB_IN_B17_valid_in(SB_T1_SOUTH_SB_IN_B17_valid),
    .SB_T1_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_OUT_B17_enable),
    .SB_T1_SOUTH_SB_OUT_B17_ready_in(SB_T1_SOUTH_SB_OUT_B17_ready_and_Z),
    .SB_T1_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_OUT_B17_valid_out),
    .SB_T1_WEST_SB_IN_B17(SB_T1_WEST_SB_IN_B17),
    .SB_T1_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_IN_B17_enable),
    .SB_T1_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_IN_B17_ready_out),
    .SB_T1_WEST_SB_IN_B17_valid_in(SB_T1_WEST_SB_IN_B17_valid),
    .SB_T1_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_OUT_B17_enable),
    .SB_T1_WEST_SB_OUT_B17_ready_in(SB_T1_WEST_SB_OUT_B17_ready_and_Z),
    .SB_T1_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_OUT_B17_valid_out),
    .SB_T2_EAST_SB_IN_B17(SB_T2_EAST_SB_IN_B17),
    .SB_T2_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_IN_B17_enable),
    .SB_T2_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_IN_B17_ready_out),
    .SB_T2_EAST_SB_IN_B17_valid_in(SB_T2_EAST_SB_IN_B17_valid),
    .SB_T2_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_OUT_B17_enable),
    .SB_T2_EAST_SB_OUT_B17_ready_in(SB_T2_EAST_SB_OUT_B17_ready_and_Z),
    .SB_T2_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_OUT_B17_valid_out),
    .SB_T2_NORTH_SB_IN_B17(SB_T2_NORTH_SB_IN_B17),
    .SB_T2_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_IN_B17_enable),
    .SB_T2_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_IN_B17_ready_out),
    .SB_T2_NORTH_SB_IN_B17_valid_in(SB_T2_NORTH_SB_IN_B17_valid),
    .SB_T2_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_OUT_B17_enable),
    .SB_T2_NORTH_SB_OUT_B17_ready_in(SB_T2_NORTH_SB_OUT_B17_ready_and_Z),
    .SB_T2_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_OUT_B17_valid_out),
    .SB_T2_SOUTH_SB_IN_B17(SB_T2_SOUTH_SB_IN_B17),
    .SB_T2_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_IN_B17_enable),
    .SB_T2_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_IN_B17_ready_out),
    .SB_T2_SOUTH_SB_IN_B17_valid_in(SB_T2_SOUTH_SB_IN_B17_valid),
    .SB_T2_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_OUT_B17_enable),
    .SB_T2_SOUTH_SB_OUT_B17_ready_in(SB_T2_SOUTH_SB_OUT_B17_ready_and_Z),
    .SB_T2_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_OUT_B17_valid_out),
    .SB_T2_WEST_SB_IN_B17(SB_T2_WEST_SB_IN_B17),
    .SB_T2_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_IN_B17_enable),
    .SB_T2_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_IN_B17_ready_out),
    .SB_T2_WEST_SB_IN_B17_valid_in(SB_T2_WEST_SB_IN_B17_valid),
    .SB_T2_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_OUT_B17_enable),
    .SB_T2_WEST_SB_OUT_B17_ready_in(SB_T2_WEST_SB_OUT_B17_ready_and_Z),
    .SB_T2_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_OUT_B17_valid_out),
    .SB_T3_EAST_SB_IN_B17(SB_T3_EAST_SB_IN_B17),
    .SB_T3_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_IN_B17_enable),
    .SB_T3_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_IN_B17_ready_out),
    .SB_T3_EAST_SB_IN_B17_valid_in(SB_T3_EAST_SB_IN_B17_valid),
    .SB_T3_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_OUT_B17_enable),
    .SB_T3_EAST_SB_OUT_B17_ready_in(SB_T3_EAST_SB_OUT_B17_ready_and_Z),
    .SB_T3_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_OUT_B17_valid_out),
    .SB_T3_NORTH_SB_IN_B17(SB_T3_NORTH_SB_IN_B17),
    .SB_T3_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_IN_B17_enable),
    .SB_T3_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_IN_B17_ready_out),
    .SB_T3_NORTH_SB_IN_B17_valid_in(SB_T3_NORTH_SB_IN_B17_valid),
    .SB_T3_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_OUT_B17_enable),
    .SB_T3_NORTH_SB_OUT_B17_ready_in(SB_T3_NORTH_SB_OUT_B17_ready_and_Z),
    .SB_T3_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_OUT_B17_valid_out),
    .SB_T3_SOUTH_SB_IN_B17(SB_T3_SOUTH_SB_IN_B17),
    .SB_T3_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_IN_B17_enable),
    .SB_T3_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_IN_B17_ready_out),
    .SB_T3_SOUTH_SB_IN_B17_valid_in(SB_T3_SOUTH_SB_IN_B17_valid),
    .SB_T3_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_OUT_B17_enable),
    .SB_T3_SOUTH_SB_OUT_B17_ready_in(SB_T3_SOUTH_SB_OUT_B17_ready_and_Z),
    .SB_T3_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_OUT_B17_valid_out),
    .SB_T3_WEST_SB_IN_B17(SB_T3_WEST_SB_IN_B17),
    .SB_T3_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_IN_B17_enable),
    .SB_T3_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_IN_B17_ready_out),
    .SB_T3_WEST_SB_IN_B17_valid_in(SB_T3_WEST_SB_IN_B17_valid),
    .SB_T3_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_OUT_B17_enable),
    .SB_T3_WEST_SB_OUT_B17_ready_in(SB_T3_WEST_SB_OUT_B17_ready_and_Z),
    .SB_T3_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_OUT_B17_valid_out),
    .SB_T4_EAST_SB_IN_B17(SB_T4_EAST_SB_IN_B17),
    .SB_T4_EAST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_IN_B17_enable),
    .SB_T4_EAST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_IN_B17_ready_out),
    .SB_T4_EAST_SB_IN_B17_valid_in(SB_T4_EAST_SB_IN_B17_valid),
    .SB_T4_EAST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_EAST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_OUT_B17_enable),
    .SB_T4_EAST_SB_OUT_B17_ready_in(SB_T4_EAST_SB_OUT_B17_ready_and_Z),
    .SB_T4_EAST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_OUT_B17_valid_out),
    .SB_T4_NORTH_SB_IN_B17(SB_T4_NORTH_SB_IN_B17),
    .SB_T4_NORTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_IN_B17_enable),
    .SB_T4_NORTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_IN_B17_ready_out),
    .SB_T4_NORTH_SB_IN_B17_valid_in(SB_T4_NORTH_SB_IN_B17_valid),
    .SB_T4_NORTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_OUT_B17_enable),
    .SB_T4_NORTH_SB_OUT_B17_ready_in(SB_T4_NORTH_SB_OUT_B17_ready_and_Z),
    .SB_T4_NORTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_OUT_B17_valid_out),
    .SB_T4_SOUTH_SB_IN_B17(SB_T4_SOUTH_SB_IN_B17),
    .SB_T4_SOUTH_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_IN_B17_enable),
    .SB_T4_SOUTH_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_IN_B17_ready_out),
    .SB_T4_SOUTH_SB_IN_B17_valid_in(SB_T4_SOUTH_SB_IN_B17_valid),
    .SB_T4_SOUTH_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_OUT_B17_enable),
    .SB_T4_SOUTH_SB_OUT_B17_ready_in(SB_T4_SOUTH_SB_OUT_B17_ready_and_Z),
    .SB_T4_SOUTH_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_OUT_B17_valid_out),
    .SB_T4_WEST_SB_IN_B17(SB_T4_WEST_SB_IN_B17),
    .SB_T4_WEST_SB_IN_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_IN_B17_enable),
    .SB_T4_WEST_SB_IN_B17_ready_out(SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_IN_B17_ready_out),
    .SB_T4_WEST_SB_IN_B17_valid_in(SB_T4_WEST_SB_IN_B17_valid),
    .SB_T4_WEST_SB_OUT_B17(SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_WEST_SB_OUT_B17_enable(SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_OUT_B17_enable),
    .SB_T4_WEST_SB_OUT_B17_ready_in(SB_T4_WEST_SB_OUT_B17_ready_and_Z),
    .SB_T4_WEST_SB_OUT_B17_valid_out(SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_OUT_B17_valid_out),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_11_out),
    .read_config_data(SB_ID0_5TRACKS_B17_MemCore_read_config_data),
    .reset(reset),
    .stall(stall)
);
SB_ID0_5TRACKS_B1_MemCore SB_ID0_5TRACKS_B1_MemCore (
    .MEM_input_width_1_num_0_enable(CB_MEM_input_width_1_num_0_enable),
    .MEM_input_width_1_num_0_out_sel(CB_MEM_input_width_1_num_0_out_sel),
    .MEM_input_width_1_num_0_ready(CB_MEM_input_width_1_num_0_ready_out),
    .MEM_input_width_1_num_1_enable(CB_MEM_input_width_1_num_1_enable),
    .MEM_input_width_1_num_1_out_sel(CB_MEM_input_width_1_num_1_out_sel),
    .MEM_input_width_1_num_1_ready(CB_MEM_input_width_1_num_1_ready_out),
    .MEM_output_width_1_num_0(MemCore_inst0_MEM_output_width_1_num_0),
    .MEM_output_width_1_num_0_ready_out(SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_0_ready_out),
    .MEM_output_width_1_num_0_valid(MEM_output_width_1_num_0_loopback_valid_out[0]),
    .MEM_output_width_1_num_1(MemCore_inst0_MEM_output_width_1_num_1),
    .MEM_output_width_1_num_1_ready_out(SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_1_ready_out),
    .MEM_output_width_1_num_1_valid(MEM_output_width_1_num_1_loopback_valid_out[0]),
    .MEM_output_width_1_num_2(MemCore_inst0_MEM_output_width_1_num_2),
    .MEM_output_width_1_num_2_ready_out(SB_ID0_5TRACKS_B1_MemCore_MEM_output_width_1_num_2_ready_out),
    .MEM_output_width_1_num_2_valid(MEM_output_width_1_num_2_loopback_valid_out[0]),
    .SB_T0_EAST_SB_IN_B1(SB_T0_EAST_SB_IN_B1),
    .SB_T0_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_IN_B1_enable),
    .SB_T0_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_IN_B1_ready_out),
    .SB_T0_EAST_SB_IN_B1_valid_in(SB_T0_EAST_SB_IN_B1_valid),
    .SB_T0_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1_enable),
    .SB_T0_EAST_SB_OUT_B1_ready_in(SB_T0_EAST_SB_OUT_B1_ready_and_Z),
    .SB_T0_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1_valid_out),
    .SB_T0_NORTH_SB_IN_B1(SB_T0_NORTH_SB_IN_B1),
    .SB_T0_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_IN_B1_enable),
    .SB_T0_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_IN_B1_ready_out),
    .SB_T0_NORTH_SB_IN_B1_valid_in(SB_T0_NORTH_SB_IN_B1_valid),
    .SB_T0_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1_enable),
    .SB_T0_NORTH_SB_OUT_B1_ready_in(SB_T0_NORTH_SB_OUT_B1_ready_and_Z),
    .SB_T0_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1_valid_out),
    .SB_T0_SOUTH_SB_IN_B1(SB_T0_SOUTH_SB_IN_B1),
    .SB_T0_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_IN_B1_enable),
    .SB_T0_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_IN_B1_ready_out),
    .SB_T0_SOUTH_SB_IN_B1_valid_in(SB_T0_SOUTH_SB_IN_B1_valid),
    .SB_T0_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1_enable),
    .SB_T0_SOUTH_SB_OUT_B1_ready_in(SB_T0_SOUTH_SB_OUT_B1_ready_and_Z),
    .SB_T0_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1_valid_out),
    .SB_T0_WEST_SB_IN_B1(SB_T0_WEST_SB_IN_B1),
    .SB_T0_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_IN_B1_enable),
    .SB_T0_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_IN_B1_ready_out),
    .SB_T0_WEST_SB_IN_B1_valid_in(SB_T0_WEST_SB_IN_B1_valid),
    .SB_T0_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1_enable),
    .SB_T0_WEST_SB_OUT_B1_ready_in(SB_T0_WEST_SB_OUT_B1_ready_and_Z),
    .SB_T0_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1_valid_out),
    .SB_T1_EAST_SB_IN_B1(SB_T1_EAST_SB_IN_B1),
    .SB_T1_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_IN_B1_enable),
    .SB_T1_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_IN_B1_ready_out),
    .SB_T1_EAST_SB_IN_B1_valid_in(SB_T1_EAST_SB_IN_B1_valid),
    .SB_T1_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1_enable),
    .SB_T1_EAST_SB_OUT_B1_ready_in(SB_T1_EAST_SB_OUT_B1_ready_and_Z),
    .SB_T1_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1_valid_out),
    .SB_T1_NORTH_SB_IN_B1(SB_T1_NORTH_SB_IN_B1),
    .SB_T1_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_IN_B1_enable),
    .SB_T1_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_IN_B1_ready_out),
    .SB_T1_NORTH_SB_IN_B1_valid_in(SB_T1_NORTH_SB_IN_B1_valid),
    .SB_T1_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1_enable),
    .SB_T1_NORTH_SB_OUT_B1_ready_in(SB_T1_NORTH_SB_OUT_B1_ready_and_Z),
    .SB_T1_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1_valid_out),
    .SB_T1_SOUTH_SB_IN_B1(SB_T1_SOUTH_SB_IN_B1),
    .SB_T1_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_IN_B1_enable),
    .SB_T1_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_IN_B1_ready_out),
    .SB_T1_SOUTH_SB_IN_B1_valid_in(SB_T1_SOUTH_SB_IN_B1_valid),
    .SB_T1_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1_enable),
    .SB_T1_SOUTH_SB_OUT_B1_ready_in(SB_T1_SOUTH_SB_OUT_B1_ready_and_Z),
    .SB_T1_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1_valid_out),
    .SB_T1_WEST_SB_IN_B1(SB_T1_WEST_SB_IN_B1),
    .SB_T1_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_IN_B1_enable),
    .SB_T1_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_IN_B1_ready_out),
    .SB_T1_WEST_SB_IN_B1_valid_in(SB_T1_WEST_SB_IN_B1_valid),
    .SB_T1_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1_enable),
    .SB_T1_WEST_SB_OUT_B1_ready_in(SB_T1_WEST_SB_OUT_B1_ready_and_Z),
    .SB_T1_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1_valid_out),
    .SB_T2_EAST_SB_IN_B1(SB_T2_EAST_SB_IN_B1),
    .SB_T2_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_IN_B1_enable),
    .SB_T2_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_IN_B1_ready_out),
    .SB_T2_EAST_SB_IN_B1_valid_in(SB_T2_EAST_SB_IN_B1_valid),
    .SB_T2_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1_enable),
    .SB_T2_EAST_SB_OUT_B1_ready_in(SB_T2_EAST_SB_OUT_B1_ready_and_Z),
    .SB_T2_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1_valid_out),
    .SB_T2_NORTH_SB_IN_B1(SB_T2_NORTH_SB_IN_B1),
    .SB_T2_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_IN_B1_enable),
    .SB_T2_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_IN_B1_ready_out),
    .SB_T2_NORTH_SB_IN_B1_valid_in(SB_T2_NORTH_SB_IN_B1_valid),
    .SB_T2_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1_enable),
    .SB_T2_NORTH_SB_OUT_B1_ready_in(SB_T2_NORTH_SB_OUT_B1_ready_and_Z),
    .SB_T2_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1_valid_out),
    .SB_T2_SOUTH_SB_IN_B1(SB_T2_SOUTH_SB_IN_B1),
    .SB_T2_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_IN_B1_enable),
    .SB_T2_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_IN_B1_ready_out),
    .SB_T2_SOUTH_SB_IN_B1_valid_in(SB_T2_SOUTH_SB_IN_B1_valid),
    .SB_T2_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1_enable),
    .SB_T2_SOUTH_SB_OUT_B1_ready_in(SB_T2_SOUTH_SB_OUT_B1_ready_and_Z),
    .SB_T2_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1_valid_out),
    .SB_T2_WEST_SB_IN_B1(SB_T2_WEST_SB_IN_B1),
    .SB_T2_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_IN_B1_enable),
    .SB_T2_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_IN_B1_ready_out),
    .SB_T2_WEST_SB_IN_B1_valid_in(SB_T2_WEST_SB_IN_B1_valid),
    .SB_T2_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1_enable),
    .SB_T2_WEST_SB_OUT_B1_ready_in(SB_T2_WEST_SB_OUT_B1_ready_and_Z),
    .SB_T2_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1_valid_out),
    .SB_T3_EAST_SB_IN_B1(SB_T3_EAST_SB_IN_B1),
    .SB_T3_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_IN_B1_enable),
    .SB_T3_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_IN_B1_ready_out),
    .SB_T3_EAST_SB_IN_B1_valid_in(SB_T3_EAST_SB_IN_B1_valid),
    .SB_T3_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1_enable),
    .SB_T3_EAST_SB_OUT_B1_ready_in(SB_T3_EAST_SB_OUT_B1_ready_and_Z),
    .SB_T3_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1_valid_out),
    .SB_T3_NORTH_SB_IN_B1(SB_T3_NORTH_SB_IN_B1),
    .SB_T3_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_IN_B1_enable),
    .SB_T3_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_IN_B1_ready_out),
    .SB_T3_NORTH_SB_IN_B1_valid_in(SB_T3_NORTH_SB_IN_B1_valid),
    .SB_T3_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1_enable),
    .SB_T3_NORTH_SB_OUT_B1_ready_in(SB_T3_NORTH_SB_OUT_B1_ready_and_Z),
    .SB_T3_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1_valid_out),
    .SB_T3_SOUTH_SB_IN_B1(SB_T3_SOUTH_SB_IN_B1),
    .SB_T3_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_IN_B1_enable),
    .SB_T3_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_IN_B1_ready_out),
    .SB_T3_SOUTH_SB_IN_B1_valid_in(SB_T3_SOUTH_SB_IN_B1_valid),
    .SB_T3_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1_enable),
    .SB_T3_SOUTH_SB_OUT_B1_ready_in(SB_T3_SOUTH_SB_OUT_B1_ready_and_Z),
    .SB_T3_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1_valid_out),
    .SB_T3_WEST_SB_IN_B1(SB_T3_WEST_SB_IN_B1),
    .SB_T3_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_IN_B1_enable),
    .SB_T3_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_IN_B1_ready_out),
    .SB_T3_WEST_SB_IN_B1_valid_in(SB_T3_WEST_SB_IN_B1_valid),
    .SB_T3_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1_enable),
    .SB_T3_WEST_SB_OUT_B1_ready_in(SB_T3_WEST_SB_OUT_B1_ready_and_Z),
    .SB_T3_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1_valid_out),
    .SB_T4_EAST_SB_IN_B1(SB_T4_EAST_SB_IN_B1),
    .SB_T4_EAST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_IN_B1_enable),
    .SB_T4_EAST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_IN_B1_ready_out),
    .SB_T4_EAST_SB_IN_B1_valid_in(SB_T4_EAST_SB_IN_B1_valid),
    .SB_T4_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1_enable),
    .SB_T4_EAST_SB_OUT_B1_ready_in(SB_T4_EAST_SB_OUT_B1_ready_and_Z),
    .SB_T4_EAST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1_valid_out),
    .SB_T4_NORTH_SB_IN_B1(SB_T4_NORTH_SB_IN_B1),
    .SB_T4_NORTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_IN_B1_enable),
    .SB_T4_NORTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_IN_B1_ready_out),
    .SB_T4_NORTH_SB_IN_B1_valid_in(SB_T4_NORTH_SB_IN_B1_valid),
    .SB_T4_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1_enable),
    .SB_T4_NORTH_SB_OUT_B1_ready_in(SB_T4_NORTH_SB_OUT_B1_ready_and_Z),
    .SB_T4_NORTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1_valid_out),
    .SB_T4_SOUTH_SB_IN_B1(SB_T4_SOUTH_SB_IN_B1),
    .SB_T4_SOUTH_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_IN_B1_enable),
    .SB_T4_SOUTH_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_IN_B1_ready_out),
    .SB_T4_SOUTH_SB_IN_B1_valid_in(SB_T4_SOUTH_SB_IN_B1_valid),
    .SB_T4_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1_enable),
    .SB_T4_SOUTH_SB_OUT_B1_ready_in(SB_T4_SOUTH_SB_OUT_B1_ready_and_Z),
    .SB_T4_SOUTH_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1_valid_out),
    .SB_T4_WEST_SB_IN_B1(SB_T4_WEST_SB_IN_B1),
    .SB_T4_WEST_SB_IN_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_IN_B1_enable),
    .SB_T4_WEST_SB_IN_B1_ready_out(SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_IN_B1_ready_out),
    .SB_T4_WEST_SB_IN_B1_valid_in(SB_T4_WEST_SB_IN_B1_valid),
    .SB_T4_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B1_enable(SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1_enable),
    .SB_T4_WEST_SB_OUT_B1_ready_in(SB_T4_WEST_SB_OUT_B1_ready_and_Z),
    .SB_T4_WEST_SB_OUT_B1_valid_out(SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1_valid_out),
    .clk(clk),
    .config_config_addr(self_config_config_addr_out[31:24]),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_10_out),
    .read_config_data(SB_ID0_5TRACKS_B1_MemCore_read_config_data),
    .reset(reset),
    .stall(stall)
);
and_cell SB_T0_EAST_SB_OUT_B17_ready_and (
    .A(SB_T0_EAST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_OUT_B17_enable),
    .Z(SB_T0_EAST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T0_EAST_SB_OUT_B1_ready_and (
    .A(SB_T0_EAST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1_enable),
    .Z(SB_T0_EAST_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T0_NORTH_SB_OUT_B17_ready_and (
    .A(SB_T0_NORTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_OUT_B17_enable),
    .Z(SB_T0_NORTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T0_NORTH_SB_OUT_B1_ready_and (
    .A(SB_T0_NORTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1_enable),
    .Z(SB_T0_NORTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T0_SOUTH_SB_OUT_B17_ready_and (
    .A(SB_T0_SOUTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_OUT_B17_enable),
    .Z(SB_T0_SOUTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T0_SOUTH_SB_OUT_B1_ready_and (
    .A(SB_T0_SOUTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1_enable),
    .Z(SB_T0_SOUTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T0_WEST_SB_OUT_B17_ready_and (
    .A(SB_T0_WEST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_OUT_B17_enable),
    .Z(SB_T0_WEST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T0_WEST_SB_OUT_B1_ready_and (
    .A(SB_T0_WEST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1_enable),
    .Z(SB_T0_WEST_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T1_EAST_SB_OUT_B17_ready_and (
    .A(SB_T1_EAST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_OUT_B17_enable),
    .Z(SB_T1_EAST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T1_EAST_SB_OUT_B1_ready_and (
    .A(SB_T1_EAST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1_enable),
    .Z(SB_T1_EAST_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T1_NORTH_SB_OUT_B17_ready_and (
    .A(SB_T1_NORTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_OUT_B17_enable),
    .Z(SB_T1_NORTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T1_NORTH_SB_OUT_B1_ready_and (
    .A(SB_T1_NORTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1_enable),
    .Z(SB_T1_NORTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T1_SOUTH_SB_OUT_B17_ready_and (
    .A(SB_T1_SOUTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_OUT_B17_enable),
    .Z(SB_T1_SOUTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T1_SOUTH_SB_OUT_B1_ready_and (
    .A(SB_T1_SOUTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1_enable),
    .Z(SB_T1_SOUTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T1_WEST_SB_OUT_B17_ready_and (
    .A(SB_T1_WEST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_OUT_B17_enable),
    .Z(SB_T1_WEST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T1_WEST_SB_OUT_B1_ready_and (
    .A(SB_T1_WEST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1_enable),
    .Z(SB_T1_WEST_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T2_EAST_SB_OUT_B17_ready_and (
    .A(SB_T2_EAST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_OUT_B17_enable),
    .Z(SB_T2_EAST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T2_EAST_SB_OUT_B1_ready_and (
    .A(SB_T2_EAST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1_enable),
    .Z(SB_T2_EAST_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T2_NORTH_SB_OUT_B17_ready_and (
    .A(SB_T2_NORTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_OUT_B17_enable),
    .Z(SB_T2_NORTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T2_NORTH_SB_OUT_B1_ready_and (
    .A(SB_T2_NORTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1_enable),
    .Z(SB_T2_NORTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T2_SOUTH_SB_OUT_B17_ready_and (
    .A(SB_T2_SOUTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_OUT_B17_enable),
    .Z(SB_T2_SOUTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T2_SOUTH_SB_OUT_B1_ready_and (
    .A(SB_T2_SOUTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1_enable),
    .Z(SB_T2_SOUTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T2_WEST_SB_OUT_B17_ready_and (
    .A(SB_T2_WEST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_OUT_B17_enable),
    .Z(SB_T2_WEST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T2_WEST_SB_OUT_B1_ready_and (
    .A(SB_T2_WEST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1_enable),
    .Z(SB_T2_WEST_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T3_EAST_SB_OUT_B17_ready_and (
    .A(SB_T3_EAST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_OUT_B17_enable),
    .Z(SB_T3_EAST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T3_EAST_SB_OUT_B1_ready_and (
    .A(SB_T3_EAST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1_enable),
    .Z(SB_T3_EAST_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T3_NORTH_SB_OUT_B17_ready_and (
    .A(SB_T3_NORTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_OUT_B17_enable),
    .Z(SB_T3_NORTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T3_NORTH_SB_OUT_B1_ready_and (
    .A(SB_T3_NORTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1_enable),
    .Z(SB_T3_NORTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T3_SOUTH_SB_OUT_B17_ready_and (
    .A(SB_T3_SOUTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_OUT_B17_enable),
    .Z(SB_T3_SOUTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T3_SOUTH_SB_OUT_B1_ready_and (
    .A(SB_T3_SOUTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1_enable),
    .Z(SB_T3_SOUTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T3_WEST_SB_OUT_B17_ready_and (
    .A(SB_T3_WEST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_OUT_B17_enable),
    .Z(SB_T3_WEST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T3_WEST_SB_OUT_B1_ready_and (
    .A(SB_T3_WEST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1_enable),
    .Z(SB_T3_WEST_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T4_EAST_SB_OUT_B17_ready_and (
    .A(SB_T4_EAST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_OUT_B17_enable),
    .Z(SB_T4_EAST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T4_EAST_SB_OUT_B1_ready_and (
    .A(SB_T4_EAST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1_enable),
    .Z(SB_T4_EAST_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T4_NORTH_SB_OUT_B17_ready_and (
    .A(SB_T4_NORTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_OUT_B17_enable),
    .Z(SB_T4_NORTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T4_NORTH_SB_OUT_B1_ready_and (
    .A(SB_T4_NORTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1_enable),
    .Z(SB_T4_NORTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T4_SOUTH_SB_OUT_B17_ready_and (
    .A(SB_T4_SOUTH_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_OUT_B17_enable),
    .Z(SB_T4_SOUTH_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T4_SOUTH_SB_OUT_B1_ready_and (
    .A(SB_T4_SOUTH_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1_enable),
    .Z(SB_T4_SOUTH_SB_OUT_B1_ready_and_Z)
);
and_cell SB_T4_WEST_SB_OUT_B17_ready_and (
    .A(SB_T4_WEST_SB_OUT_B17_ready),
    .B(SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_OUT_B17_enable),
    .Z(SB_T4_WEST_SB_OUT_B17_ready_and_Z)
);
and_cell SB_T4_WEST_SB_OUT_B1_ready_and (
    .A(SB_T4_WEST_SB_OUT_B1_ready),
    .B(SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1_enable),
    .Z(SB_T4_WEST_SB_OUT_B1_ready_and_Z)
);
corebit_and and_inst0 (
    .in0(coreir_eq_16_inst0_out),
    .in1(config_read[0]),
    .out(and_inst0_out)
);
corebit_and and_inst1 (
    .in0(coreir_eq_16_inst0_out),
    .in1(config_write[0]),
    .out(and_inst1_out)
);
corebit_const #(
    .value(1'b1)
) bit_const_1_None (
    .out(bit_const_1_None_out)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
coreir_const #(
    .value(9'h1ff),
    .width(9)
) const_511_9 (
    .out(const_511_9_out)
);
coreir_eq #(
    .width(16)
) coreir_eq_16_inst0 (
    .in0(tile_id),
    .in1(self_config_config_addr_out[15:0]),
    .out(coreir_eq_16_inst0_out)
);
wire [31:0] read_data_mux_I [12:0];
assign read_data_mux_I[12] = PowerDomainConfigReg_inst0_read_config_data;
assign read_data_mux_I[11] = SB_ID0_5TRACKS_B17_MemCore_read_config_data;
assign read_data_mux_I[10] = SB_ID0_5TRACKS_B1_MemCore_read_config_data;
assign read_data_mux_I[9] = CB_flush_read_config_data;
assign read_data_mux_I[8] = CB_MEM_input_width_1_num_1_read_config_data;
assign read_data_mux_I[7] = CB_MEM_input_width_1_num_0_read_config_data;
assign read_data_mux_I[6] = CB_MEM_input_width_17_num_3_read_config_data;
assign read_data_mux_I[5] = CB_MEM_input_width_17_num_2_read_config_data;
assign read_data_mux_I[4] = CB_MEM_input_width_17_num_1_read_config_data;
assign read_data_mux_I[3] = CB_MEM_input_width_17_num_0_read_config_data;
assign read_data_mux_I[2] = MemCore_inst0_read_config_data_2;
assign read_data_mux_I[1] = MemCore_inst0_read_config_data_1;
assign read_data_mux_I[0] = MemCore_inst0_read_config_data;
MuxWithDefaultWrapper_13_32_8_0 read_data_mux (
    .I(read_data_mux_I),
    .S(self_config_config_addr_out[23:16]),
    .EN(and_inst0_out),
    .O(read_data_mux_O)
);
mantle_wire__typeBit32 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
assign SB_T0_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_IN_B17_ready_out;
assign SB_T0_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_IN_B1_ready_out;
assign SB_T0_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1;
assign SB_T0_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_OUT_B17;
assign SB_T0_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T0_EAST_SB_OUT_B17_valid_out;
assign SB_T0_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1_valid_out;
assign SB_T0_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_IN_B17_ready_out;
assign SB_T0_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_IN_B1_ready_out;
assign SB_T0_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1;
assign SB_T0_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_OUT_B17;
assign SB_T0_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T0_NORTH_SB_OUT_B17_valid_out;
assign SB_T0_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1_valid_out;
assign SB_T0_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_IN_B17_ready_out;
assign SB_T0_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_IN_B1_ready_out;
assign SB_T0_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1;
assign SB_T0_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_OUT_B17;
assign SB_T0_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T0_SOUTH_SB_OUT_B17_valid_out;
assign SB_T0_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1_valid_out;
assign SB_T0_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_IN_B17_ready_out;
assign SB_T0_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_IN_B1_ready_out;
assign SB_T0_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1;
assign SB_T0_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_OUT_B17;
assign SB_T0_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T0_WEST_SB_OUT_B17_valid_out;
assign SB_T0_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1_valid_out;
assign SB_T1_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_IN_B17_ready_out;
assign SB_T1_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_IN_B1_ready_out;
assign SB_T1_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1;
assign SB_T1_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_OUT_B17;
assign SB_T1_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T1_EAST_SB_OUT_B17_valid_out;
assign SB_T1_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1_valid_out;
assign SB_T1_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_IN_B17_ready_out;
assign SB_T1_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_IN_B1_ready_out;
assign SB_T1_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1;
assign SB_T1_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_OUT_B17;
assign SB_T1_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T1_NORTH_SB_OUT_B17_valid_out;
assign SB_T1_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1_valid_out;
assign SB_T1_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_IN_B17_ready_out;
assign SB_T1_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_IN_B1_ready_out;
assign SB_T1_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1;
assign SB_T1_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_OUT_B17;
assign SB_T1_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T1_SOUTH_SB_OUT_B17_valid_out;
assign SB_T1_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1_valid_out;
assign SB_T1_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_IN_B17_ready_out;
assign SB_T1_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_IN_B1_ready_out;
assign SB_T1_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1;
assign SB_T1_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_OUT_B17;
assign SB_T1_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T1_WEST_SB_OUT_B17_valid_out;
assign SB_T1_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1_valid_out;
assign SB_T2_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_IN_B17_ready_out;
assign SB_T2_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_IN_B1_ready_out;
assign SB_T2_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1;
assign SB_T2_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_OUT_B17;
assign SB_T2_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T2_EAST_SB_OUT_B17_valid_out;
assign SB_T2_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1_valid_out;
assign SB_T2_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_IN_B17_ready_out;
assign SB_T2_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_IN_B1_ready_out;
assign SB_T2_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1;
assign SB_T2_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_OUT_B17;
assign SB_T2_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T2_NORTH_SB_OUT_B17_valid_out;
assign SB_T2_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1_valid_out;
assign SB_T2_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_IN_B17_ready_out;
assign SB_T2_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_IN_B1_ready_out;
assign SB_T2_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1;
assign SB_T2_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_OUT_B17;
assign SB_T2_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T2_SOUTH_SB_OUT_B17_valid_out;
assign SB_T2_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1_valid_out;
assign SB_T2_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_IN_B17_ready_out;
assign SB_T2_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_IN_B1_ready_out;
assign SB_T2_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1;
assign SB_T2_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_OUT_B17;
assign SB_T2_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T2_WEST_SB_OUT_B17_valid_out;
assign SB_T2_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1_valid_out;
assign SB_T3_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_IN_B17_ready_out;
assign SB_T3_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_IN_B1_ready_out;
assign SB_T3_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1;
assign SB_T3_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_OUT_B17;
assign SB_T3_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T3_EAST_SB_OUT_B17_valid_out;
assign SB_T3_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1_valid_out;
assign SB_T3_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_IN_B17_ready_out;
assign SB_T3_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_IN_B1_ready_out;
assign SB_T3_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1;
assign SB_T3_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_OUT_B17;
assign SB_T3_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T3_NORTH_SB_OUT_B17_valid_out;
assign SB_T3_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1_valid_out;
assign SB_T3_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_IN_B17_ready_out;
assign SB_T3_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_IN_B1_ready_out;
assign SB_T3_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1;
assign SB_T3_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_OUT_B17;
assign SB_T3_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T3_SOUTH_SB_OUT_B17_valid_out;
assign SB_T3_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1_valid_out;
assign SB_T3_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_IN_B17_ready_out;
assign SB_T3_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_IN_B1_ready_out;
assign SB_T3_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1;
assign SB_T3_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_OUT_B17;
assign SB_T3_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T3_WEST_SB_OUT_B17_valid_out;
assign SB_T3_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1_valid_out;
assign SB_T4_EAST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_IN_B17_ready_out;
assign SB_T4_EAST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_IN_B1_ready_out;
assign SB_T4_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1;
assign SB_T4_EAST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_OUT_B17;
assign SB_T4_EAST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T4_EAST_SB_OUT_B17_valid_out;
assign SB_T4_EAST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1_valid_out;
assign SB_T4_NORTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_IN_B17_ready_out;
assign SB_T4_NORTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_IN_B1_ready_out;
assign SB_T4_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1;
assign SB_T4_NORTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_OUT_B17;
assign SB_T4_NORTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T4_NORTH_SB_OUT_B17_valid_out;
assign SB_T4_NORTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1_valid_out;
assign SB_T4_SOUTH_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_IN_B17_ready_out;
assign SB_T4_SOUTH_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_IN_B1_ready_out;
assign SB_T4_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1;
assign SB_T4_SOUTH_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_OUT_B17;
assign SB_T4_SOUTH_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T4_SOUTH_SB_OUT_B17_valid_out;
assign SB_T4_SOUTH_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1_valid_out;
assign SB_T4_WEST_SB_IN_B17_ready = SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_IN_B17_ready_out;
assign SB_T4_WEST_SB_IN_B1_ready = SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_IN_B1_ready_out;
assign SB_T4_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1;
assign SB_T4_WEST_SB_OUT_B17 = SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_OUT_B17;
assign SB_T4_WEST_SB_OUT_B17_valid = SB_ID0_5TRACKS_B17_MemCore_SB_T4_WEST_SB_OUT_B17_valid_out;
assign SB_T4_WEST_SB_OUT_B1_valid = SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1_valid_out;
assign clk_out = clk;
assign config_out_config_addr = config_config_addr;
assign config_out_config_data = config_config_data;
assign config_out_read = config_read;
assign config_out_write = config_write;
assign flush_out = flush;
assign hi = const_511_9_out;
assign lo = const_0_8_out;
assign read_config_data = PowerDomainOR_O;
assign reset_out = reset;
assign stall_out = stall;
endmodule

module Interconnect (
    input clk,
    input [31:0] config_0_config_addr,
    input [31:0] config_0_config_data,
    input [0:0] config_0_read,
    input [0:0] config_0_write,
    input [31:0] config_1_config_addr,
    input [31:0] config_1_config_data,
    input [0:0] config_1_read,
    input [0:0] config_1_write,
    input [31:0] config_2_config_addr,
    input [31:0] config_2_config_data,
    input [0:0] config_2_read,
    input [0:0] config_2_write,
    input [31:0] config_3_config_addr,
    input [31:0] config_3_config_data,
    input [0:0] config_3_read,
    input [0:0] config_3_write,
    input [0:0] flush,
    input [16:0] glb2io_17_X00_Y00,
    output glb2io_17_X00_Y00_ready,
    input glb2io_17_X00_Y00_valid,
    input [16:0] glb2io_17_X01_Y00,
    output glb2io_17_X01_Y00_ready,
    input glb2io_17_X01_Y00_valid,
    input [16:0] glb2io_17_X02_Y00,
    output glb2io_17_X02_Y00_ready,
    input glb2io_17_X02_Y00_valid,
    input [16:0] glb2io_17_X03_Y00,
    output glb2io_17_X03_Y00_ready,
    input glb2io_17_X03_Y00_valid,
    input [0:0] glb2io_1_X00_Y00,
    output glb2io_1_X00_Y00_ready,
    input glb2io_1_X00_Y00_valid,
    input [0:0] glb2io_1_X01_Y00,
    output glb2io_1_X01_Y00_ready,
    input glb2io_1_X01_Y00_valid,
    input [0:0] glb2io_1_X02_Y00,
    output glb2io_1_X02_Y00_ready,
    input glb2io_1_X02_Y00_valid,
    input [0:0] glb2io_1_X03_Y00,
    output glb2io_1_X03_Y00_ready,
    input glb2io_1_X03_Y00_valid,
    output [16:0] io2glb_17_X00_Y00,
    input io2glb_17_X00_Y00_ready,
    output io2glb_17_X00_Y00_valid,
    output [16:0] io2glb_17_X01_Y00,
    input io2glb_17_X01_Y00_ready,
    output io2glb_17_X01_Y00_valid,
    output [16:0] io2glb_17_X02_Y00,
    input io2glb_17_X02_Y00_ready,
    output io2glb_17_X02_Y00_valid,
    output [16:0] io2glb_17_X03_Y00,
    input io2glb_17_X03_Y00_ready,
    output io2glb_17_X03_Y00_valid,
    output [0:0] io2glb_1_X00_Y00,
    input io2glb_1_X00_Y00_ready,
    output io2glb_1_X00_Y00_valid,
    output [0:0] io2glb_1_X01_Y00,
    input io2glb_1_X01_Y00_ready,
    output io2glb_1_X01_Y00_valid,
    output [0:0] io2glb_1_X02_Y00,
    input io2glb_1_X02_Y00_ready,
    output io2glb_1_X02_Y00_valid,
    output [0:0] io2glb_1_X03_Y00,
    input io2glb_1_X03_Y00_ready,
    output io2glb_1_X03_Y00_valid,
    output [31:0] read_config_data,
    input reset,
    input [3:0] stall
);
wire [0:0] PipelineRegister_inst0$Register_inst0$reg_P1_inst0_out;
wire [0:0] PipelineRegister_inst1$Register_inst0$reg_P1_inst0_out;
wire [0:0] PipelineRegister_inst2$Register_inst0$reg_P1_inst0_out;
wire [0:0] PipelineRegister_inst3$Register_inst0$reg_P1_inst0_out;
wire [65:0] PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out;
wire [65:0] PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out;
wire [65:0] PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out;
wire [65:0] PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out;
wire Tile_X00_Y00_clk_out;
wire [31:0] Tile_X00_Y00_config_out_config_addr;
wire [31:0] Tile_X00_Y00_config_out_config_data;
wire [0:0] Tile_X00_Y00_config_out_read;
wire [0:0] Tile_X00_Y00_config_out_write;
wire Tile_X00_Y00_f2io_17_ready;
wire Tile_X00_Y00_f2io_1_ready;
wire [0:0] Tile_X00_Y00_flush_out;
wire Tile_X00_Y00_glb2io_17_ready;
wire Tile_X00_Y00_glb2io_1_ready;
wire [8:0] Tile_X00_Y00_hi;
wire [0:0] Tile_X00_Y00_io2f_1;
wire [16:0] Tile_X00_Y00_io2f_17;
wire Tile_X00_Y00_io2f_17_valid;
wire Tile_X00_Y00_io2f_1_valid;
wire [0:0] Tile_X00_Y00_io2glb_1;
wire [16:0] Tile_X00_Y00_io2glb_17;
wire Tile_X00_Y00_io2glb_17_valid;
wire Tile_X00_Y00_io2glb_1_valid;
wire [7:0] Tile_X00_Y00_lo;
wire [31:0] Tile_X00_Y00_read_config_data;
wire Tile_X00_Y00_reset_out;
wire [0:0] Tile_X00_Y00_stall_out;
wire Tile_X00_Y01_SB_T0_EAST_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T0_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T0_EAST_SB_OUT_B17;
wire Tile_X00_Y01_SB_T0_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T0_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T0_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B17;
wire Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T0_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T0_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B17;
wire Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T0_WEST_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T0_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T0_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T0_WEST_SB_OUT_B17;
wire Tile_X00_Y01_SB_T0_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T0_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T1_EAST_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T1_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T1_EAST_SB_OUT_B17;
wire Tile_X00_Y01_SB_T1_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T1_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T1_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B17;
wire Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T1_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T1_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B17;
wire Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T1_WEST_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T1_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T1_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T1_WEST_SB_OUT_B17;
wire Tile_X00_Y01_SB_T1_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T1_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T2_EAST_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T2_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T2_EAST_SB_OUT_B17;
wire Tile_X00_Y01_SB_T2_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T2_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T2_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B17;
wire Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T2_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T2_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B17;
wire Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T2_WEST_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T2_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T2_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T2_WEST_SB_OUT_B17;
wire Tile_X00_Y01_SB_T2_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T2_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T3_EAST_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T3_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T3_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T3_EAST_SB_OUT_B17;
wire Tile_X00_Y01_SB_T3_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T3_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T3_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T3_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B17;
wire Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T3_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T3_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B17;
wire Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T3_WEST_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T3_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T3_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T3_WEST_SB_OUT_B17;
wire Tile_X00_Y01_SB_T3_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T3_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T4_EAST_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T4_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T4_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T4_EAST_SB_OUT_B17;
wire Tile_X00_Y01_SB_T4_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T4_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T4_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T4_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B17;
wire Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T4_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T4_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B17;
wire Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y01_SB_T4_WEST_SB_IN_B17_ready;
wire Tile_X00_Y01_SB_T4_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y01_SB_T4_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y01_SB_T4_WEST_SB_OUT_B17;
wire Tile_X00_Y01_SB_T4_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y01_SB_T4_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y01_clk_out;
wire Tile_X00_Y01_clk_pass_through_out_bot;
wire Tile_X00_Y01_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y01_config_out_config_addr;
wire [31:0] Tile_X00_Y01_config_out_config_data;
wire [0:0] Tile_X00_Y01_config_out_read;
wire [0:0] Tile_X00_Y01_config_out_write;
wire [0:0] Tile_X00_Y01_flush_out;
wire [8:0] Tile_X00_Y01_hi;
wire [7:0] Tile_X00_Y01_lo;
wire [31:0] Tile_X00_Y01_read_config_data;
wire Tile_X00_Y01_reset_out;
wire [0:0] Tile_X00_Y01_stall_out;
wire Tile_X00_Y02_SB_T0_EAST_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T0_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T0_EAST_SB_OUT_B17;
wire Tile_X00_Y02_SB_T0_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T0_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T0_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B17;
wire Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T0_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T0_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B17;
wire Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T0_WEST_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T0_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T0_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T0_WEST_SB_OUT_B17;
wire Tile_X00_Y02_SB_T0_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T0_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T1_EAST_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T1_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T1_EAST_SB_OUT_B17;
wire Tile_X00_Y02_SB_T1_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T1_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T1_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B17;
wire Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T1_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T1_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B17;
wire Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T1_WEST_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T1_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T1_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T1_WEST_SB_OUT_B17;
wire Tile_X00_Y02_SB_T1_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T1_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T2_EAST_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T2_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T2_EAST_SB_OUT_B17;
wire Tile_X00_Y02_SB_T2_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T2_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T2_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B17;
wire Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T2_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T2_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B17;
wire Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T2_WEST_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T2_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T2_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T2_WEST_SB_OUT_B17;
wire Tile_X00_Y02_SB_T2_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T2_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T3_EAST_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T3_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T3_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T3_EAST_SB_OUT_B17;
wire Tile_X00_Y02_SB_T3_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T3_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T3_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T3_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B17;
wire Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T3_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T3_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B17;
wire Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T3_WEST_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T3_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T3_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T3_WEST_SB_OUT_B17;
wire Tile_X00_Y02_SB_T3_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T3_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T4_EAST_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T4_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T4_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T4_EAST_SB_OUT_B17;
wire Tile_X00_Y02_SB_T4_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T4_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T4_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T4_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B17;
wire Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T4_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T4_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B17;
wire Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y02_SB_T4_WEST_SB_IN_B17_ready;
wire Tile_X00_Y02_SB_T4_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y02_SB_T4_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y02_SB_T4_WEST_SB_OUT_B17;
wire Tile_X00_Y02_SB_T4_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y02_SB_T4_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y02_clk_out;
wire Tile_X00_Y02_clk_pass_through_out_bot;
wire Tile_X00_Y02_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y02_config_out_config_addr;
wire [31:0] Tile_X00_Y02_config_out_config_data;
wire [0:0] Tile_X00_Y02_config_out_read;
wire [0:0] Tile_X00_Y02_config_out_write;
wire [0:0] Tile_X00_Y02_flush_out;
wire [8:0] Tile_X00_Y02_hi;
wire [7:0] Tile_X00_Y02_lo;
wire [31:0] Tile_X00_Y02_read_config_data;
wire Tile_X00_Y02_reset_out;
wire [0:0] Tile_X00_Y02_stall_out;
wire Tile_X00_Y03_SB_T0_EAST_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T0_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T0_EAST_SB_OUT_B17;
wire Tile_X00_Y03_SB_T0_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T0_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T0_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B17;
wire Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T0_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T0_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B17;
wire Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T0_WEST_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T0_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T0_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T0_WEST_SB_OUT_B17;
wire Tile_X00_Y03_SB_T0_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T0_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T1_EAST_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T1_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T1_EAST_SB_OUT_B17;
wire Tile_X00_Y03_SB_T1_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T1_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T1_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B17;
wire Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T1_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T1_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B17;
wire Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T1_WEST_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T1_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T1_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T1_WEST_SB_OUT_B17;
wire Tile_X00_Y03_SB_T1_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T1_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T2_EAST_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T2_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T2_EAST_SB_OUT_B17;
wire Tile_X00_Y03_SB_T2_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T2_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T2_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B17;
wire Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T2_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T2_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B17;
wire Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T2_WEST_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T2_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T2_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T2_WEST_SB_OUT_B17;
wire Tile_X00_Y03_SB_T2_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T2_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T3_EAST_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T3_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T3_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T3_EAST_SB_OUT_B17;
wire Tile_X00_Y03_SB_T3_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T3_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T3_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T3_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B17;
wire Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T3_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T3_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B17;
wire Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T3_WEST_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T3_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T3_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T3_WEST_SB_OUT_B17;
wire Tile_X00_Y03_SB_T3_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T3_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T4_EAST_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T4_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T4_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T4_EAST_SB_OUT_B17;
wire Tile_X00_Y03_SB_T4_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T4_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T4_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T4_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B17;
wire Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T4_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T4_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B17;
wire Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y03_SB_T4_WEST_SB_IN_B17_ready;
wire Tile_X00_Y03_SB_T4_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y03_SB_T4_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y03_SB_T4_WEST_SB_OUT_B17;
wire Tile_X00_Y03_SB_T4_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y03_SB_T4_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y03_clk_out;
wire Tile_X00_Y03_clk_pass_through_out_bot;
wire Tile_X00_Y03_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y03_config_out_config_addr;
wire [31:0] Tile_X00_Y03_config_out_config_data;
wire [0:0] Tile_X00_Y03_config_out_read;
wire [0:0] Tile_X00_Y03_config_out_write;
wire [0:0] Tile_X00_Y03_flush_out;
wire [8:0] Tile_X00_Y03_hi;
wire [7:0] Tile_X00_Y03_lo;
wire [31:0] Tile_X00_Y03_read_config_data;
wire Tile_X00_Y03_reset_out;
wire [0:0] Tile_X00_Y03_stall_out;
wire Tile_X00_Y04_SB_T0_EAST_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T0_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T0_EAST_SB_OUT_B17;
wire Tile_X00_Y04_SB_T0_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T0_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T0_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B17;
wire Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T0_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T0_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B17;
wire Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T0_WEST_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T0_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T0_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T0_WEST_SB_OUT_B17;
wire Tile_X00_Y04_SB_T0_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T0_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T1_EAST_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T1_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T1_EAST_SB_OUT_B17;
wire Tile_X00_Y04_SB_T1_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T1_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T1_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B17;
wire Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T1_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T1_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B17;
wire Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T1_WEST_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T1_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T1_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T1_WEST_SB_OUT_B17;
wire Tile_X00_Y04_SB_T1_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T1_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T2_EAST_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T2_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T2_EAST_SB_OUT_B17;
wire Tile_X00_Y04_SB_T2_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T2_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T2_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B17;
wire Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T2_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T2_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B17;
wire Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T2_WEST_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T2_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T2_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T2_WEST_SB_OUT_B17;
wire Tile_X00_Y04_SB_T2_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T2_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T3_EAST_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T3_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T3_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T3_EAST_SB_OUT_B17;
wire Tile_X00_Y04_SB_T3_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T3_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T3_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T3_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B17;
wire Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T3_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T3_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B17;
wire Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T3_WEST_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T3_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T3_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T3_WEST_SB_OUT_B17;
wire Tile_X00_Y04_SB_T3_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T3_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T4_EAST_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T4_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T4_EAST_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T4_EAST_SB_OUT_B17;
wire Tile_X00_Y04_SB_T4_EAST_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T4_EAST_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T4_NORTH_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T4_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B17;
wire Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T4_SOUTH_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T4_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B17;
wire Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B1_valid;
wire Tile_X00_Y04_SB_T4_WEST_SB_IN_B17_ready;
wire Tile_X00_Y04_SB_T4_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X00_Y04_SB_T4_WEST_SB_OUT_B1;
wire [16:0] Tile_X00_Y04_SB_T4_WEST_SB_OUT_B17;
wire Tile_X00_Y04_SB_T4_WEST_SB_OUT_B17_valid;
wire Tile_X00_Y04_SB_T4_WEST_SB_OUT_B1_valid;
wire Tile_X00_Y04_clk_out;
wire Tile_X00_Y04_clk_pass_through_out_bot;
wire Tile_X00_Y04_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y04_config_out_config_addr;
wire [31:0] Tile_X00_Y04_config_out_config_data;
wire [0:0] Tile_X00_Y04_config_out_read;
wire [0:0] Tile_X00_Y04_config_out_write;
wire [0:0] Tile_X00_Y04_flush_out;
wire [8:0] Tile_X00_Y04_hi;
wire [7:0] Tile_X00_Y04_lo;
wire [31:0] Tile_X00_Y04_read_config_data;
wire Tile_X00_Y04_reset_out;
wire [0:0] Tile_X00_Y04_stall_out;
wire Tile_X01_Y00_clk_out;
wire [31:0] Tile_X01_Y00_config_out_config_addr;
wire [31:0] Tile_X01_Y00_config_out_config_data;
wire [0:0] Tile_X01_Y00_config_out_read;
wire [0:0] Tile_X01_Y00_config_out_write;
wire Tile_X01_Y00_f2io_17_ready;
wire Tile_X01_Y00_f2io_1_ready;
wire [0:0] Tile_X01_Y00_flush_out;
wire Tile_X01_Y00_glb2io_17_ready;
wire Tile_X01_Y00_glb2io_1_ready;
wire [8:0] Tile_X01_Y00_hi;
wire [0:0] Tile_X01_Y00_io2f_1;
wire [16:0] Tile_X01_Y00_io2f_17;
wire Tile_X01_Y00_io2f_17_valid;
wire Tile_X01_Y00_io2f_1_valid;
wire [0:0] Tile_X01_Y00_io2glb_1;
wire [16:0] Tile_X01_Y00_io2glb_17;
wire Tile_X01_Y00_io2glb_17_valid;
wire Tile_X01_Y00_io2glb_1_valid;
wire [7:0] Tile_X01_Y00_lo;
wire [31:0] Tile_X01_Y00_read_config_data;
wire Tile_X01_Y00_reset_out;
wire [0:0] Tile_X01_Y00_stall_out;
wire Tile_X01_Y01_SB_T0_EAST_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T0_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T0_EAST_SB_OUT_B17;
wire Tile_X01_Y01_SB_T0_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T0_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T0_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B17;
wire Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T0_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T0_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B17;
wire Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T0_WEST_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T0_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T0_WEST_SB_OUT_B17;
wire Tile_X01_Y01_SB_T0_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T1_EAST_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T1_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T1_EAST_SB_OUT_B17;
wire Tile_X01_Y01_SB_T1_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T1_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T1_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B17;
wire Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T1_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T1_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B17;
wire Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T1_WEST_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T1_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T1_WEST_SB_OUT_B17;
wire Tile_X01_Y01_SB_T1_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T2_EAST_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T2_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T2_EAST_SB_OUT_B17;
wire Tile_X01_Y01_SB_T2_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T2_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T2_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B17;
wire Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T2_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T2_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B17;
wire Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T2_WEST_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T2_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T2_WEST_SB_OUT_B17;
wire Tile_X01_Y01_SB_T2_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T3_EAST_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T3_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T3_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T3_EAST_SB_OUT_B17;
wire Tile_X01_Y01_SB_T3_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T3_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T3_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T3_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B17;
wire Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T3_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T3_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B17;
wire Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T3_WEST_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T3_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T3_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T3_WEST_SB_OUT_B17;
wire Tile_X01_Y01_SB_T3_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T3_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T4_EAST_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T4_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T4_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T4_EAST_SB_OUT_B17;
wire Tile_X01_Y01_SB_T4_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T4_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T4_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T4_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B17;
wire Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T4_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T4_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B17;
wire Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y01_SB_T4_WEST_SB_IN_B17_ready;
wire Tile_X01_Y01_SB_T4_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y01_SB_T4_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y01_SB_T4_WEST_SB_OUT_B17;
wire Tile_X01_Y01_SB_T4_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y01_SB_T4_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y01_clk_out;
wire Tile_X01_Y01_clk_pass_through_out_bot;
wire Tile_X01_Y01_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y01_config_out_config_addr;
wire [31:0] Tile_X01_Y01_config_out_config_data;
wire [0:0] Tile_X01_Y01_config_out_read;
wire [0:0] Tile_X01_Y01_config_out_write;
wire [0:0] Tile_X01_Y01_flush_out;
wire [8:0] Tile_X01_Y01_hi;
wire [7:0] Tile_X01_Y01_lo;
wire [31:0] Tile_X01_Y01_read_config_data;
wire Tile_X01_Y01_reset_out;
wire [0:0] Tile_X01_Y01_stall_out;
wire Tile_X01_Y02_SB_T0_EAST_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T0_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T0_EAST_SB_OUT_B17;
wire Tile_X01_Y02_SB_T0_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T0_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T0_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B17;
wire Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T0_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T0_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B17;
wire Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T0_WEST_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T0_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T0_WEST_SB_OUT_B17;
wire Tile_X01_Y02_SB_T0_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T1_EAST_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T1_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T1_EAST_SB_OUT_B17;
wire Tile_X01_Y02_SB_T1_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T1_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T1_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B17;
wire Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T1_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T1_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B17;
wire Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T1_WEST_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T1_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T1_WEST_SB_OUT_B17;
wire Tile_X01_Y02_SB_T1_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T2_EAST_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T2_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T2_EAST_SB_OUT_B17;
wire Tile_X01_Y02_SB_T2_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T2_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T2_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B17;
wire Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T2_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T2_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B17;
wire Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T2_WEST_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T2_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T2_WEST_SB_OUT_B17;
wire Tile_X01_Y02_SB_T2_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T3_EAST_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T3_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T3_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T3_EAST_SB_OUT_B17;
wire Tile_X01_Y02_SB_T3_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T3_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T3_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T3_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B17;
wire Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T3_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T3_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B17;
wire Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T3_WEST_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T3_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T3_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T3_WEST_SB_OUT_B17;
wire Tile_X01_Y02_SB_T3_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T3_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T4_EAST_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T4_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T4_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T4_EAST_SB_OUT_B17;
wire Tile_X01_Y02_SB_T4_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T4_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T4_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T4_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B17;
wire Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T4_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T4_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B17;
wire Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y02_SB_T4_WEST_SB_IN_B17_ready;
wire Tile_X01_Y02_SB_T4_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y02_SB_T4_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y02_SB_T4_WEST_SB_OUT_B17;
wire Tile_X01_Y02_SB_T4_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y02_SB_T4_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y02_clk_out;
wire Tile_X01_Y02_clk_pass_through_out_bot;
wire Tile_X01_Y02_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y02_config_out_config_addr;
wire [31:0] Tile_X01_Y02_config_out_config_data;
wire [0:0] Tile_X01_Y02_config_out_read;
wire [0:0] Tile_X01_Y02_config_out_write;
wire [0:0] Tile_X01_Y02_flush_out;
wire [8:0] Tile_X01_Y02_hi;
wire [7:0] Tile_X01_Y02_lo;
wire [31:0] Tile_X01_Y02_read_config_data;
wire Tile_X01_Y02_reset_out;
wire [0:0] Tile_X01_Y02_stall_out;
wire Tile_X01_Y03_SB_T0_EAST_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T0_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T0_EAST_SB_OUT_B17;
wire Tile_X01_Y03_SB_T0_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T0_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T0_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B17;
wire Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T0_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T0_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B17;
wire Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T0_WEST_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T0_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T0_WEST_SB_OUT_B17;
wire Tile_X01_Y03_SB_T0_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T1_EAST_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T1_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T1_EAST_SB_OUT_B17;
wire Tile_X01_Y03_SB_T1_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T1_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T1_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B17;
wire Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T1_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T1_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B17;
wire Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T1_WEST_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T1_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T1_WEST_SB_OUT_B17;
wire Tile_X01_Y03_SB_T1_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T2_EAST_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T2_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T2_EAST_SB_OUT_B17;
wire Tile_X01_Y03_SB_T2_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T2_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T2_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B17;
wire Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T2_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T2_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B17;
wire Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T2_WEST_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T2_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T2_WEST_SB_OUT_B17;
wire Tile_X01_Y03_SB_T2_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T3_EAST_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T3_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T3_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T3_EAST_SB_OUT_B17;
wire Tile_X01_Y03_SB_T3_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T3_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T3_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T3_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B17;
wire Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T3_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T3_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B17;
wire Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T3_WEST_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T3_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T3_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T3_WEST_SB_OUT_B17;
wire Tile_X01_Y03_SB_T3_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T3_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T4_EAST_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T4_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T4_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T4_EAST_SB_OUT_B17;
wire Tile_X01_Y03_SB_T4_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T4_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T4_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T4_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B17;
wire Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T4_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T4_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B17;
wire Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y03_SB_T4_WEST_SB_IN_B17_ready;
wire Tile_X01_Y03_SB_T4_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y03_SB_T4_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y03_SB_T4_WEST_SB_OUT_B17;
wire Tile_X01_Y03_SB_T4_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y03_SB_T4_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y03_clk_out;
wire Tile_X01_Y03_clk_pass_through_out_bot;
wire Tile_X01_Y03_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y03_config_out_config_addr;
wire [31:0] Tile_X01_Y03_config_out_config_data;
wire [0:0] Tile_X01_Y03_config_out_read;
wire [0:0] Tile_X01_Y03_config_out_write;
wire [0:0] Tile_X01_Y03_flush_out;
wire [8:0] Tile_X01_Y03_hi;
wire [7:0] Tile_X01_Y03_lo;
wire [31:0] Tile_X01_Y03_read_config_data;
wire Tile_X01_Y03_reset_out;
wire [0:0] Tile_X01_Y03_stall_out;
wire Tile_X01_Y04_SB_T0_EAST_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T0_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T0_EAST_SB_OUT_B17;
wire Tile_X01_Y04_SB_T0_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T0_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T0_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B17;
wire Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T0_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T0_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B17;
wire Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T0_WEST_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T0_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T0_WEST_SB_OUT_B17;
wire Tile_X01_Y04_SB_T0_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T1_EAST_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T1_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T1_EAST_SB_OUT_B17;
wire Tile_X01_Y04_SB_T1_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T1_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T1_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B17;
wire Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T1_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T1_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B17;
wire Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T1_WEST_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T1_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T1_WEST_SB_OUT_B17;
wire Tile_X01_Y04_SB_T1_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T2_EAST_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T2_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T2_EAST_SB_OUT_B17;
wire Tile_X01_Y04_SB_T2_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T2_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T2_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B17;
wire Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T2_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T2_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B17;
wire Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T2_WEST_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T2_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T2_WEST_SB_OUT_B17;
wire Tile_X01_Y04_SB_T2_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T3_EAST_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T3_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T3_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T3_EAST_SB_OUT_B17;
wire Tile_X01_Y04_SB_T3_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T3_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T3_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T3_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B17;
wire Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T3_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T3_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B17;
wire Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T3_WEST_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T3_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T3_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T3_WEST_SB_OUT_B17;
wire Tile_X01_Y04_SB_T3_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T3_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T4_EAST_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T4_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T4_EAST_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T4_EAST_SB_OUT_B17;
wire Tile_X01_Y04_SB_T4_EAST_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T4_EAST_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T4_NORTH_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T4_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B17;
wire Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T4_SOUTH_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T4_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B17;
wire Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B1_valid;
wire Tile_X01_Y04_SB_T4_WEST_SB_IN_B17_ready;
wire Tile_X01_Y04_SB_T4_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X01_Y04_SB_T4_WEST_SB_OUT_B1;
wire [16:0] Tile_X01_Y04_SB_T4_WEST_SB_OUT_B17;
wire Tile_X01_Y04_SB_T4_WEST_SB_OUT_B17_valid;
wire Tile_X01_Y04_SB_T4_WEST_SB_OUT_B1_valid;
wire Tile_X01_Y04_clk_out;
wire Tile_X01_Y04_clk_pass_through_out_bot;
wire Tile_X01_Y04_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y04_config_out_config_addr;
wire [31:0] Tile_X01_Y04_config_out_config_data;
wire [0:0] Tile_X01_Y04_config_out_read;
wire [0:0] Tile_X01_Y04_config_out_write;
wire [0:0] Tile_X01_Y04_flush_out;
wire [8:0] Tile_X01_Y04_hi;
wire [7:0] Tile_X01_Y04_lo;
wire [31:0] Tile_X01_Y04_read_config_data;
wire Tile_X01_Y04_reset_out;
wire [0:0] Tile_X01_Y04_stall_out;
wire Tile_X02_Y00_clk_out;
wire [31:0] Tile_X02_Y00_config_out_config_addr;
wire [31:0] Tile_X02_Y00_config_out_config_data;
wire [0:0] Tile_X02_Y00_config_out_read;
wire [0:0] Tile_X02_Y00_config_out_write;
wire Tile_X02_Y00_f2io_17_ready;
wire Tile_X02_Y00_f2io_1_ready;
wire [0:0] Tile_X02_Y00_flush_out;
wire Tile_X02_Y00_glb2io_17_ready;
wire Tile_X02_Y00_glb2io_1_ready;
wire [8:0] Tile_X02_Y00_hi;
wire [0:0] Tile_X02_Y00_io2f_1;
wire [16:0] Tile_X02_Y00_io2f_17;
wire Tile_X02_Y00_io2f_17_valid;
wire Tile_X02_Y00_io2f_1_valid;
wire [0:0] Tile_X02_Y00_io2glb_1;
wire [16:0] Tile_X02_Y00_io2glb_17;
wire Tile_X02_Y00_io2glb_17_valid;
wire Tile_X02_Y00_io2glb_1_valid;
wire [7:0] Tile_X02_Y00_lo;
wire [31:0] Tile_X02_Y00_read_config_data;
wire Tile_X02_Y00_reset_out;
wire [0:0] Tile_X02_Y00_stall_out;
wire Tile_X02_Y01_SB_T0_EAST_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T0_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T0_EAST_SB_OUT_B17;
wire Tile_X02_Y01_SB_T0_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T0_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T0_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B17;
wire Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T0_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T0_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B17;
wire Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T0_WEST_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T0_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T0_WEST_SB_OUT_B17;
wire Tile_X02_Y01_SB_T0_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T1_EAST_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T1_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T1_EAST_SB_OUT_B17;
wire Tile_X02_Y01_SB_T1_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T1_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T1_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B17;
wire Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T1_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T1_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B17;
wire Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T1_WEST_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T1_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T1_WEST_SB_OUT_B17;
wire Tile_X02_Y01_SB_T1_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T2_EAST_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T2_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T2_EAST_SB_OUT_B17;
wire Tile_X02_Y01_SB_T2_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T2_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T2_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B17;
wire Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T2_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T2_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B17;
wire Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T2_WEST_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T2_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T2_WEST_SB_OUT_B17;
wire Tile_X02_Y01_SB_T2_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T3_EAST_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T3_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T3_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T3_EAST_SB_OUT_B17;
wire Tile_X02_Y01_SB_T3_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T3_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T3_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T3_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B17;
wire Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T3_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T3_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B17;
wire Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T3_WEST_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T3_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T3_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T3_WEST_SB_OUT_B17;
wire Tile_X02_Y01_SB_T3_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T3_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T4_EAST_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T4_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T4_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T4_EAST_SB_OUT_B17;
wire Tile_X02_Y01_SB_T4_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T4_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T4_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T4_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B17;
wire Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T4_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T4_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B17;
wire Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y01_SB_T4_WEST_SB_IN_B17_ready;
wire Tile_X02_Y01_SB_T4_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y01_SB_T4_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y01_SB_T4_WEST_SB_OUT_B17;
wire Tile_X02_Y01_SB_T4_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y01_SB_T4_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y01_clk_out;
wire Tile_X02_Y01_clk_pass_through_out_bot;
wire Tile_X02_Y01_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y01_config_out_config_addr;
wire [31:0] Tile_X02_Y01_config_out_config_data;
wire [0:0] Tile_X02_Y01_config_out_read;
wire [0:0] Tile_X02_Y01_config_out_write;
wire [0:0] Tile_X02_Y01_flush_out;
wire [8:0] Tile_X02_Y01_hi;
wire [7:0] Tile_X02_Y01_lo;
wire [31:0] Tile_X02_Y01_read_config_data;
wire Tile_X02_Y01_reset_out;
wire [0:0] Tile_X02_Y01_stall_out;
wire Tile_X02_Y02_SB_T0_EAST_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T0_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T0_EAST_SB_OUT_B17;
wire Tile_X02_Y02_SB_T0_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T0_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T0_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B17;
wire Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T0_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T0_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B17;
wire Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T0_WEST_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T0_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T0_WEST_SB_OUT_B17;
wire Tile_X02_Y02_SB_T0_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T1_EAST_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T1_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T1_EAST_SB_OUT_B17;
wire Tile_X02_Y02_SB_T1_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T1_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T1_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B17;
wire Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T1_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T1_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B17;
wire Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T1_WEST_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T1_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T1_WEST_SB_OUT_B17;
wire Tile_X02_Y02_SB_T1_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T2_EAST_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T2_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T2_EAST_SB_OUT_B17;
wire Tile_X02_Y02_SB_T2_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T2_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T2_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B17;
wire Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T2_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T2_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B17;
wire Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T2_WEST_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T2_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T2_WEST_SB_OUT_B17;
wire Tile_X02_Y02_SB_T2_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T3_EAST_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T3_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T3_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T3_EAST_SB_OUT_B17;
wire Tile_X02_Y02_SB_T3_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T3_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T3_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T3_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B17;
wire Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T3_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T3_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B17;
wire Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T3_WEST_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T3_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T3_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T3_WEST_SB_OUT_B17;
wire Tile_X02_Y02_SB_T3_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T3_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T4_EAST_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T4_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T4_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T4_EAST_SB_OUT_B17;
wire Tile_X02_Y02_SB_T4_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T4_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T4_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T4_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B17;
wire Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T4_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T4_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B17;
wire Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y02_SB_T4_WEST_SB_IN_B17_ready;
wire Tile_X02_Y02_SB_T4_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y02_SB_T4_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y02_SB_T4_WEST_SB_OUT_B17;
wire Tile_X02_Y02_SB_T4_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y02_SB_T4_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y02_clk_out;
wire Tile_X02_Y02_clk_pass_through_out_bot;
wire Tile_X02_Y02_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y02_config_out_config_addr;
wire [31:0] Tile_X02_Y02_config_out_config_data;
wire [0:0] Tile_X02_Y02_config_out_read;
wire [0:0] Tile_X02_Y02_config_out_write;
wire [0:0] Tile_X02_Y02_flush_out;
wire [8:0] Tile_X02_Y02_hi;
wire [7:0] Tile_X02_Y02_lo;
wire [31:0] Tile_X02_Y02_read_config_data;
wire Tile_X02_Y02_reset_out;
wire [0:0] Tile_X02_Y02_stall_out;
wire Tile_X02_Y03_SB_T0_EAST_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T0_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T0_EAST_SB_OUT_B17;
wire Tile_X02_Y03_SB_T0_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T0_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T0_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B17;
wire Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T0_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T0_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B17;
wire Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T0_WEST_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T0_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T0_WEST_SB_OUT_B17;
wire Tile_X02_Y03_SB_T0_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T1_EAST_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T1_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T1_EAST_SB_OUT_B17;
wire Tile_X02_Y03_SB_T1_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T1_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T1_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B17;
wire Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T1_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T1_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B17;
wire Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T1_WEST_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T1_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T1_WEST_SB_OUT_B17;
wire Tile_X02_Y03_SB_T1_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T2_EAST_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T2_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T2_EAST_SB_OUT_B17;
wire Tile_X02_Y03_SB_T2_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T2_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T2_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B17;
wire Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T2_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T2_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B17;
wire Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T2_WEST_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T2_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T2_WEST_SB_OUT_B17;
wire Tile_X02_Y03_SB_T2_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T3_EAST_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T3_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T3_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T3_EAST_SB_OUT_B17;
wire Tile_X02_Y03_SB_T3_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T3_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T3_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T3_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B17;
wire Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T3_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T3_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B17;
wire Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T3_WEST_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T3_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T3_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T3_WEST_SB_OUT_B17;
wire Tile_X02_Y03_SB_T3_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T3_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T4_EAST_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T4_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T4_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T4_EAST_SB_OUT_B17;
wire Tile_X02_Y03_SB_T4_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T4_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T4_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T4_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B17;
wire Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T4_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T4_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B17;
wire Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y03_SB_T4_WEST_SB_IN_B17_ready;
wire Tile_X02_Y03_SB_T4_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y03_SB_T4_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y03_SB_T4_WEST_SB_OUT_B17;
wire Tile_X02_Y03_SB_T4_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y03_SB_T4_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y03_clk_out;
wire Tile_X02_Y03_clk_pass_through_out_bot;
wire Tile_X02_Y03_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y03_config_out_config_addr;
wire [31:0] Tile_X02_Y03_config_out_config_data;
wire [0:0] Tile_X02_Y03_config_out_read;
wire [0:0] Tile_X02_Y03_config_out_write;
wire [0:0] Tile_X02_Y03_flush_out;
wire [8:0] Tile_X02_Y03_hi;
wire [7:0] Tile_X02_Y03_lo;
wire [31:0] Tile_X02_Y03_read_config_data;
wire Tile_X02_Y03_reset_out;
wire [0:0] Tile_X02_Y03_stall_out;
wire Tile_X02_Y04_SB_T0_EAST_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T0_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T0_EAST_SB_OUT_B17;
wire Tile_X02_Y04_SB_T0_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T0_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T0_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B17;
wire Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T0_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T0_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B17;
wire Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T0_WEST_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T0_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T0_WEST_SB_OUT_B17;
wire Tile_X02_Y04_SB_T0_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T1_EAST_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T1_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T1_EAST_SB_OUT_B17;
wire Tile_X02_Y04_SB_T1_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T1_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T1_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B17;
wire Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T1_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T1_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B17;
wire Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T1_WEST_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T1_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T1_WEST_SB_OUT_B17;
wire Tile_X02_Y04_SB_T1_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T2_EAST_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T2_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T2_EAST_SB_OUT_B17;
wire Tile_X02_Y04_SB_T2_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T2_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T2_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B17;
wire Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T2_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T2_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B17;
wire Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T2_WEST_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T2_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T2_WEST_SB_OUT_B17;
wire Tile_X02_Y04_SB_T2_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T3_EAST_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T3_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T3_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T3_EAST_SB_OUT_B17;
wire Tile_X02_Y04_SB_T3_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T3_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T3_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T3_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B17;
wire Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T3_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T3_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B17;
wire Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T3_WEST_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T3_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T3_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T3_WEST_SB_OUT_B17;
wire Tile_X02_Y04_SB_T3_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T3_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T4_EAST_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T4_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T4_EAST_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T4_EAST_SB_OUT_B17;
wire Tile_X02_Y04_SB_T4_EAST_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T4_EAST_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T4_NORTH_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T4_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B17;
wire Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T4_SOUTH_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T4_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B17;
wire Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B1_valid;
wire Tile_X02_Y04_SB_T4_WEST_SB_IN_B17_ready;
wire Tile_X02_Y04_SB_T4_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X02_Y04_SB_T4_WEST_SB_OUT_B1;
wire [16:0] Tile_X02_Y04_SB_T4_WEST_SB_OUT_B17;
wire Tile_X02_Y04_SB_T4_WEST_SB_OUT_B17_valid;
wire Tile_X02_Y04_SB_T4_WEST_SB_OUT_B1_valid;
wire Tile_X02_Y04_clk_out;
wire Tile_X02_Y04_clk_pass_through_out_bot;
wire Tile_X02_Y04_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y04_config_out_config_addr;
wire [31:0] Tile_X02_Y04_config_out_config_data;
wire [0:0] Tile_X02_Y04_config_out_read;
wire [0:0] Tile_X02_Y04_config_out_write;
wire [0:0] Tile_X02_Y04_flush_out;
wire [8:0] Tile_X02_Y04_hi;
wire [7:0] Tile_X02_Y04_lo;
wire [31:0] Tile_X02_Y04_read_config_data;
wire Tile_X02_Y04_reset_out;
wire [0:0] Tile_X02_Y04_stall_out;
wire Tile_X03_Y00_clk_out;
wire [31:0] Tile_X03_Y00_config_out_config_addr;
wire [31:0] Tile_X03_Y00_config_out_config_data;
wire [0:0] Tile_X03_Y00_config_out_read;
wire [0:0] Tile_X03_Y00_config_out_write;
wire Tile_X03_Y00_f2io_17_ready;
wire Tile_X03_Y00_f2io_1_ready;
wire [0:0] Tile_X03_Y00_flush_out;
wire Tile_X03_Y00_glb2io_17_ready;
wire Tile_X03_Y00_glb2io_1_ready;
wire [8:0] Tile_X03_Y00_hi;
wire [0:0] Tile_X03_Y00_io2f_1;
wire [16:0] Tile_X03_Y00_io2f_17;
wire Tile_X03_Y00_io2f_17_valid;
wire Tile_X03_Y00_io2f_1_valid;
wire [0:0] Tile_X03_Y00_io2glb_1;
wire [16:0] Tile_X03_Y00_io2glb_17;
wire Tile_X03_Y00_io2glb_17_valid;
wire Tile_X03_Y00_io2glb_1_valid;
wire [7:0] Tile_X03_Y00_lo;
wire [31:0] Tile_X03_Y00_read_config_data;
wire Tile_X03_Y00_reset_out;
wire [0:0] Tile_X03_Y00_stall_out;
wire Tile_X03_Y01_SB_T0_EAST_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T0_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T0_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T0_EAST_SB_OUT_B17;
wire Tile_X03_Y01_SB_T0_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T0_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T0_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T0_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B17;
wire Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T0_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T0_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B17;
wire Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T0_WEST_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T0_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T0_WEST_SB_OUT_B17;
wire Tile_X03_Y01_SB_T0_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T1_EAST_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T1_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T1_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T1_EAST_SB_OUT_B17;
wire Tile_X03_Y01_SB_T1_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T1_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T1_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T1_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B17;
wire Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T1_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T1_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B17;
wire Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T1_WEST_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T1_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T1_WEST_SB_OUT_B17;
wire Tile_X03_Y01_SB_T1_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T2_EAST_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T2_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T2_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T2_EAST_SB_OUT_B17;
wire Tile_X03_Y01_SB_T2_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T2_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T2_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T2_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B17;
wire Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T2_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T2_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B17;
wire Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T2_WEST_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T2_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T2_WEST_SB_OUT_B17;
wire Tile_X03_Y01_SB_T2_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T3_EAST_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T3_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T3_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T3_EAST_SB_OUT_B17;
wire Tile_X03_Y01_SB_T3_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T3_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T3_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T3_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B17;
wire Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T3_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T3_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B17;
wire Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T3_WEST_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T3_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T3_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T3_WEST_SB_OUT_B17;
wire Tile_X03_Y01_SB_T3_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T3_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T4_EAST_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T4_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T4_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T4_EAST_SB_OUT_B17;
wire Tile_X03_Y01_SB_T4_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T4_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T4_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T4_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B17;
wire Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T4_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T4_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B17;
wire Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y01_SB_T4_WEST_SB_IN_B17_ready;
wire Tile_X03_Y01_SB_T4_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y01_SB_T4_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y01_SB_T4_WEST_SB_OUT_B17;
wire Tile_X03_Y01_SB_T4_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y01_SB_T4_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y01_clk_out;
wire [31:0] Tile_X03_Y01_config_out_config_addr;
wire [31:0] Tile_X03_Y01_config_out_config_data;
wire [0:0] Tile_X03_Y01_config_out_read;
wire [0:0] Tile_X03_Y01_config_out_write;
wire [0:0] Tile_X03_Y01_flush_out;
wire [8:0] Tile_X03_Y01_hi;
wire [7:0] Tile_X03_Y01_lo;
wire [31:0] Tile_X03_Y01_read_config_data;
wire Tile_X03_Y01_reset_out;
wire [0:0] Tile_X03_Y01_stall_out;
wire Tile_X03_Y02_SB_T0_EAST_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T0_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T0_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T0_EAST_SB_OUT_B17;
wire Tile_X03_Y02_SB_T0_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T0_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T0_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T0_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B17;
wire Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T0_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T0_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B17;
wire Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T0_WEST_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T0_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T0_WEST_SB_OUT_B17;
wire Tile_X03_Y02_SB_T0_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T1_EAST_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T1_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T1_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T1_EAST_SB_OUT_B17;
wire Tile_X03_Y02_SB_T1_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T1_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T1_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T1_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B17;
wire Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T1_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T1_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B17;
wire Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T1_WEST_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T1_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T1_WEST_SB_OUT_B17;
wire Tile_X03_Y02_SB_T1_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T2_EAST_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T2_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T2_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T2_EAST_SB_OUT_B17;
wire Tile_X03_Y02_SB_T2_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T2_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T2_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T2_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B17;
wire Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T2_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T2_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B17;
wire Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T2_WEST_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T2_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T2_WEST_SB_OUT_B17;
wire Tile_X03_Y02_SB_T2_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T3_EAST_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T3_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T3_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T3_EAST_SB_OUT_B17;
wire Tile_X03_Y02_SB_T3_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T3_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T3_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T3_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B17;
wire Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T3_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T3_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B17;
wire Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T3_WEST_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T3_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T3_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T3_WEST_SB_OUT_B17;
wire Tile_X03_Y02_SB_T3_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T3_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T4_EAST_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T4_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T4_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T4_EAST_SB_OUT_B17;
wire Tile_X03_Y02_SB_T4_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T4_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T4_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T4_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B17;
wire Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T4_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T4_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B17;
wire Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y02_SB_T4_WEST_SB_IN_B17_ready;
wire Tile_X03_Y02_SB_T4_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y02_SB_T4_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y02_SB_T4_WEST_SB_OUT_B17;
wire Tile_X03_Y02_SB_T4_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y02_SB_T4_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y02_clk_out;
wire [31:0] Tile_X03_Y02_config_out_config_addr;
wire [31:0] Tile_X03_Y02_config_out_config_data;
wire [0:0] Tile_X03_Y02_config_out_read;
wire [0:0] Tile_X03_Y02_config_out_write;
wire [0:0] Tile_X03_Y02_flush_out;
wire [8:0] Tile_X03_Y02_hi;
wire [7:0] Tile_X03_Y02_lo;
wire [31:0] Tile_X03_Y02_read_config_data;
wire Tile_X03_Y02_reset_out;
wire [0:0] Tile_X03_Y02_stall_out;
wire Tile_X03_Y03_SB_T0_EAST_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T0_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T0_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T0_EAST_SB_OUT_B17;
wire Tile_X03_Y03_SB_T0_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T0_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T0_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T0_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B17;
wire Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T0_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T0_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B17;
wire Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T0_WEST_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T0_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T0_WEST_SB_OUT_B17;
wire Tile_X03_Y03_SB_T0_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T1_EAST_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T1_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T1_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T1_EAST_SB_OUT_B17;
wire Tile_X03_Y03_SB_T1_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T1_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T1_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T1_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B17;
wire Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T1_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T1_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B17;
wire Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T1_WEST_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T1_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T1_WEST_SB_OUT_B17;
wire Tile_X03_Y03_SB_T1_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T2_EAST_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T2_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T2_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T2_EAST_SB_OUT_B17;
wire Tile_X03_Y03_SB_T2_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T2_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T2_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T2_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B17;
wire Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T2_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T2_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B17;
wire Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T2_WEST_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T2_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T2_WEST_SB_OUT_B17;
wire Tile_X03_Y03_SB_T2_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T3_EAST_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T3_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T3_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T3_EAST_SB_OUT_B17;
wire Tile_X03_Y03_SB_T3_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T3_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T3_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T3_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B17;
wire Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T3_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T3_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B17;
wire Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T3_WEST_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T3_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T3_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T3_WEST_SB_OUT_B17;
wire Tile_X03_Y03_SB_T3_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T3_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T4_EAST_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T4_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T4_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T4_EAST_SB_OUT_B17;
wire Tile_X03_Y03_SB_T4_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T4_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T4_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T4_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B17;
wire Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T4_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T4_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B17;
wire Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y03_SB_T4_WEST_SB_IN_B17_ready;
wire Tile_X03_Y03_SB_T4_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y03_SB_T4_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y03_SB_T4_WEST_SB_OUT_B17;
wire Tile_X03_Y03_SB_T4_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y03_SB_T4_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y03_clk_out;
wire [31:0] Tile_X03_Y03_config_out_config_addr;
wire [31:0] Tile_X03_Y03_config_out_config_data;
wire [0:0] Tile_X03_Y03_config_out_read;
wire [0:0] Tile_X03_Y03_config_out_write;
wire [0:0] Tile_X03_Y03_flush_out;
wire [8:0] Tile_X03_Y03_hi;
wire [7:0] Tile_X03_Y03_lo;
wire [31:0] Tile_X03_Y03_read_config_data;
wire Tile_X03_Y03_reset_out;
wire [0:0] Tile_X03_Y03_stall_out;
wire Tile_X03_Y04_SB_T0_EAST_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T0_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T0_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T0_EAST_SB_OUT_B17;
wire Tile_X03_Y04_SB_T0_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T0_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T0_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T0_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B17;
wire Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T0_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T0_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B17;
wire Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T0_WEST_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T0_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T0_WEST_SB_OUT_B17;
wire Tile_X03_Y04_SB_T0_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T1_EAST_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T1_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T1_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T1_EAST_SB_OUT_B17;
wire Tile_X03_Y04_SB_T1_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T1_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T1_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T1_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B17;
wire Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T1_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T1_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B17;
wire Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T1_WEST_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T1_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T1_WEST_SB_OUT_B17;
wire Tile_X03_Y04_SB_T1_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T2_EAST_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T2_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T2_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T2_EAST_SB_OUT_B17;
wire Tile_X03_Y04_SB_T2_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T2_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T2_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T2_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B17;
wire Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T2_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T2_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B17;
wire Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T2_WEST_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T2_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T2_WEST_SB_OUT_B17;
wire Tile_X03_Y04_SB_T2_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T3_EAST_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T3_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T3_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T3_EAST_SB_OUT_B17;
wire Tile_X03_Y04_SB_T3_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T3_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T3_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T3_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B17;
wire Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T3_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T3_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B17;
wire Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T3_WEST_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T3_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T3_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T3_WEST_SB_OUT_B17;
wire Tile_X03_Y04_SB_T3_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T3_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T4_EAST_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T4_EAST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T4_EAST_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T4_EAST_SB_OUT_B17;
wire Tile_X03_Y04_SB_T4_EAST_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T4_EAST_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T4_NORTH_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T4_NORTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B17;
wire Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T4_SOUTH_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T4_SOUTH_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B17;
wire Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B1_valid;
wire Tile_X03_Y04_SB_T4_WEST_SB_IN_B17_ready;
wire Tile_X03_Y04_SB_T4_WEST_SB_IN_B1_ready;
wire [0:0] Tile_X03_Y04_SB_T4_WEST_SB_OUT_B1;
wire [16:0] Tile_X03_Y04_SB_T4_WEST_SB_OUT_B17;
wire Tile_X03_Y04_SB_T4_WEST_SB_OUT_B17_valid;
wire Tile_X03_Y04_SB_T4_WEST_SB_OUT_B1_valid;
wire Tile_X03_Y04_clk_out;
wire [31:0] Tile_X03_Y04_config_out_config_addr;
wire [31:0] Tile_X03_Y04_config_out_config_data;
wire [0:0] Tile_X03_Y04_config_out_read;
wire [0:0] Tile_X03_Y04_config_out_write;
wire [0:0] Tile_X03_Y04_flush_out;
wire [8:0] Tile_X03_Y04_hi;
wire [7:0] Tile_X03_Y04_lo;
wire [31:0] Tile_X03_Y04_read_config_data;
wire Tile_X03_Y04_reset_out;
wire [0:0] Tile_X03_Y04_stall_out;
wire bit_const_0_None_out;
wire [0:0] const_0_1_out;
wire [16:0] const_0_17_out;
wire [31:0] const_0_32_out;
wire coreir_wrapInClock_inst0_out;
wire coreir_wrapInClock_inst1_out;
wire coreir_wrapInClock_inst2_out;
wire [31:0] read_config_data_or_final_O;
wire [3:0] self_stall_out;
coreir_reg #(
    .clk_posedge(1'b1),
    .init(1'h0),
    .width(1)
) PipelineRegister_inst0$Register_inst0$reg_P1_inst0 (
    .clk(clk),
    .in(flush),
    .out(PipelineRegister_inst0$Register_inst0$reg_P1_inst0_out)
);
coreir_reg #(
    .clk_posedge(1'b1),
    .init(1'h0),
    .width(1)
) PipelineRegister_inst1$Register_inst0$reg_P1_inst0 (
    .clk(clk),
    .in(flush),
    .out(PipelineRegister_inst1$Register_inst0$reg_P1_inst0_out)
);
coreir_reg #(
    .clk_posedge(1'b1),
    .init(1'h0),
    .width(1)
) PipelineRegister_inst2$Register_inst0$reg_P1_inst0 (
    .clk(clk),
    .in(flush),
    .out(PipelineRegister_inst2$Register_inst0$reg_P1_inst0_out)
);
coreir_reg #(
    .clk_posedge(1'b1),
    .init(1'h0),
    .width(1)
) PipelineRegister_inst3$Register_inst0$reg_P1_inst0 (
    .clk(clk),
    .in(flush),
    .out(PipelineRegister_inst3$Register_inst0$reg_P1_inst0_out)
);
wire [65:0] PipelineRegister_inst4$Register_inst0$reg_P66_inst0_in;
assign PipelineRegister_inst4$Register_inst0$reg_P66_inst0_in = {config_0_write[0],config_0_read[0],config_0_config_data,config_0_config_addr};
coreir_reg #(
    .clk_posedge(1'b1),
    .init(66'h00000000000000000),
    .width(66)
) PipelineRegister_inst4$Register_inst0$reg_P66_inst0 (
    .clk(clk),
    .in(PipelineRegister_inst4$Register_inst0$reg_P66_inst0_in),
    .out(PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out)
);
wire [65:0] PipelineRegister_inst5$Register_inst0$reg_P66_inst0_in;
assign PipelineRegister_inst5$Register_inst0$reg_P66_inst0_in = {config_1_write[0],config_1_read[0],config_1_config_data,config_1_config_addr};
coreir_reg #(
    .clk_posedge(1'b1),
    .init(66'h00000000000000000),
    .width(66)
) PipelineRegister_inst5$Register_inst0$reg_P66_inst0 (
    .clk(clk),
    .in(PipelineRegister_inst5$Register_inst0$reg_P66_inst0_in),
    .out(PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out)
);
wire [65:0] PipelineRegister_inst6$Register_inst0$reg_P66_inst0_in;
assign PipelineRegister_inst6$Register_inst0$reg_P66_inst0_in = {config_2_write[0],config_2_read[0],config_2_config_data,config_2_config_addr};
coreir_reg #(
    .clk_posedge(1'b1),
    .init(66'h00000000000000000),
    .width(66)
) PipelineRegister_inst6$Register_inst0$reg_P66_inst0 (
    .clk(clk),
    .in(PipelineRegister_inst6$Register_inst0$reg_P66_inst0_in),
    .out(PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out)
);
wire [65:0] PipelineRegister_inst7$Register_inst0$reg_P66_inst0_in;
assign PipelineRegister_inst7$Register_inst0$reg_P66_inst0_in = {config_3_write[0],config_3_read[0],config_3_config_data,config_3_config_addr};
coreir_reg #(
    .clk_posedge(1'b1),
    .init(66'h00000000000000000),
    .width(66)
) PipelineRegister_inst7$Register_inst0$reg_P66_inst0 (
    .clk(clk),
    .in(PipelineRegister_inst7$Register_inst0$reg_P66_inst0_in),
    .out(PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out)
);
wire [31:0] Tile_X00_Y00_config_config_addr;
assign Tile_X00_Y00_config_config_addr = {PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[31],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[30],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[29],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[28],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[27],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[26],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[25],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[24],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[23],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[22],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[21],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[20],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[19],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[18],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[17],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[16],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[15],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[14],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[13],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[12],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[11],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[10],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[9],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[8],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[7],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[6],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[5],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[4],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[3],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[2],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[1],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[0]};
wire [31:0] Tile_X00_Y00_config_config_data;
assign Tile_X00_Y00_config_config_data = {PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[63],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[62],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[61],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[60],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[59],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[58],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[57],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[56],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[55],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[54],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[53],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[52],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[51],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[50],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[49],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[48],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[47],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[46],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[45],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[44],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[43],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[42],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[41],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[40],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[39],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[38],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[37],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[36],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[35],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[34],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[33],PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[32]};
wire [4:0] Tile_X00_Y00_io2f_17_ready;
assign Tile_X00_Y00_io2f_17_ready = {Tile_X00_Y01_SB_T4_NORTH_SB_IN_B17_ready,Tile_X00_Y01_SB_T3_NORTH_SB_IN_B17_ready,Tile_X00_Y01_SB_T2_NORTH_SB_IN_B17_ready,Tile_X00_Y01_SB_T1_NORTH_SB_IN_B17_ready,Tile_X00_Y01_SB_T0_NORTH_SB_IN_B17_ready};
wire [4:0] Tile_X00_Y00_io2f_1_ready;
assign Tile_X00_Y00_io2f_1_ready = {Tile_X00_Y01_SB_T4_NORTH_SB_IN_B1_ready,Tile_X00_Y01_SB_T3_NORTH_SB_IN_B1_ready,Tile_X00_Y01_SB_T2_NORTH_SB_IN_B1_ready,Tile_X00_Y01_SB_T1_NORTH_SB_IN_B1_ready,Tile_X00_Y01_SB_T0_NORTH_SB_IN_B1_ready};
wire [15:0] Tile_X00_Y00_tile_id;
assign Tile_X00_Y00_tile_id = {Tile_X00_Y00_lo[7],Tile_X00_Y00_lo[7],Tile_X00_Y00_lo[6],Tile_X00_Y00_lo[6],Tile_X00_Y00_lo[5],Tile_X00_Y00_lo[5],Tile_X00_Y00_lo[4],Tile_X00_Y00_lo[4],Tile_X00_Y00_lo[3],Tile_X00_Y00_lo[3],Tile_X00_Y00_lo[2],Tile_X00_Y00_lo[2],Tile_X00_Y00_lo[1],Tile_X00_Y00_lo[1],Tile_X00_Y00_lo[0],Tile_X00_Y00_lo[0]};
Tile_IOCoreReadyValid Tile_X00_Y00 (
    .clk(clk),
    .clk_out(Tile_X00_Y00_clk_out),
    .config_config_addr(Tile_X00_Y00_config_config_addr),
    .config_config_data(Tile_X00_Y00_config_config_data),
    .config_out_config_addr(Tile_X00_Y00_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y00_config_out_config_data),
    .config_out_read(Tile_X00_Y00_config_out_read),
    .config_out_write(Tile_X00_Y00_config_out_write),
    .config_read(PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[64]),
    .config_write(PipelineRegister_inst4$Register_inst0$reg_P66_inst0_out[65]),
    .f2io_1(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1),
    .f2io_17(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B17),
    .f2io_17_ready(Tile_X00_Y00_f2io_17_ready),
    .f2io_17_valid(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B17_valid),
    .f2io_1_ready(Tile_X00_Y00_f2io_1_ready),
    .f2io_1_valid(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1_valid),
    .flush(PipelineRegister_inst0$Register_inst0$reg_P1_inst0_out),
    .flush_out(Tile_X00_Y00_flush_out),
    .glb2io_1(glb2io_1_X00_Y00),
    .glb2io_17(glb2io_17_X00_Y00),
    .glb2io_17_ready(Tile_X00_Y00_glb2io_17_ready),
    .glb2io_17_valid(glb2io_17_X00_Y00_valid),
    .glb2io_1_ready(Tile_X00_Y00_glb2io_1_ready),
    .glb2io_1_valid(glb2io_1_X00_Y00_valid),
    .hi(Tile_X00_Y00_hi),
    .io2f_1(Tile_X00_Y00_io2f_1),
    .io2f_17(Tile_X00_Y00_io2f_17),
    .io2f_17_ready(Tile_X00_Y00_io2f_17_ready),
    .io2f_17_valid(Tile_X00_Y00_io2f_17_valid),
    .io2f_1_ready(Tile_X00_Y00_io2f_1_ready),
    .io2f_1_valid(Tile_X00_Y00_io2f_1_valid),
    .io2glb_1(Tile_X00_Y00_io2glb_1),
    .io2glb_17(Tile_X00_Y00_io2glb_17),
    .io2glb_17_ready(io2glb_17_X00_Y00_ready),
    .io2glb_17_valid(Tile_X00_Y00_io2glb_17_valid),
    .io2glb_1_ready(io2glb_1_X00_Y00_ready),
    .io2glb_1_valid(Tile_X00_Y00_io2glb_1_valid),
    .lo(Tile_X00_Y00_lo),
    .read_config_data(Tile_X00_Y00_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X00_Y00_reset_out),
    .stall(self_stall_out[0:0]),
    .stall_out(Tile_X00_Y00_stall_out),
    .tile_id(Tile_X00_Y00_tile_id)
);
wire [15:0] Tile_X00_Y01_tile_id;
assign Tile_X00_Y01_tile_id = {Tile_X00_Y01_lo[7],Tile_X00_Y01_lo[7],Tile_X00_Y01_lo[6],Tile_X00_Y01_lo[6],Tile_X00_Y01_lo[5],Tile_X00_Y01_lo[5],Tile_X00_Y01_lo[4],Tile_X00_Y01_lo[4],Tile_X00_Y01_lo[3],Tile_X00_Y01_lo[3],Tile_X00_Y01_lo[2],Tile_X00_Y01_lo[2],Tile_X00_Y01_lo[1],Tile_X00_Y01_lo[1],Tile_X00_Y01_lo[0],Tile_X00_Y01_hi[0]};
Tile_PE Tile_X00_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B17(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_EAST_SB_IN_B17_ready(Tile_X00_Y01_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_IN_B17_valid(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_IN_B1_ready(Tile_X00_Y01_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_IN_B1_valid(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B17(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_EAST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B17(Tile_X00_Y00_io2f_17),
    .SB_T0_NORTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_IN_B17_valid(Tile_X00_Y00_io2f_17_valid),
    .SB_T0_NORTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_IN_B1_valid(Tile_X00_Y00_io2f_1_valid),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B17(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_OUT_B17_ready(Tile_X00_Y00_f2io_17_ready),
    .SB_T0_NORTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_OUT_B1_ready(Tile_X00_Y00_f2io_1_ready),
    .SB_T0_NORTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B17(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B17(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B17(const_0_17_out),
    .SB_T0_WEST_SB_IN_B17_ready(Tile_X00_Y01_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T0_WEST_SB_IN_B1_ready(Tile_X00_Y01_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B17(Tile_X00_Y01_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T0_WEST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T0_WEST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B17(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_EAST_SB_IN_B17_ready(Tile_X00_Y01_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_IN_B17_valid(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_IN_B1_ready(Tile_X00_Y01_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_IN_B1_valid(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B17(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_EAST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B17(Tile_X00_Y00_io2f_17),
    .SB_T1_NORTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_IN_B17_valid(Tile_X00_Y00_io2f_17_valid),
    .SB_T1_NORTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_IN_B1_valid(Tile_X00_Y00_io2f_1_valid),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B17(Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T1_NORTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T1_NORTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B17(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B17(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B17(const_0_17_out),
    .SB_T1_WEST_SB_IN_B17_ready(Tile_X00_Y01_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T1_WEST_SB_IN_B1_ready(Tile_X00_Y01_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B17(Tile_X00_Y01_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T1_WEST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T1_WEST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B17(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_EAST_SB_IN_B17_ready(Tile_X00_Y01_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_IN_B17_valid(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_IN_B1_ready(Tile_X00_Y01_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_IN_B1_valid(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B17(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_EAST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B17(Tile_X00_Y00_io2f_17),
    .SB_T2_NORTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_IN_B17_valid(Tile_X00_Y00_io2f_17_valid),
    .SB_T2_NORTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_IN_B1_valid(Tile_X00_Y00_io2f_1_valid),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B17(Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T2_NORTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T2_NORTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B17(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B17(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B17(const_0_17_out),
    .SB_T2_WEST_SB_IN_B17_ready(Tile_X00_Y01_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T2_WEST_SB_IN_B1_ready(Tile_X00_Y01_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B17(Tile_X00_Y01_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T2_WEST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T2_WEST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B17(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_EAST_SB_IN_B17_ready(Tile_X00_Y01_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_IN_B17_valid(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_IN_B1_ready(Tile_X00_Y01_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_IN_B1_valid(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B17(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_EAST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B17(Tile_X00_Y00_io2f_17),
    .SB_T3_NORTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_IN_B17_valid(Tile_X00_Y00_io2f_17_valid),
    .SB_T3_NORTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_IN_B1_valid(Tile_X00_Y00_io2f_1_valid),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B17(Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T3_NORTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T3_NORTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B17(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B17(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B17(const_0_17_out),
    .SB_T3_WEST_SB_IN_B17_ready(Tile_X00_Y01_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T3_WEST_SB_IN_B1_ready(Tile_X00_Y01_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B17(Tile_X00_Y01_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T3_WEST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T3_WEST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B17(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_EAST_SB_IN_B17_ready(Tile_X00_Y01_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_IN_B17_valid(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_IN_B1_ready(Tile_X00_Y01_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_IN_B1_valid(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B17(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_EAST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B17(Tile_X00_Y00_io2f_17),
    .SB_T4_NORTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_IN_B17_valid(Tile_X00_Y00_io2f_17_valid),
    .SB_T4_NORTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_IN_B1_valid(Tile_X00_Y00_io2f_1_valid),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B17(Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T4_NORTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T4_NORTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B17(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_IN_B17_ready(Tile_X00_Y01_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_IN_B1_ready(Tile_X00_Y01_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B17(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B17(const_0_17_out),
    .SB_T4_WEST_SB_IN_B17_ready(Tile_X00_Y01_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T4_WEST_SB_IN_B1_ready(Tile_X00_Y01_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B17(Tile_X00_Y01_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T4_WEST_SB_OUT_B17_valid(Tile_X00_Y01_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T4_WEST_SB_OUT_B1_valid(Tile_X00_Y01_SB_T4_WEST_SB_OUT_B1_valid),
    .clk(Tile_X00_Y00_clk_out),
    .clk_out(Tile_X00_Y01_clk_out),
    .clk_pass_through(coreir_wrapInClock_inst0_out),
    .clk_pass_through_out_bot(Tile_X00_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y01_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y00_config_out_config_addr),
    .config_config_data(Tile_X00_Y00_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y01_config_out_config_data),
    .config_out_read(Tile_X00_Y01_config_out_read),
    .config_out_write(Tile_X00_Y01_config_out_write),
    .config_read(Tile_X00_Y00_config_out_read),
    .config_write(Tile_X00_Y00_config_out_write),
    .flush(Tile_X00_Y00_flush_out),
    .flush_out(Tile_X00_Y01_flush_out),
    .hi(Tile_X00_Y01_hi),
    .lo(Tile_X00_Y01_lo),
    .read_config_data(Tile_X00_Y01_read_config_data),
    .read_config_data_in(Tile_X00_Y00_read_config_data),
    .reset(Tile_X00_Y00_reset_out),
    .reset_out(Tile_X00_Y01_reset_out),
    .stall(Tile_X00_Y00_stall_out),
    .stall_out(Tile_X00_Y01_stall_out),
    .tile_id(Tile_X00_Y01_tile_id)
);
wire [15:0] Tile_X00_Y02_tile_id;
assign Tile_X00_Y02_tile_id = {Tile_X00_Y02_lo[7],Tile_X00_Y02_lo[7],Tile_X00_Y02_lo[6],Tile_X00_Y02_lo[6],Tile_X00_Y02_lo[5],Tile_X00_Y02_lo[5],Tile_X00_Y02_lo[4],Tile_X00_Y02_lo[4],Tile_X00_Y02_lo[3],Tile_X00_Y02_lo[3],Tile_X00_Y02_lo[2],Tile_X00_Y02_lo[2],Tile_X00_Y02_lo[1],Tile_X00_Y02_lo[1],Tile_X00_Y02_hi[1],Tile_X00_Y02_lo[0]};
Tile_PE Tile_X00_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B17(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_EAST_SB_IN_B17_ready(Tile_X00_Y02_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_IN_B17_valid(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_IN_B1_ready(Tile_X00_Y02_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_IN_B1_valid(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B17(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_EAST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B17(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_IN_B17_valid(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_IN_B1_valid(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B17(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_OUT_B17_ready(Tile_X00_Y01_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_OUT_B1_ready(Tile_X00_Y01_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B17(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B17(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B17(const_0_17_out),
    .SB_T0_WEST_SB_IN_B17_ready(Tile_X00_Y02_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T0_WEST_SB_IN_B1_ready(Tile_X00_Y02_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B17(Tile_X00_Y02_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T0_WEST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T0_WEST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B17(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_EAST_SB_IN_B17_ready(Tile_X00_Y02_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_IN_B17_valid(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_IN_B1_ready(Tile_X00_Y02_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_IN_B1_valid(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B17(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_EAST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B17(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_IN_B17_valid(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_IN_B1_valid(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B17(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_OUT_B17_ready(Tile_X00_Y01_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_OUT_B1_ready(Tile_X00_Y01_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B17(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B17(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B17(const_0_17_out),
    .SB_T1_WEST_SB_IN_B17_ready(Tile_X00_Y02_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T1_WEST_SB_IN_B1_ready(Tile_X00_Y02_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B17(Tile_X00_Y02_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T1_WEST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T1_WEST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B17(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_EAST_SB_IN_B17_ready(Tile_X00_Y02_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_IN_B17_valid(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_IN_B1_ready(Tile_X00_Y02_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_IN_B1_valid(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B17(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_EAST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B17(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_IN_B17_valid(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_IN_B1_valid(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B17(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_OUT_B17_ready(Tile_X00_Y01_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_OUT_B1_ready(Tile_X00_Y01_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B17(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B17(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B17(const_0_17_out),
    .SB_T2_WEST_SB_IN_B17_ready(Tile_X00_Y02_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T2_WEST_SB_IN_B1_ready(Tile_X00_Y02_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B17(Tile_X00_Y02_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T2_WEST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T2_WEST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B17(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_EAST_SB_IN_B17_ready(Tile_X00_Y02_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_IN_B17_valid(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_IN_B1_ready(Tile_X00_Y02_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_IN_B1_valid(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B17(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_EAST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B17(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_IN_B17_valid(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_IN_B1_valid(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B17(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_OUT_B17_ready(Tile_X00_Y01_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_OUT_B1_ready(Tile_X00_Y01_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B17(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B17(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B17(const_0_17_out),
    .SB_T3_WEST_SB_IN_B17_ready(Tile_X00_Y02_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T3_WEST_SB_IN_B1_ready(Tile_X00_Y02_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B17(Tile_X00_Y02_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T3_WEST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T3_WEST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B17(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_EAST_SB_IN_B17_ready(Tile_X00_Y02_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_IN_B17_valid(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_IN_B1_ready(Tile_X00_Y02_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_IN_B1_valid(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B17(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_EAST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B17(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_IN_B17_valid(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_IN_B1_valid(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B17(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_OUT_B17_ready(Tile_X00_Y01_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_OUT_B1_ready(Tile_X00_Y01_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B17(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_IN_B17_ready(Tile_X00_Y02_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_IN_B1_ready(Tile_X00_Y02_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B17(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B17(const_0_17_out),
    .SB_T4_WEST_SB_IN_B17_ready(Tile_X00_Y02_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T4_WEST_SB_IN_B1_ready(Tile_X00_Y02_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B17(Tile_X00_Y02_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T4_WEST_SB_OUT_B17_valid(Tile_X00_Y02_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T4_WEST_SB_OUT_B1_valid(Tile_X00_Y02_SB_T4_WEST_SB_OUT_B1_valid),
    .clk(Tile_X00_Y01_clk_out),
    .clk_out(Tile_X00_Y02_clk_out),
    .clk_pass_through(Tile_X00_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y02_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y01_config_out_config_addr),
    .config_config_data(Tile_X00_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y02_config_out_config_data),
    .config_out_read(Tile_X00_Y02_config_out_read),
    .config_out_write(Tile_X00_Y02_config_out_write),
    .config_read(Tile_X00_Y01_config_out_read),
    .config_write(Tile_X00_Y01_config_out_write),
    .flush(Tile_X00_Y01_flush_out),
    .flush_out(Tile_X00_Y02_flush_out),
    .hi(Tile_X00_Y02_hi),
    .lo(Tile_X00_Y02_lo),
    .read_config_data(Tile_X00_Y02_read_config_data),
    .read_config_data_in(Tile_X00_Y01_read_config_data),
    .reset(Tile_X00_Y01_reset_out),
    .reset_out(Tile_X00_Y02_reset_out),
    .stall(Tile_X00_Y01_stall_out),
    .stall_out(Tile_X00_Y02_stall_out),
    .tile_id(Tile_X00_Y02_tile_id)
);
wire [15:0] Tile_X00_Y03_tile_id;
assign Tile_X00_Y03_tile_id = {Tile_X00_Y03_lo[7],Tile_X00_Y03_lo[7],Tile_X00_Y03_lo[6],Tile_X00_Y03_lo[6],Tile_X00_Y03_lo[5],Tile_X00_Y03_lo[5],Tile_X00_Y03_lo[4],Tile_X00_Y03_lo[4],Tile_X00_Y03_lo[3],Tile_X00_Y03_lo[3],Tile_X00_Y03_lo[2],Tile_X00_Y03_lo[2],Tile_X00_Y03_lo[1],Tile_X00_Y03_lo[1],Tile_X00_Y03_hi[1],Tile_X00_Y03_hi[0]};
Tile_PE Tile_X00_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B17(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_EAST_SB_IN_B17_ready(Tile_X00_Y03_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_IN_B17_valid(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_IN_B1_ready(Tile_X00_Y03_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_IN_B1_valid(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B17(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_EAST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B17(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B17(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B17(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_IN_B17_valid(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_IN_B1_valid(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B17(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X00_Y04_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X00_Y04_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B17(const_0_17_out),
    .SB_T0_WEST_SB_IN_B17_ready(Tile_X00_Y03_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T0_WEST_SB_IN_B1_ready(Tile_X00_Y03_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B17(Tile_X00_Y03_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T0_WEST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T0_WEST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B17(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_EAST_SB_IN_B17_ready(Tile_X00_Y03_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_IN_B17_valid(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_IN_B1_ready(Tile_X00_Y03_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_IN_B1_valid(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B17(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_EAST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B17(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B17(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B17(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_IN_B17_valid(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_IN_B1_valid(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B17(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X00_Y04_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X00_Y04_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B17(const_0_17_out),
    .SB_T1_WEST_SB_IN_B17_ready(Tile_X00_Y03_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T1_WEST_SB_IN_B1_ready(Tile_X00_Y03_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B17(Tile_X00_Y03_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T1_WEST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T1_WEST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B17(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_EAST_SB_IN_B17_ready(Tile_X00_Y03_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_IN_B17_valid(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_IN_B1_ready(Tile_X00_Y03_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_IN_B1_valid(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B17(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_EAST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B17(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B17(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B17(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_IN_B17_valid(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_IN_B1_valid(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B17(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X00_Y04_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X00_Y04_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B17(const_0_17_out),
    .SB_T2_WEST_SB_IN_B17_ready(Tile_X00_Y03_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T2_WEST_SB_IN_B1_ready(Tile_X00_Y03_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B17(Tile_X00_Y03_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T2_WEST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T2_WEST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B17(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_EAST_SB_IN_B17_ready(Tile_X00_Y03_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_IN_B17_valid(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_IN_B1_ready(Tile_X00_Y03_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_IN_B1_valid(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B17(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_EAST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B17(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B17(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B17(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_IN_B17_valid(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_IN_B1_valid(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B17(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X00_Y04_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X00_Y04_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B17(const_0_17_out),
    .SB_T3_WEST_SB_IN_B17_ready(Tile_X00_Y03_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T3_WEST_SB_IN_B1_ready(Tile_X00_Y03_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B17(Tile_X00_Y03_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T3_WEST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T3_WEST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B17(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_EAST_SB_IN_B17_ready(Tile_X00_Y03_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_IN_B17_valid(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_IN_B1_ready(Tile_X00_Y03_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_IN_B1_valid(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B17(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_EAST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B17(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_IN_B17_valid(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_IN_B1_valid(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B17(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_OUT_B17_ready(Tile_X00_Y02_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_OUT_B1_ready(Tile_X00_Y02_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B17(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_IN_B17_ready(Tile_X00_Y03_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_IN_B17_valid(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_IN_B1_ready(Tile_X00_Y03_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_IN_B1_valid(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B17(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X00_Y04_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X00_Y04_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B17(const_0_17_out),
    .SB_T4_WEST_SB_IN_B17_ready(Tile_X00_Y03_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T4_WEST_SB_IN_B1_ready(Tile_X00_Y03_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B17(Tile_X00_Y03_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T4_WEST_SB_OUT_B17_valid(Tile_X00_Y03_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T4_WEST_SB_OUT_B1_valid(Tile_X00_Y03_SB_T4_WEST_SB_OUT_B1_valid),
    .clk(Tile_X00_Y02_clk_out),
    .clk_out(Tile_X00_Y03_clk_out),
    .clk_pass_through(Tile_X00_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y03_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y02_config_out_config_addr),
    .config_config_data(Tile_X00_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y03_config_out_config_data),
    .config_out_read(Tile_X00_Y03_config_out_read),
    .config_out_write(Tile_X00_Y03_config_out_write),
    .config_read(Tile_X00_Y02_config_out_read),
    .config_write(Tile_X00_Y02_config_out_write),
    .flush(Tile_X00_Y02_flush_out),
    .flush_out(Tile_X00_Y03_flush_out),
    .hi(Tile_X00_Y03_hi),
    .lo(Tile_X00_Y03_lo),
    .read_config_data(Tile_X00_Y03_read_config_data),
    .read_config_data_in(Tile_X00_Y02_read_config_data),
    .reset(Tile_X00_Y02_reset_out),
    .reset_out(Tile_X00_Y03_reset_out),
    .stall(Tile_X00_Y02_stall_out),
    .stall_out(Tile_X00_Y03_stall_out),
    .tile_id(Tile_X00_Y03_tile_id)
);
wire [15:0] Tile_X00_Y04_tile_id;
assign Tile_X00_Y04_tile_id = {Tile_X00_Y04_lo[7],Tile_X00_Y04_lo[7],Tile_X00_Y04_lo[6],Tile_X00_Y04_lo[6],Tile_X00_Y04_lo[5],Tile_X00_Y04_lo[5],Tile_X00_Y04_lo[4],Tile_X00_Y04_lo[4],Tile_X00_Y04_lo[3],Tile_X00_Y04_lo[3],Tile_X00_Y04_lo[2],Tile_X00_Y04_lo[2],Tile_X00_Y04_lo[1],Tile_X00_Y04_hi[1],Tile_X00_Y04_lo[0],Tile_X00_Y04_lo[0]};
Tile_PE Tile_X00_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B17(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_EAST_SB_IN_B17_ready(Tile_X00_Y04_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_IN_B17_valid(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_IN_B1_ready(Tile_X00_Y04_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_IN_B1_valid(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B17(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_EAST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B17(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B17(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T0_SOUTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T0_SOUTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B17(Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B17(const_0_17_out),
    .SB_T0_WEST_SB_IN_B17_ready(Tile_X00_Y04_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T0_WEST_SB_IN_B1_ready(Tile_X00_Y04_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B17(Tile_X00_Y04_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T0_WEST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T0_WEST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B17(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_EAST_SB_IN_B17_ready(Tile_X00_Y04_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_IN_B17_valid(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_IN_B1_ready(Tile_X00_Y04_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_IN_B1_valid(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B17(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_EAST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B17(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B17(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T1_SOUTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T1_SOUTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B17(Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B17(const_0_17_out),
    .SB_T1_WEST_SB_IN_B17_ready(Tile_X00_Y04_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T1_WEST_SB_IN_B1_ready(Tile_X00_Y04_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B17(Tile_X00_Y04_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T1_WEST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T1_WEST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B17(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_EAST_SB_IN_B17_ready(Tile_X00_Y04_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_IN_B17_valid(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_IN_B1_ready(Tile_X00_Y04_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_IN_B1_valid(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B17(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_EAST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B17(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B17(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T2_SOUTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T2_SOUTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B17(Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B17(const_0_17_out),
    .SB_T2_WEST_SB_IN_B17_ready(Tile_X00_Y04_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T2_WEST_SB_IN_B1_ready(Tile_X00_Y04_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B17(Tile_X00_Y04_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T2_WEST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T2_WEST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B17(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_EAST_SB_IN_B17_ready(Tile_X00_Y04_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_IN_B17_valid(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_IN_B1_ready(Tile_X00_Y04_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_IN_B1_valid(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B17(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_EAST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B17(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B17(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T3_SOUTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T3_SOUTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B17(Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B17(const_0_17_out),
    .SB_T3_WEST_SB_IN_B17_ready(Tile_X00_Y04_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T3_WEST_SB_IN_B1_ready(Tile_X00_Y04_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B17(Tile_X00_Y04_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T3_WEST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T3_WEST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B17(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_EAST_SB_IN_B17_ready(Tile_X00_Y04_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_IN_B17_valid(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_IN_B1_ready(Tile_X00_Y04_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_IN_B1_valid(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B17(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_EAST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B17(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_IN_B17_valid(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_IN_B1_valid(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B17(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_OUT_B17_ready(Tile_X00_Y03_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_OUT_B1_ready(Tile_X00_Y03_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T4_SOUTH_SB_IN_B17_ready(Tile_X00_Y04_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T4_SOUTH_SB_IN_B1_ready(Tile_X00_Y04_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B17(Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B17(const_0_17_out),
    .SB_T4_WEST_SB_IN_B17_ready(Tile_X00_Y04_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T4_WEST_SB_IN_B1_ready(Tile_X00_Y04_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B17(Tile_X00_Y04_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_WEST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T4_WEST_SB_OUT_B17_valid(Tile_X00_Y04_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T4_WEST_SB_OUT_B1_valid(Tile_X00_Y04_SB_T4_WEST_SB_OUT_B1_valid),
    .clk(Tile_X00_Y03_clk_out),
    .clk_out(Tile_X00_Y04_clk_out),
    .clk_pass_through(Tile_X00_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y04_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y03_config_out_config_addr),
    .config_config_data(Tile_X00_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y04_config_out_config_data),
    .config_out_read(Tile_X00_Y04_config_out_read),
    .config_out_write(Tile_X00_Y04_config_out_write),
    .config_read(Tile_X00_Y03_config_out_read),
    .config_write(Tile_X00_Y03_config_out_write),
    .flush(Tile_X00_Y03_flush_out),
    .flush_out(Tile_X00_Y04_flush_out),
    .hi(Tile_X00_Y04_hi),
    .lo(Tile_X00_Y04_lo),
    .read_config_data(Tile_X00_Y04_read_config_data),
    .read_config_data_in(Tile_X00_Y03_read_config_data),
    .reset(Tile_X00_Y03_reset_out),
    .reset_out(Tile_X00_Y04_reset_out),
    .stall(Tile_X00_Y03_stall_out),
    .stall_out(Tile_X00_Y04_stall_out),
    .tile_id(Tile_X00_Y04_tile_id)
);
wire [31:0] Tile_X01_Y00_config_config_addr;
assign Tile_X01_Y00_config_config_addr = {PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[31],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[30],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[29],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[28],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[27],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[26],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[25],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[24],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[23],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[22],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[21],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[20],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[19],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[18],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[17],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[16],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[15],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[14],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[13],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[12],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[11],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[10],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[9],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[8],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[7],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[6],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[5],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[4],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[3],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[2],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[1],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[0]};
wire [31:0] Tile_X01_Y00_config_config_data;
assign Tile_X01_Y00_config_config_data = {PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[63],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[62],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[61],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[60],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[59],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[58],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[57],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[56],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[55],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[54],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[53],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[52],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[51],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[50],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[49],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[48],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[47],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[46],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[45],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[44],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[43],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[42],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[41],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[40],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[39],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[38],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[37],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[36],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[35],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[34],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[33],PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[32]};
wire [4:0] Tile_X01_Y00_io2f_17_ready;
assign Tile_X01_Y00_io2f_17_ready = {Tile_X01_Y01_SB_T4_NORTH_SB_IN_B17_ready,Tile_X01_Y01_SB_T3_NORTH_SB_IN_B17_ready,Tile_X01_Y01_SB_T2_NORTH_SB_IN_B17_ready,Tile_X01_Y01_SB_T1_NORTH_SB_IN_B17_ready,Tile_X01_Y01_SB_T0_NORTH_SB_IN_B17_ready};
wire [4:0] Tile_X01_Y00_io2f_1_ready;
assign Tile_X01_Y00_io2f_1_ready = {Tile_X01_Y01_SB_T4_NORTH_SB_IN_B1_ready,Tile_X01_Y01_SB_T3_NORTH_SB_IN_B1_ready,Tile_X01_Y01_SB_T2_NORTH_SB_IN_B1_ready,Tile_X01_Y01_SB_T1_NORTH_SB_IN_B1_ready,Tile_X01_Y01_SB_T0_NORTH_SB_IN_B1_ready};
wire [15:0] Tile_X01_Y00_tile_id;
assign Tile_X01_Y00_tile_id = {Tile_X01_Y00_lo[7],Tile_X01_Y00_lo[7],Tile_X01_Y00_lo[6],Tile_X01_Y00_lo[6],Tile_X01_Y00_lo[5],Tile_X01_Y00_lo[5],Tile_X01_Y00_lo[4],Tile_X01_Y00_hi[4],Tile_X01_Y00_lo[3],Tile_X01_Y00_lo[3],Tile_X01_Y00_lo[2],Tile_X01_Y00_lo[2],Tile_X01_Y00_lo[1],Tile_X01_Y00_lo[1],Tile_X01_Y00_lo[0],Tile_X01_Y00_lo[0]};
Tile_IOCoreReadyValid Tile_X01_Y00 (
    .clk(clk),
    .clk_out(Tile_X01_Y00_clk_out),
    .config_config_addr(Tile_X01_Y00_config_config_addr),
    .config_config_data(Tile_X01_Y00_config_config_data),
    .config_out_config_addr(Tile_X01_Y00_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y00_config_out_config_data),
    .config_out_read(Tile_X01_Y00_config_out_read),
    .config_out_write(Tile_X01_Y00_config_out_write),
    .config_read(PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[64]),
    .config_write(PipelineRegister_inst5$Register_inst0$reg_P66_inst0_out[65]),
    .f2io_1(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1),
    .f2io_17(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B17),
    .f2io_17_ready(Tile_X01_Y00_f2io_17_ready),
    .f2io_17_valid(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B17_valid),
    .f2io_1_ready(Tile_X01_Y00_f2io_1_ready),
    .f2io_1_valid(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1_valid),
    .flush(PipelineRegister_inst1$Register_inst0$reg_P1_inst0_out),
    .flush_out(Tile_X01_Y00_flush_out),
    .glb2io_1(glb2io_1_X01_Y00),
    .glb2io_17(glb2io_17_X01_Y00),
    .glb2io_17_ready(Tile_X01_Y00_glb2io_17_ready),
    .glb2io_17_valid(glb2io_17_X01_Y00_valid),
    .glb2io_1_ready(Tile_X01_Y00_glb2io_1_ready),
    .glb2io_1_valid(glb2io_1_X01_Y00_valid),
    .hi(Tile_X01_Y00_hi),
    .io2f_1(Tile_X01_Y00_io2f_1),
    .io2f_17(Tile_X01_Y00_io2f_17),
    .io2f_17_ready(Tile_X01_Y00_io2f_17_ready),
    .io2f_17_valid(Tile_X01_Y00_io2f_17_valid),
    .io2f_1_ready(Tile_X01_Y00_io2f_1_ready),
    .io2f_1_valid(Tile_X01_Y00_io2f_1_valid),
    .io2glb_1(Tile_X01_Y00_io2glb_1),
    .io2glb_17(Tile_X01_Y00_io2glb_17),
    .io2glb_17_ready(io2glb_17_X01_Y00_ready),
    .io2glb_17_valid(Tile_X01_Y00_io2glb_17_valid),
    .io2glb_1_ready(io2glb_1_X01_Y00_ready),
    .io2glb_1_valid(Tile_X01_Y00_io2glb_1_valid),
    .lo(Tile_X01_Y00_lo),
    .read_config_data(Tile_X01_Y00_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X01_Y00_reset_out),
    .stall(self_stall_out[1:1]),
    .stall_out(Tile_X01_Y00_stall_out),
    .tile_id(Tile_X01_Y00_tile_id)
);
wire [15:0] Tile_X01_Y01_tile_id;
assign Tile_X01_Y01_tile_id = {Tile_X01_Y01_lo[7],Tile_X01_Y01_lo[7],Tile_X01_Y01_lo[6],Tile_X01_Y01_lo[6],Tile_X01_Y01_lo[5],Tile_X01_Y01_lo[5],Tile_X01_Y01_lo[4],Tile_X01_Y01_hi[4],Tile_X01_Y01_lo[3],Tile_X01_Y01_lo[3],Tile_X01_Y01_lo[2],Tile_X01_Y01_lo[2],Tile_X01_Y01_lo[1],Tile_X01_Y01_lo[1],Tile_X01_Y01_lo[0],Tile_X01_Y01_hi[0]};
Tile_PE Tile_X01_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B17(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_EAST_SB_IN_B17_ready(Tile_X01_Y01_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_IN_B17_valid(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_IN_B1_ready(Tile_X01_Y01_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_IN_B1_valid(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B17(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_EAST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B17(Tile_X01_Y00_io2f_17),
    .SB_T0_NORTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_IN_B17_valid(Tile_X01_Y00_io2f_17_valid),
    .SB_T0_NORTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_IN_B1_valid(Tile_X01_Y00_io2f_1_valid),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B17(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_OUT_B17_ready(Tile_X01_Y00_f2io_17_ready),
    .SB_T0_NORTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_OUT_B1_ready(Tile_X01_Y00_f2io_1_ready),
    .SB_T0_NORTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B17(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B17(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B17(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_WEST_SB_IN_B17_ready(Tile_X01_Y01_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_IN_B17_valid(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_IN_B1_ready(Tile_X01_Y01_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_IN_B1_valid(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B17(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_WEST_SB_OUT_B17_ready(Tile_X00_Y01_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_OUT_B1_ready(Tile_X00_Y01_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B17(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_EAST_SB_IN_B17_ready(Tile_X01_Y01_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_IN_B17_valid(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_IN_B1_ready(Tile_X01_Y01_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_IN_B1_valid(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B17(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_EAST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B17(Tile_X01_Y00_io2f_17),
    .SB_T1_NORTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_IN_B17_valid(Tile_X01_Y00_io2f_17_valid),
    .SB_T1_NORTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_IN_B1_valid(Tile_X01_Y00_io2f_1_valid),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B17(Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T1_NORTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T1_NORTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B17(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B17(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B17(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_WEST_SB_IN_B17_ready(Tile_X01_Y01_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_IN_B17_valid(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_IN_B1_ready(Tile_X01_Y01_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_IN_B1_valid(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B17(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_WEST_SB_OUT_B17_ready(Tile_X00_Y01_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_OUT_B1_ready(Tile_X00_Y01_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B17(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_EAST_SB_IN_B17_ready(Tile_X01_Y01_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_IN_B17_valid(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_IN_B1_ready(Tile_X01_Y01_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_IN_B1_valid(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B17(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_EAST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B17(Tile_X01_Y00_io2f_17),
    .SB_T2_NORTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_IN_B17_valid(Tile_X01_Y00_io2f_17_valid),
    .SB_T2_NORTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_IN_B1_valid(Tile_X01_Y00_io2f_1_valid),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B17(Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T2_NORTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T2_NORTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B17(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B17(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B17(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_WEST_SB_IN_B17_ready(Tile_X01_Y01_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_IN_B17_valid(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_IN_B1_ready(Tile_X01_Y01_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_IN_B1_valid(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B17(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_WEST_SB_OUT_B17_ready(Tile_X00_Y01_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_OUT_B1_ready(Tile_X00_Y01_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B17(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_EAST_SB_IN_B17_ready(Tile_X01_Y01_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_IN_B17_valid(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_IN_B1_ready(Tile_X01_Y01_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_IN_B1_valid(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B17(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_EAST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B17(Tile_X01_Y00_io2f_17),
    .SB_T3_NORTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_IN_B17_valid(Tile_X01_Y00_io2f_17_valid),
    .SB_T3_NORTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_IN_B1_valid(Tile_X01_Y00_io2f_1_valid),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B17(Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T3_NORTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T3_NORTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B17(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B17(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B17(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_WEST_SB_IN_B17_ready(Tile_X01_Y01_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_IN_B17_valid(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_IN_B1_ready(Tile_X01_Y01_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_IN_B1_valid(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B17(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_WEST_SB_OUT_B17_ready(Tile_X00_Y01_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_OUT_B1_ready(Tile_X00_Y01_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B17(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_EAST_SB_IN_B17_ready(Tile_X01_Y01_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_IN_B17_valid(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_IN_B1_ready(Tile_X01_Y01_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_IN_B1_valid(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B17(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_EAST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B17(Tile_X01_Y00_io2f_17),
    .SB_T4_NORTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_IN_B17_valid(Tile_X01_Y00_io2f_17_valid),
    .SB_T4_NORTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_IN_B1_valid(Tile_X01_Y00_io2f_1_valid),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B17(Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T4_NORTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T4_NORTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B17(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_IN_B17_ready(Tile_X01_Y01_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_IN_B1_ready(Tile_X01_Y01_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B17(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B17(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_WEST_SB_IN_B17_ready(Tile_X01_Y01_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_IN_B17_valid(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_IN_B1_ready(Tile_X01_Y01_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_IN_B1_valid(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B17(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_WEST_SB_OUT_B17_ready(Tile_X00_Y01_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_OUT_B17_valid(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_OUT_B1_ready(Tile_X00_Y01_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_OUT_B1_valid(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B1_valid),
    .clk(Tile_X01_Y00_clk_out),
    .clk_out(Tile_X01_Y01_clk_out),
    .clk_pass_through(coreir_wrapInClock_inst1_out),
    .clk_pass_through_out_bot(Tile_X01_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y01_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y00_config_out_config_addr),
    .config_config_data(Tile_X01_Y00_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y01_config_out_config_data),
    .config_out_read(Tile_X01_Y01_config_out_read),
    .config_out_write(Tile_X01_Y01_config_out_write),
    .config_read(Tile_X01_Y00_config_out_read),
    .config_write(Tile_X01_Y00_config_out_write),
    .flush(Tile_X01_Y00_flush_out),
    .flush_out(Tile_X01_Y01_flush_out),
    .hi(Tile_X01_Y01_hi),
    .lo(Tile_X01_Y01_lo),
    .read_config_data(Tile_X01_Y01_read_config_data),
    .read_config_data_in(Tile_X01_Y00_read_config_data),
    .reset(Tile_X01_Y00_reset_out),
    .reset_out(Tile_X01_Y01_reset_out),
    .stall(Tile_X01_Y00_stall_out),
    .stall_out(Tile_X01_Y01_stall_out),
    .tile_id(Tile_X01_Y01_tile_id)
);
wire [15:0] Tile_X01_Y02_tile_id;
assign Tile_X01_Y02_tile_id = {Tile_X01_Y02_lo[7],Tile_X01_Y02_lo[7],Tile_X01_Y02_lo[6],Tile_X01_Y02_lo[6],Tile_X01_Y02_lo[5],Tile_X01_Y02_lo[5],Tile_X01_Y02_lo[4],Tile_X01_Y02_hi[4],Tile_X01_Y02_lo[3],Tile_X01_Y02_lo[3],Tile_X01_Y02_lo[2],Tile_X01_Y02_lo[2],Tile_X01_Y02_lo[1],Tile_X01_Y02_lo[1],Tile_X01_Y02_hi[1],Tile_X01_Y02_lo[0]};
Tile_PE Tile_X01_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B17(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_EAST_SB_IN_B17_ready(Tile_X01_Y02_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_IN_B17_valid(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_IN_B1_ready(Tile_X01_Y02_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_IN_B1_valid(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B17(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_EAST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B17(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_IN_B17_valid(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_IN_B1_valid(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B17(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_OUT_B17_ready(Tile_X01_Y01_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_OUT_B1_ready(Tile_X01_Y01_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B17(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B17(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B17(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_WEST_SB_IN_B17_ready(Tile_X01_Y02_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_IN_B17_valid(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_IN_B1_ready(Tile_X01_Y02_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_IN_B1_valid(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B17(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_WEST_SB_OUT_B17_ready(Tile_X00_Y02_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_OUT_B1_ready(Tile_X00_Y02_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B17(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_EAST_SB_IN_B17_ready(Tile_X01_Y02_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_IN_B17_valid(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_IN_B1_ready(Tile_X01_Y02_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_IN_B1_valid(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B17(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_EAST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B17(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_IN_B17_valid(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_IN_B1_valid(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B17(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_OUT_B17_ready(Tile_X01_Y01_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_OUT_B1_ready(Tile_X01_Y01_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B17(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B17(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B17(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_WEST_SB_IN_B17_ready(Tile_X01_Y02_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_IN_B17_valid(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_IN_B1_ready(Tile_X01_Y02_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_IN_B1_valid(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B17(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_WEST_SB_OUT_B17_ready(Tile_X00_Y02_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_OUT_B1_ready(Tile_X00_Y02_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B17(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_EAST_SB_IN_B17_ready(Tile_X01_Y02_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_IN_B17_valid(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_IN_B1_ready(Tile_X01_Y02_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_IN_B1_valid(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B17(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_EAST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B17(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_IN_B17_valid(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_IN_B1_valid(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B17(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_OUT_B17_ready(Tile_X01_Y01_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_OUT_B1_ready(Tile_X01_Y01_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B17(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B17(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B17(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_WEST_SB_IN_B17_ready(Tile_X01_Y02_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_IN_B17_valid(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_IN_B1_ready(Tile_X01_Y02_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_IN_B1_valid(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B17(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_WEST_SB_OUT_B17_ready(Tile_X00_Y02_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_OUT_B1_ready(Tile_X00_Y02_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B17(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_EAST_SB_IN_B17_ready(Tile_X01_Y02_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_IN_B17_valid(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_IN_B1_ready(Tile_X01_Y02_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_IN_B1_valid(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B17(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_EAST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B17(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_IN_B17_valid(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_IN_B1_valid(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B17(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_OUT_B17_ready(Tile_X01_Y01_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_OUT_B1_ready(Tile_X01_Y01_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B17(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B17(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B17(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_WEST_SB_IN_B17_ready(Tile_X01_Y02_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_IN_B17_valid(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_IN_B1_ready(Tile_X01_Y02_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_IN_B1_valid(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B17(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_WEST_SB_OUT_B17_ready(Tile_X00_Y02_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_OUT_B1_ready(Tile_X00_Y02_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B17(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_EAST_SB_IN_B17_ready(Tile_X01_Y02_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_IN_B17_valid(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_IN_B1_ready(Tile_X01_Y02_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_IN_B1_valid(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B17(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_EAST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B17(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_IN_B17_valid(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_IN_B1_valid(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B17(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_OUT_B17_ready(Tile_X01_Y01_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_OUT_B1_ready(Tile_X01_Y01_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B17(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_IN_B17_ready(Tile_X01_Y02_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_IN_B1_ready(Tile_X01_Y02_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B17(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B17(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_WEST_SB_IN_B17_ready(Tile_X01_Y02_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_IN_B17_valid(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_IN_B1_ready(Tile_X01_Y02_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_IN_B1_valid(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B17(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_WEST_SB_OUT_B17_ready(Tile_X00_Y02_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_OUT_B17_valid(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_OUT_B1_ready(Tile_X00_Y02_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_OUT_B1_valid(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B1_valid),
    .clk(Tile_X01_Y01_clk_out),
    .clk_out(Tile_X01_Y02_clk_out),
    .clk_pass_through(Tile_X01_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y02_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y01_config_out_config_addr),
    .config_config_data(Tile_X01_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y02_config_out_config_data),
    .config_out_read(Tile_X01_Y02_config_out_read),
    .config_out_write(Tile_X01_Y02_config_out_write),
    .config_read(Tile_X01_Y01_config_out_read),
    .config_write(Tile_X01_Y01_config_out_write),
    .flush(Tile_X01_Y01_flush_out),
    .flush_out(Tile_X01_Y02_flush_out),
    .hi(Tile_X01_Y02_hi),
    .lo(Tile_X01_Y02_lo),
    .read_config_data(Tile_X01_Y02_read_config_data),
    .read_config_data_in(Tile_X01_Y01_read_config_data),
    .reset(Tile_X01_Y01_reset_out),
    .reset_out(Tile_X01_Y02_reset_out),
    .stall(Tile_X01_Y01_stall_out),
    .stall_out(Tile_X01_Y02_stall_out),
    .tile_id(Tile_X01_Y02_tile_id)
);
wire [15:0] Tile_X01_Y03_tile_id;
assign Tile_X01_Y03_tile_id = {Tile_X01_Y03_lo[7],Tile_X01_Y03_lo[7],Tile_X01_Y03_lo[6],Tile_X01_Y03_lo[6],Tile_X01_Y03_lo[5],Tile_X01_Y03_lo[5],Tile_X01_Y03_lo[4],Tile_X01_Y03_hi[4],Tile_X01_Y03_lo[3],Tile_X01_Y03_lo[3],Tile_X01_Y03_lo[2],Tile_X01_Y03_lo[2],Tile_X01_Y03_lo[1],Tile_X01_Y03_lo[1],Tile_X01_Y03_hi[1],Tile_X01_Y03_hi[0]};
Tile_PE Tile_X01_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B17(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_EAST_SB_IN_B17_ready(Tile_X01_Y03_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_IN_B17_valid(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_IN_B1_ready(Tile_X01_Y03_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_IN_B1_valid(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B17(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_EAST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B17(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B17(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B17(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_IN_B17_valid(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_IN_B1_valid(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B17(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X01_Y04_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X01_Y04_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B17(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_WEST_SB_IN_B17_ready(Tile_X01_Y03_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_IN_B17_valid(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_IN_B1_ready(Tile_X01_Y03_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_IN_B1_valid(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B17(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_WEST_SB_OUT_B17_ready(Tile_X00_Y03_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_OUT_B1_ready(Tile_X00_Y03_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B17(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_EAST_SB_IN_B17_ready(Tile_X01_Y03_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_IN_B17_valid(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_IN_B1_ready(Tile_X01_Y03_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_IN_B1_valid(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B17(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_EAST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B17(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B17(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B17(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_IN_B17_valid(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_IN_B1_valid(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B17(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X01_Y04_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X01_Y04_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B17(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_WEST_SB_IN_B17_ready(Tile_X01_Y03_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_IN_B17_valid(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_IN_B1_ready(Tile_X01_Y03_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_IN_B1_valid(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B17(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_WEST_SB_OUT_B17_ready(Tile_X00_Y03_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_OUT_B1_ready(Tile_X00_Y03_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B17(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_EAST_SB_IN_B17_ready(Tile_X01_Y03_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_IN_B17_valid(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_IN_B1_ready(Tile_X01_Y03_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_IN_B1_valid(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B17(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_EAST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B17(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B17(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B17(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_IN_B17_valid(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_IN_B1_valid(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B17(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X01_Y04_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X01_Y04_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B17(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_WEST_SB_IN_B17_ready(Tile_X01_Y03_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_IN_B17_valid(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_IN_B1_ready(Tile_X01_Y03_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_IN_B1_valid(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B17(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_WEST_SB_OUT_B17_ready(Tile_X00_Y03_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_OUT_B1_ready(Tile_X00_Y03_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B17(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_EAST_SB_IN_B17_ready(Tile_X01_Y03_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_IN_B17_valid(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_IN_B1_ready(Tile_X01_Y03_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_IN_B1_valid(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B17(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_EAST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B17(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B17(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B17(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_IN_B17_valid(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_IN_B1_valid(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B17(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X01_Y04_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X01_Y04_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B17(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_WEST_SB_IN_B17_ready(Tile_X01_Y03_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_IN_B17_valid(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_IN_B1_ready(Tile_X01_Y03_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_IN_B1_valid(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B17(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_WEST_SB_OUT_B17_ready(Tile_X00_Y03_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_OUT_B1_ready(Tile_X00_Y03_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B17(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_EAST_SB_IN_B17_ready(Tile_X01_Y03_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_IN_B17_valid(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_IN_B1_ready(Tile_X01_Y03_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_IN_B1_valid(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B17(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_EAST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B17(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_IN_B17_valid(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_IN_B1_valid(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B17(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_OUT_B17_ready(Tile_X01_Y02_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_OUT_B1_ready(Tile_X01_Y02_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B17(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_IN_B17_ready(Tile_X01_Y03_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_IN_B17_valid(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_IN_B1_ready(Tile_X01_Y03_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_IN_B1_valid(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B17(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X01_Y04_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X01_Y04_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B17(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_WEST_SB_IN_B17_ready(Tile_X01_Y03_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_IN_B17_valid(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_IN_B1_ready(Tile_X01_Y03_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_IN_B1_valid(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B17(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_WEST_SB_OUT_B17_ready(Tile_X00_Y03_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_OUT_B17_valid(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_OUT_B1_ready(Tile_X00_Y03_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_OUT_B1_valid(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B1_valid),
    .clk(Tile_X01_Y02_clk_out),
    .clk_out(Tile_X01_Y03_clk_out),
    .clk_pass_through(Tile_X01_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y03_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y02_config_out_config_addr),
    .config_config_data(Tile_X01_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y03_config_out_config_data),
    .config_out_read(Tile_X01_Y03_config_out_read),
    .config_out_write(Tile_X01_Y03_config_out_write),
    .config_read(Tile_X01_Y02_config_out_read),
    .config_write(Tile_X01_Y02_config_out_write),
    .flush(Tile_X01_Y02_flush_out),
    .flush_out(Tile_X01_Y03_flush_out),
    .hi(Tile_X01_Y03_hi),
    .lo(Tile_X01_Y03_lo),
    .read_config_data(Tile_X01_Y03_read_config_data),
    .read_config_data_in(Tile_X01_Y02_read_config_data),
    .reset(Tile_X01_Y02_reset_out),
    .reset_out(Tile_X01_Y03_reset_out),
    .stall(Tile_X01_Y02_stall_out),
    .stall_out(Tile_X01_Y03_stall_out),
    .tile_id(Tile_X01_Y03_tile_id)
);
wire [15:0] Tile_X01_Y04_tile_id;
assign Tile_X01_Y04_tile_id = {Tile_X01_Y04_lo[7],Tile_X01_Y04_lo[7],Tile_X01_Y04_lo[6],Tile_X01_Y04_lo[6],Tile_X01_Y04_lo[5],Tile_X01_Y04_lo[5],Tile_X01_Y04_lo[4],Tile_X01_Y04_hi[4],Tile_X01_Y04_lo[3],Tile_X01_Y04_lo[3],Tile_X01_Y04_lo[2],Tile_X01_Y04_lo[2],Tile_X01_Y04_lo[1],Tile_X01_Y04_hi[1],Tile_X01_Y04_lo[0],Tile_X01_Y04_lo[0]};
Tile_PE Tile_X01_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B17(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_EAST_SB_IN_B17_ready(Tile_X01_Y04_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_IN_B17_valid(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_IN_B1_ready(Tile_X01_Y04_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_IN_B1_valid(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B17(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_EAST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B17(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B17(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T0_SOUTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T0_SOUTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B17(Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B17(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_WEST_SB_IN_B17_ready(Tile_X01_Y04_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_IN_B17_valid(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_IN_B1_ready(Tile_X01_Y04_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_IN_B1_valid(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B17(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_WEST_SB_OUT_B17_ready(Tile_X00_Y04_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_OUT_B1_ready(Tile_X00_Y04_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B17(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_EAST_SB_IN_B17_ready(Tile_X01_Y04_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_IN_B17_valid(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_IN_B1_ready(Tile_X01_Y04_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_IN_B1_valid(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B17(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_EAST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B17(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B17(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T1_SOUTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T1_SOUTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B17(Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B17(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_WEST_SB_IN_B17_ready(Tile_X01_Y04_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_IN_B17_valid(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_IN_B1_ready(Tile_X01_Y04_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_IN_B1_valid(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B17(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_WEST_SB_OUT_B17_ready(Tile_X00_Y04_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_OUT_B1_ready(Tile_X00_Y04_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B17(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_EAST_SB_IN_B17_ready(Tile_X01_Y04_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_IN_B17_valid(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_IN_B1_ready(Tile_X01_Y04_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_IN_B1_valid(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B17(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_EAST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B17(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B17(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T2_SOUTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T2_SOUTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B17(Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B17(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_WEST_SB_IN_B17_ready(Tile_X01_Y04_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_IN_B17_valid(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_IN_B1_ready(Tile_X01_Y04_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_IN_B1_valid(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B17(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_WEST_SB_OUT_B17_ready(Tile_X00_Y04_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_OUT_B1_ready(Tile_X00_Y04_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B17(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_EAST_SB_IN_B17_ready(Tile_X01_Y04_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_IN_B17_valid(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_IN_B1_ready(Tile_X01_Y04_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_IN_B1_valid(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B17(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_EAST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B17(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B17(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T3_SOUTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T3_SOUTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B17(Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B17(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_WEST_SB_IN_B17_ready(Tile_X01_Y04_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_IN_B17_valid(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_IN_B1_ready(Tile_X01_Y04_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_IN_B1_valid(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B17(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_WEST_SB_OUT_B17_ready(Tile_X00_Y04_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_OUT_B1_ready(Tile_X00_Y04_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B17(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_EAST_SB_IN_B17_ready(Tile_X01_Y04_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_IN_B17_valid(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_IN_B1_ready(Tile_X01_Y04_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_IN_B1_valid(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B17(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_EAST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B17(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_IN_B17_valid(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_IN_B1_valid(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B17(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_OUT_B17_ready(Tile_X01_Y03_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_OUT_B1_ready(Tile_X01_Y03_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T4_SOUTH_SB_IN_B17_ready(Tile_X01_Y04_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T4_SOUTH_SB_IN_B1_ready(Tile_X01_Y04_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B17(Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B17(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_WEST_SB_IN_B17_ready(Tile_X01_Y04_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_IN_B17_valid(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_IN_B1_ready(Tile_X01_Y04_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_IN_B1_valid(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B17(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_WEST_SB_OUT_B17_ready(Tile_X00_Y04_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_OUT_B17_valid(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_OUT_B1_ready(Tile_X00_Y04_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_OUT_B1_valid(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B1_valid),
    .clk(Tile_X01_Y03_clk_out),
    .clk_out(Tile_X01_Y04_clk_out),
    .clk_pass_through(Tile_X01_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y04_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y03_config_out_config_addr),
    .config_config_data(Tile_X01_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y04_config_out_config_data),
    .config_out_read(Tile_X01_Y04_config_out_read),
    .config_out_write(Tile_X01_Y04_config_out_write),
    .config_read(Tile_X01_Y03_config_out_read),
    .config_write(Tile_X01_Y03_config_out_write),
    .flush(Tile_X01_Y03_flush_out),
    .flush_out(Tile_X01_Y04_flush_out),
    .hi(Tile_X01_Y04_hi),
    .lo(Tile_X01_Y04_lo),
    .read_config_data(Tile_X01_Y04_read_config_data),
    .read_config_data_in(Tile_X01_Y03_read_config_data),
    .reset(Tile_X01_Y03_reset_out),
    .reset_out(Tile_X01_Y04_reset_out),
    .stall(Tile_X01_Y03_stall_out),
    .stall_out(Tile_X01_Y04_stall_out),
    .tile_id(Tile_X01_Y04_tile_id)
);
wire [31:0] Tile_X02_Y00_config_config_addr;
assign Tile_X02_Y00_config_config_addr = {PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[31],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[30],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[29],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[28],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[27],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[26],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[25],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[24],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[23],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[22],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[21],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[20],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[19],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[18],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[17],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[16],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[15],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[14],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[13],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[12],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[11],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[10],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[9],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[8],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[7],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[6],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[5],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[4],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[3],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[2],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[1],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[0]};
wire [31:0] Tile_X02_Y00_config_config_data;
assign Tile_X02_Y00_config_config_data = {PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[63],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[62],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[61],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[60],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[59],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[58],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[57],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[56],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[55],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[54],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[53],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[52],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[51],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[50],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[49],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[48],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[47],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[46],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[45],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[44],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[43],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[42],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[41],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[40],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[39],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[38],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[37],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[36],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[35],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[34],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[33],PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[32]};
wire [4:0] Tile_X02_Y00_io2f_17_ready;
assign Tile_X02_Y00_io2f_17_ready = {Tile_X02_Y01_SB_T4_NORTH_SB_IN_B17_ready,Tile_X02_Y01_SB_T3_NORTH_SB_IN_B17_ready,Tile_X02_Y01_SB_T2_NORTH_SB_IN_B17_ready,Tile_X02_Y01_SB_T1_NORTH_SB_IN_B17_ready,Tile_X02_Y01_SB_T0_NORTH_SB_IN_B17_ready};
wire [4:0] Tile_X02_Y00_io2f_1_ready;
assign Tile_X02_Y00_io2f_1_ready = {Tile_X02_Y01_SB_T4_NORTH_SB_IN_B1_ready,Tile_X02_Y01_SB_T3_NORTH_SB_IN_B1_ready,Tile_X02_Y01_SB_T2_NORTH_SB_IN_B1_ready,Tile_X02_Y01_SB_T1_NORTH_SB_IN_B1_ready,Tile_X02_Y01_SB_T0_NORTH_SB_IN_B1_ready};
wire [15:0] Tile_X02_Y00_tile_id;
assign Tile_X02_Y00_tile_id = {Tile_X02_Y00_lo[7],Tile_X02_Y00_lo[7],Tile_X02_Y00_lo[6],Tile_X02_Y00_lo[6],Tile_X02_Y00_lo[5],Tile_X02_Y00_lo[5],Tile_X02_Y00_hi[5],Tile_X02_Y00_lo[4],Tile_X02_Y00_lo[3],Tile_X02_Y00_lo[3],Tile_X02_Y00_lo[2],Tile_X02_Y00_lo[2],Tile_X02_Y00_lo[1],Tile_X02_Y00_lo[1],Tile_X02_Y00_lo[0],Tile_X02_Y00_lo[0]};
Tile_IOCoreReadyValid Tile_X02_Y00 (
    .clk(clk),
    .clk_out(Tile_X02_Y00_clk_out),
    .config_config_addr(Tile_X02_Y00_config_config_addr),
    .config_config_data(Tile_X02_Y00_config_config_data),
    .config_out_config_addr(Tile_X02_Y00_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y00_config_out_config_data),
    .config_out_read(Tile_X02_Y00_config_out_read),
    .config_out_write(Tile_X02_Y00_config_out_write),
    .config_read(PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[64]),
    .config_write(PipelineRegister_inst6$Register_inst0$reg_P66_inst0_out[65]),
    .f2io_1(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1),
    .f2io_17(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B17),
    .f2io_17_ready(Tile_X02_Y00_f2io_17_ready),
    .f2io_17_valid(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B17_valid),
    .f2io_1_ready(Tile_X02_Y00_f2io_1_ready),
    .f2io_1_valid(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1_valid),
    .flush(PipelineRegister_inst2$Register_inst0$reg_P1_inst0_out),
    .flush_out(Tile_X02_Y00_flush_out),
    .glb2io_1(glb2io_1_X02_Y00),
    .glb2io_17(glb2io_17_X02_Y00),
    .glb2io_17_ready(Tile_X02_Y00_glb2io_17_ready),
    .glb2io_17_valid(glb2io_17_X02_Y00_valid),
    .glb2io_1_ready(Tile_X02_Y00_glb2io_1_ready),
    .glb2io_1_valid(glb2io_1_X02_Y00_valid),
    .hi(Tile_X02_Y00_hi),
    .io2f_1(Tile_X02_Y00_io2f_1),
    .io2f_17(Tile_X02_Y00_io2f_17),
    .io2f_17_ready(Tile_X02_Y00_io2f_17_ready),
    .io2f_17_valid(Tile_X02_Y00_io2f_17_valid),
    .io2f_1_ready(Tile_X02_Y00_io2f_1_ready),
    .io2f_1_valid(Tile_X02_Y00_io2f_1_valid),
    .io2glb_1(Tile_X02_Y00_io2glb_1),
    .io2glb_17(Tile_X02_Y00_io2glb_17),
    .io2glb_17_ready(io2glb_17_X02_Y00_ready),
    .io2glb_17_valid(Tile_X02_Y00_io2glb_17_valid),
    .io2glb_1_ready(io2glb_1_X02_Y00_ready),
    .io2glb_1_valid(Tile_X02_Y00_io2glb_1_valid),
    .lo(Tile_X02_Y00_lo),
    .read_config_data(Tile_X02_Y00_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X02_Y00_reset_out),
    .stall(self_stall_out[2:2]),
    .stall_out(Tile_X02_Y00_stall_out),
    .tile_id(Tile_X02_Y00_tile_id)
);
wire [15:0] Tile_X02_Y01_tile_id;
assign Tile_X02_Y01_tile_id = {Tile_X02_Y01_lo[7],Tile_X02_Y01_lo[7],Tile_X02_Y01_lo[6],Tile_X02_Y01_lo[6],Tile_X02_Y01_lo[5],Tile_X02_Y01_lo[5],Tile_X02_Y01_hi[5],Tile_X02_Y01_lo[4],Tile_X02_Y01_lo[3],Tile_X02_Y01_lo[3],Tile_X02_Y01_lo[2],Tile_X02_Y01_lo[2],Tile_X02_Y01_lo[1],Tile_X02_Y01_lo[1],Tile_X02_Y01_lo[0],Tile_X02_Y01_hi[0]};
Tile_PE Tile_X02_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B17(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_EAST_SB_IN_B17_ready(Tile_X02_Y01_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_IN_B17_valid(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_IN_B1_ready(Tile_X02_Y01_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_IN_B1_valid(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B17(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_EAST_SB_OUT_B17_ready(Tile_X03_Y01_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_OUT_B1_ready(Tile_X03_Y01_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B17(Tile_X02_Y00_io2f_17),
    .SB_T0_NORTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_IN_B17_valid(Tile_X02_Y00_io2f_17_valid),
    .SB_T0_NORTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_IN_B1_valid(Tile_X02_Y00_io2f_1_valid),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B17(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_OUT_B17_ready(Tile_X02_Y00_f2io_17_ready),
    .SB_T0_NORTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_OUT_B1_ready(Tile_X02_Y00_f2io_1_ready),
    .SB_T0_NORTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B17(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B17(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B17(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_WEST_SB_IN_B17_ready(Tile_X02_Y01_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_IN_B17_valid(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_IN_B1_ready(Tile_X02_Y01_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_IN_B1_valid(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B17(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_WEST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B17(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_EAST_SB_IN_B17_ready(Tile_X02_Y01_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_IN_B17_valid(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_IN_B1_ready(Tile_X02_Y01_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_IN_B1_valid(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B17(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_EAST_SB_OUT_B17_ready(Tile_X03_Y01_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_OUT_B1_ready(Tile_X03_Y01_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B17(Tile_X02_Y00_io2f_17),
    .SB_T1_NORTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_IN_B17_valid(Tile_X02_Y00_io2f_17_valid),
    .SB_T1_NORTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_IN_B1_valid(Tile_X02_Y00_io2f_1_valid),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B17(Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T1_NORTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T1_NORTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B17(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B17(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B17(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_WEST_SB_IN_B17_ready(Tile_X02_Y01_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_IN_B17_valid(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_IN_B1_ready(Tile_X02_Y01_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_IN_B1_valid(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B17(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_WEST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B17(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_EAST_SB_IN_B17_ready(Tile_X02_Y01_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_IN_B17_valid(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_IN_B1_ready(Tile_X02_Y01_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_IN_B1_valid(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B17(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_EAST_SB_OUT_B17_ready(Tile_X03_Y01_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_OUT_B1_ready(Tile_X03_Y01_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B17(Tile_X02_Y00_io2f_17),
    .SB_T2_NORTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_IN_B17_valid(Tile_X02_Y00_io2f_17_valid),
    .SB_T2_NORTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_IN_B1_valid(Tile_X02_Y00_io2f_1_valid),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B17(Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T2_NORTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T2_NORTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B17(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B17(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B17(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_WEST_SB_IN_B17_ready(Tile_X02_Y01_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_IN_B17_valid(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_IN_B1_ready(Tile_X02_Y01_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_IN_B1_valid(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B17(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_WEST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B17(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_EAST_SB_IN_B17_ready(Tile_X02_Y01_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_IN_B17_valid(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_IN_B1_ready(Tile_X02_Y01_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_IN_B1_valid(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B17(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_EAST_SB_OUT_B17_ready(Tile_X03_Y01_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_OUT_B1_ready(Tile_X03_Y01_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B17(Tile_X02_Y00_io2f_17),
    .SB_T3_NORTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_IN_B17_valid(Tile_X02_Y00_io2f_17_valid),
    .SB_T3_NORTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_IN_B1_valid(Tile_X02_Y00_io2f_1_valid),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B17(Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T3_NORTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T3_NORTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B17(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B17(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B17(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_WEST_SB_IN_B17_ready(Tile_X02_Y01_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_IN_B17_valid(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_IN_B1_ready(Tile_X02_Y01_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_IN_B1_valid(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B17(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_WEST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B17(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_EAST_SB_IN_B17_ready(Tile_X02_Y01_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_IN_B17_valid(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_IN_B1_ready(Tile_X02_Y01_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_IN_B1_valid(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B17(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_EAST_SB_OUT_B17_ready(Tile_X03_Y01_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_OUT_B1_ready(Tile_X03_Y01_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B17(Tile_X02_Y00_io2f_17),
    .SB_T4_NORTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_IN_B17_valid(Tile_X02_Y00_io2f_17_valid),
    .SB_T4_NORTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_IN_B1_valid(Tile_X02_Y00_io2f_1_valid),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B17(Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T4_NORTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T4_NORTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B17(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_IN_B17_ready(Tile_X02_Y01_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_IN_B1_ready(Tile_X02_Y01_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B17(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B17(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_WEST_SB_IN_B17_ready(Tile_X02_Y01_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_IN_B17_valid(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_IN_B1_ready(Tile_X02_Y01_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_IN_B1_valid(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B17(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_WEST_SB_OUT_B17_ready(Tile_X01_Y01_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_OUT_B17_valid(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_OUT_B1_ready(Tile_X01_Y01_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_OUT_B1_valid(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B1_valid),
    .clk(Tile_X02_Y00_clk_out),
    .clk_out(Tile_X02_Y01_clk_out),
    .clk_pass_through(coreir_wrapInClock_inst2_out),
    .clk_pass_through_out_bot(Tile_X02_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y01_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y00_config_out_config_addr),
    .config_config_data(Tile_X02_Y00_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y01_config_out_config_data),
    .config_out_read(Tile_X02_Y01_config_out_read),
    .config_out_write(Tile_X02_Y01_config_out_write),
    .config_read(Tile_X02_Y00_config_out_read),
    .config_write(Tile_X02_Y00_config_out_write),
    .flush(Tile_X02_Y00_flush_out),
    .flush_out(Tile_X02_Y01_flush_out),
    .hi(Tile_X02_Y01_hi),
    .lo(Tile_X02_Y01_lo),
    .read_config_data(Tile_X02_Y01_read_config_data),
    .read_config_data_in(Tile_X02_Y00_read_config_data),
    .reset(Tile_X02_Y00_reset_out),
    .reset_out(Tile_X02_Y01_reset_out),
    .stall(Tile_X02_Y00_stall_out),
    .stall_out(Tile_X02_Y01_stall_out),
    .tile_id(Tile_X02_Y01_tile_id)
);
wire [15:0] Tile_X02_Y02_tile_id;
assign Tile_X02_Y02_tile_id = {Tile_X02_Y02_lo[7],Tile_X02_Y02_lo[7],Tile_X02_Y02_lo[6],Tile_X02_Y02_lo[6],Tile_X02_Y02_lo[5],Tile_X02_Y02_lo[5],Tile_X02_Y02_hi[5],Tile_X02_Y02_lo[4],Tile_X02_Y02_lo[3],Tile_X02_Y02_lo[3],Tile_X02_Y02_lo[2],Tile_X02_Y02_lo[2],Tile_X02_Y02_lo[1],Tile_X02_Y02_lo[1],Tile_X02_Y02_hi[1],Tile_X02_Y02_lo[0]};
Tile_PE Tile_X02_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B17(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_EAST_SB_IN_B17_ready(Tile_X02_Y02_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_IN_B17_valid(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_IN_B1_ready(Tile_X02_Y02_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_IN_B1_valid(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B17(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_EAST_SB_OUT_B17_ready(Tile_X03_Y02_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_OUT_B1_ready(Tile_X03_Y02_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B17(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_IN_B17_valid(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_IN_B1_valid(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B17(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_OUT_B17_ready(Tile_X02_Y01_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_OUT_B1_ready(Tile_X02_Y01_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B17(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B17(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B17(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_WEST_SB_IN_B17_ready(Tile_X02_Y02_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_IN_B17_valid(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_IN_B1_ready(Tile_X02_Y02_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_IN_B1_valid(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B17(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_WEST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B17(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_EAST_SB_IN_B17_ready(Tile_X02_Y02_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_IN_B17_valid(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_IN_B1_ready(Tile_X02_Y02_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_IN_B1_valid(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B17(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_EAST_SB_OUT_B17_ready(Tile_X03_Y02_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_OUT_B1_ready(Tile_X03_Y02_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B17(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_IN_B17_valid(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_IN_B1_valid(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B17(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_OUT_B17_ready(Tile_X02_Y01_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_OUT_B1_ready(Tile_X02_Y01_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B17(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B17(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B17(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_WEST_SB_IN_B17_ready(Tile_X02_Y02_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_IN_B17_valid(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_IN_B1_ready(Tile_X02_Y02_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_IN_B1_valid(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B17(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_WEST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B17(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_EAST_SB_IN_B17_ready(Tile_X02_Y02_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_IN_B17_valid(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_IN_B1_ready(Tile_X02_Y02_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_IN_B1_valid(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B17(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_EAST_SB_OUT_B17_ready(Tile_X03_Y02_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_OUT_B1_ready(Tile_X03_Y02_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B17(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_IN_B17_valid(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_IN_B1_valid(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B17(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_OUT_B17_ready(Tile_X02_Y01_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_OUT_B1_ready(Tile_X02_Y01_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B17(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B17(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B17(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_WEST_SB_IN_B17_ready(Tile_X02_Y02_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_IN_B17_valid(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_IN_B1_ready(Tile_X02_Y02_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_IN_B1_valid(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B17(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_WEST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B17(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_EAST_SB_IN_B17_ready(Tile_X02_Y02_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_IN_B17_valid(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_IN_B1_ready(Tile_X02_Y02_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_IN_B1_valid(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B17(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_EAST_SB_OUT_B17_ready(Tile_X03_Y02_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_OUT_B1_ready(Tile_X03_Y02_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B17(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_IN_B17_valid(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_IN_B1_valid(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B17(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_OUT_B17_ready(Tile_X02_Y01_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_OUT_B1_ready(Tile_X02_Y01_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B17(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B17(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B17(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_WEST_SB_IN_B17_ready(Tile_X02_Y02_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_IN_B17_valid(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_IN_B1_ready(Tile_X02_Y02_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_IN_B1_valid(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B17(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_WEST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B17(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_EAST_SB_IN_B17_ready(Tile_X02_Y02_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_IN_B17_valid(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_IN_B1_ready(Tile_X02_Y02_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_IN_B1_valid(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B17(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_EAST_SB_OUT_B17_ready(Tile_X03_Y02_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_OUT_B1_ready(Tile_X03_Y02_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B17(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_IN_B17_valid(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_IN_B1_valid(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B17(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_OUT_B17_ready(Tile_X02_Y01_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_OUT_B1_ready(Tile_X02_Y01_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B17(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_IN_B17_ready(Tile_X02_Y02_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_IN_B1_ready(Tile_X02_Y02_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B17(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B17(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_WEST_SB_IN_B17_ready(Tile_X02_Y02_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_IN_B17_valid(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_IN_B1_ready(Tile_X02_Y02_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_IN_B1_valid(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B17(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_WEST_SB_OUT_B17_ready(Tile_X01_Y02_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_OUT_B17_valid(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_OUT_B1_ready(Tile_X01_Y02_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_OUT_B1_valid(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B1_valid),
    .clk(Tile_X02_Y01_clk_out),
    .clk_out(Tile_X02_Y02_clk_out),
    .clk_pass_through(Tile_X02_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y02_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y01_config_out_config_addr),
    .config_config_data(Tile_X02_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y02_config_out_config_data),
    .config_out_read(Tile_X02_Y02_config_out_read),
    .config_out_write(Tile_X02_Y02_config_out_write),
    .config_read(Tile_X02_Y01_config_out_read),
    .config_write(Tile_X02_Y01_config_out_write),
    .flush(Tile_X02_Y01_flush_out),
    .flush_out(Tile_X02_Y02_flush_out),
    .hi(Tile_X02_Y02_hi),
    .lo(Tile_X02_Y02_lo),
    .read_config_data(Tile_X02_Y02_read_config_data),
    .read_config_data_in(Tile_X02_Y01_read_config_data),
    .reset(Tile_X02_Y01_reset_out),
    .reset_out(Tile_X02_Y02_reset_out),
    .stall(Tile_X02_Y01_stall_out),
    .stall_out(Tile_X02_Y02_stall_out),
    .tile_id(Tile_X02_Y02_tile_id)
);
wire [15:0] Tile_X02_Y03_tile_id;
assign Tile_X02_Y03_tile_id = {Tile_X02_Y03_lo[7],Tile_X02_Y03_lo[7],Tile_X02_Y03_lo[6],Tile_X02_Y03_lo[6],Tile_X02_Y03_lo[5],Tile_X02_Y03_lo[5],Tile_X02_Y03_hi[5],Tile_X02_Y03_lo[4],Tile_X02_Y03_lo[3],Tile_X02_Y03_lo[3],Tile_X02_Y03_lo[2],Tile_X02_Y03_lo[2],Tile_X02_Y03_lo[1],Tile_X02_Y03_lo[1],Tile_X02_Y03_hi[1],Tile_X02_Y03_hi[0]};
Tile_PE Tile_X02_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B17(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_EAST_SB_IN_B17_ready(Tile_X02_Y03_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_IN_B17_valid(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_IN_B1_ready(Tile_X02_Y03_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_IN_B1_valid(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B17(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_EAST_SB_OUT_B17_ready(Tile_X03_Y03_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_OUT_B1_ready(Tile_X03_Y03_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B17(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B17(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B17(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_IN_B17_valid(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_IN_B1_valid(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B17(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X02_Y04_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X02_Y04_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B17(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_WEST_SB_IN_B17_ready(Tile_X02_Y03_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_IN_B17_valid(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_IN_B1_ready(Tile_X02_Y03_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_IN_B1_valid(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B17(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_WEST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B17(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_EAST_SB_IN_B17_ready(Tile_X02_Y03_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_IN_B17_valid(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_IN_B1_ready(Tile_X02_Y03_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_IN_B1_valid(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B17(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_EAST_SB_OUT_B17_ready(Tile_X03_Y03_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_OUT_B1_ready(Tile_X03_Y03_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B17(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B17(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B17(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_IN_B17_valid(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_IN_B1_valid(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B17(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X02_Y04_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X02_Y04_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B17(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_WEST_SB_IN_B17_ready(Tile_X02_Y03_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_IN_B17_valid(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_IN_B1_ready(Tile_X02_Y03_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_IN_B1_valid(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B17(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_WEST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B17(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_EAST_SB_IN_B17_ready(Tile_X02_Y03_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_IN_B17_valid(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_IN_B1_ready(Tile_X02_Y03_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_IN_B1_valid(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B17(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_EAST_SB_OUT_B17_ready(Tile_X03_Y03_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_OUT_B1_ready(Tile_X03_Y03_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B17(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B17(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B17(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_IN_B17_valid(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_IN_B1_valid(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B17(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X02_Y04_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X02_Y04_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B17(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_WEST_SB_IN_B17_ready(Tile_X02_Y03_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_IN_B17_valid(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_IN_B1_ready(Tile_X02_Y03_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_IN_B1_valid(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B17(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_WEST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B17(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_EAST_SB_IN_B17_ready(Tile_X02_Y03_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_IN_B17_valid(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_IN_B1_ready(Tile_X02_Y03_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_IN_B1_valid(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B17(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_EAST_SB_OUT_B17_ready(Tile_X03_Y03_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_OUT_B1_ready(Tile_X03_Y03_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B17(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B17(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B17(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_IN_B17_valid(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_IN_B1_valid(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B17(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X02_Y04_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X02_Y04_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B17(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_WEST_SB_IN_B17_ready(Tile_X02_Y03_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_IN_B17_valid(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_IN_B1_ready(Tile_X02_Y03_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_IN_B1_valid(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B17(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_WEST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B17(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_EAST_SB_IN_B17_ready(Tile_X02_Y03_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_IN_B17_valid(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_IN_B1_ready(Tile_X02_Y03_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_IN_B1_valid(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B17(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_EAST_SB_OUT_B17_ready(Tile_X03_Y03_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_OUT_B1_ready(Tile_X03_Y03_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B17(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_IN_B17_valid(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_IN_B1_valid(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B17(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_OUT_B17_ready(Tile_X02_Y02_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_OUT_B1_ready(Tile_X02_Y02_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B17(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_IN_B17_ready(Tile_X02_Y03_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_IN_B17_valid(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_IN_B1_ready(Tile_X02_Y03_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_IN_B1_valid(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B17(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X02_Y04_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X02_Y04_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B17(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_WEST_SB_IN_B17_ready(Tile_X02_Y03_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_IN_B17_valid(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_IN_B1_ready(Tile_X02_Y03_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_IN_B1_valid(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B17(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_WEST_SB_OUT_B17_ready(Tile_X01_Y03_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_OUT_B17_valid(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_OUT_B1_ready(Tile_X01_Y03_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_OUT_B1_valid(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B1_valid),
    .clk(Tile_X02_Y02_clk_out),
    .clk_out(Tile_X02_Y03_clk_out),
    .clk_pass_through(Tile_X02_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y03_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y02_config_out_config_addr),
    .config_config_data(Tile_X02_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y03_config_out_config_data),
    .config_out_read(Tile_X02_Y03_config_out_read),
    .config_out_write(Tile_X02_Y03_config_out_write),
    .config_read(Tile_X02_Y02_config_out_read),
    .config_write(Tile_X02_Y02_config_out_write),
    .flush(Tile_X02_Y02_flush_out),
    .flush_out(Tile_X02_Y03_flush_out),
    .hi(Tile_X02_Y03_hi),
    .lo(Tile_X02_Y03_lo),
    .read_config_data(Tile_X02_Y03_read_config_data),
    .read_config_data_in(Tile_X02_Y02_read_config_data),
    .reset(Tile_X02_Y02_reset_out),
    .reset_out(Tile_X02_Y03_reset_out),
    .stall(Tile_X02_Y02_stall_out),
    .stall_out(Tile_X02_Y03_stall_out),
    .tile_id(Tile_X02_Y03_tile_id)
);
wire [15:0] Tile_X02_Y04_tile_id;
assign Tile_X02_Y04_tile_id = {Tile_X02_Y04_lo[7],Tile_X02_Y04_lo[7],Tile_X02_Y04_lo[6],Tile_X02_Y04_lo[6],Tile_X02_Y04_lo[5],Tile_X02_Y04_lo[5],Tile_X02_Y04_hi[5],Tile_X02_Y04_lo[4],Tile_X02_Y04_lo[3],Tile_X02_Y04_lo[3],Tile_X02_Y04_lo[2],Tile_X02_Y04_lo[2],Tile_X02_Y04_lo[1],Tile_X02_Y04_hi[1],Tile_X02_Y04_lo[0],Tile_X02_Y04_lo[0]};
Tile_PE Tile_X02_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B17(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_EAST_SB_IN_B17_ready(Tile_X02_Y04_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_IN_B17_valid(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_IN_B1_ready(Tile_X02_Y04_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_IN_B1_valid(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B17(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_EAST_SB_OUT_B17_ready(Tile_X03_Y04_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_OUT_B1_ready(Tile_X03_Y04_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B17(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B17(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T0_SOUTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T0_SOUTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B17(Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B17(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_WEST_SB_IN_B17_ready(Tile_X02_Y04_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_IN_B17_valid(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_IN_B1_ready(Tile_X02_Y04_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_IN_B1_valid(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B17(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_WEST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B17(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_EAST_SB_IN_B17_ready(Tile_X02_Y04_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_IN_B17_valid(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_IN_B1_ready(Tile_X02_Y04_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_IN_B1_valid(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B17(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_EAST_SB_OUT_B17_ready(Tile_X03_Y04_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_OUT_B1_ready(Tile_X03_Y04_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B17(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B17(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T1_SOUTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T1_SOUTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B17(Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B17(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_WEST_SB_IN_B17_ready(Tile_X02_Y04_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_IN_B17_valid(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_IN_B1_ready(Tile_X02_Y04_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_IN_B1_valid(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B17(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_WEST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B17(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_EAST_SB_IN_B17_ready(Tile_X02_Y04_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_IN_B17_valid(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_IN_B1_ready(Tile_X02_Y04_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_IN_B1_valid(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B17(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_EAST_SB_OUT_B17_ready(Tile_X03_Y04_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_OUT_B1_ready(Tile_X03_Y04_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B17(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B17(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T2_SOUTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T2_SOUTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B17(Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B17(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_WEST_SB_IN_B17_ready(Tile_X02_Y04_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_IN_B17_valid(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_IN_B1_ready(Tile_X02_Y04_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_IN_B1_valid(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B17(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_WEST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B17(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_EAST_SB_IN_B17_ready(Tile_X02_Y04_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_IN_B17_valid(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_IN_B1_ready(Tile_X02_Y04_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_IN_B1_valid(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B17(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_EAST_SB_OUT_B17_ready(Tile_X03_Y04_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_OUT_B1_ready(Tile_X03_Y04_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B17(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B17(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T3_SOUTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T3_SOUTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B17(Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B17(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_WEST_SB_IN_B17_ready(Tile_X02_Y04_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_IN_B17_valid(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_IN_B1_ready(Tile_X02_Y04_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_IN_B1_valid(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B17(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_WEST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B17(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_EAST_SB_IN_B17_ready(Tile_X02_Y04_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_IN_B17_valid(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_IN_B1_ready(Tile_X02_Y04_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_IN_B1_valid(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B17(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_EAST_SB_OUT_B17_ready(Tile_X03_Y04_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_OUT_B1_ready(Tile_X03_Y04_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B17(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_IN_B17_valid(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_IN_B1_valid(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B17(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_OUT_B17_ready(Tile_X02_Y03_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_OUT_B1_ready(Tile_X02_Y03_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T4_SOUTH_SB_IN_B17_ready(Tile_X02_Y04_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T4_SOUTH_SB_IN_B1_ready(Tile_X02_Y04_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B17(Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B17(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_WEST_SB_IN_B17_ready(Tile_X02_Y04_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_IN_B17_valid(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_IN_B1_ready(Tile_X02_Y04_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_IN_B1_valid(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B17(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_WEST_SB_OUT_B17_ready(Tile_X01_Y04_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_OUT_B17_valid(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_OUT_B1_ready(Tile_X01_Y04_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_OUT_B1_valid(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B1_valid),
    .clk(Tile_X02_Y03_clk_out),
    .clk_out(Tile_X02_Y04_clk_out),
    .clk_pass_through(Tile_X02_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y04_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y03_config_out_config_addr),
    .config_config_data(Tile_X02_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y04_config_out_config_data),
    .config_out_read(Tile_X02_Y04_config_out_read),
    .config_out_write(Tile_X02_Y04_config_out_write),
    .config_read(Tile_X02_Y03_config_out_read),
    .config_write(Tile_X02_Y03_config_out_write),
    .flush(Tile_X02_Y03_flush_out),
    .flush_out(Tile_X02_Y04_flush_out),
    .hi(Tile_X02_Y04_hi),
    .lo(Tile_X02_Y04_lo),
    .read_config_data(Tile_X02_Y04_read_config_data),
    .read_config_data_in(Tile_X02_Y03_read_config_data),
    .reset(Tile_X02_Y03_reset_out),
    .reset_out(Tile_X02_Y04_reset_out),
    .stall(Tile_X02_Y03_stall_out),
    .stall_out(Tile_X02_Y04_stall_out),
    .tile_id(Tile_X02_Y04_tile_id)
);
wire [31:0] Tile_X03_Y00_config_config_addr;
assign Tile_X03_Y00_config_config_addr = {PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[31],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[30],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[29],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[28],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[27],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[26],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[25],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[24],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[23],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[22],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[21],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[20],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[19],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[18],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[17],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[16],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[15],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[14],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[13],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[12],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[11],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[10],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[9],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[8],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[7],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[6],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[5],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[4],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[3],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[2],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[1],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[0]};
wire [31:0] Tile_X03_Y00_config_config_data;
assign Tile_X03_Y00_config_config_data = {PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[63],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[62],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[61],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[60],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[59],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[58],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[57],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[56],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[55],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[54],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[53],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[52],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[51],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[50],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[49],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[48],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[47],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[46],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[45],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[44],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[43],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[42],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[41],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[40],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[39],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[38],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[37],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[36],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[35],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[34],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[33],PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[32]};
wire [4:0] Tile_X03_Y00_io2f_17_ready;
assign Tile_X03_Y00_io2f_17_ready = {Tile_X03_Y01_SB_T4_NORTH_SB_IN_B17_ready,Tile_X03_Y01_SB_T3_NORTH_SB_IN_B17_ready,Tile_X03_Y01_SB_T2_NORTH_SB_IN_B17_ready,Tile_X03_Y01_SB_T1_NORTH_SB_IN_B17_ready,Tile_X03_Y01_SB_T0_NORTH_SB_IN_B17_ready};
wire [4:0] Tile_X03_Y00_io2f_1_ready;
assign Tile_X03_Y00_io2f_1_ready = {Tile_X03_Y01_SB_T4_NORTH_SB_IN_B1_ready,Tile_X03_Y01_SB_T3_NORTH_SB_IN_B1_ready,Tile_X03_Y01_SB_T2_NORTH_SB_IN_B1_ready,Tile_X03_Y01_SB_T1_NORTH_SB_IN_B1_ready,Tile_X03_Y01_SB_T0_NORTH_SB_IN_B1_ready};
wire [15:0] Tile_X03_Y00_tile_id;
assign Tile_X03_Y00_tile_id = {Tile_X03_Y00_lo[7],Tile_X03_Y00_lo[7],Tile_X03_Y00_lo[6],Tile_X03_Y00_lo[6],Tile_X03_Y00_lo[5],Tile_X03_Y00_lo[5],Tile_X03_Y00_hi[5],Tile_X03_Y00_hi[4],Tile_X03_Y00_lo[3],Tile_X03_Y00_lo[3],Tile_X03_Y00_lo[2],Tile_X03_Y00_lo[2],Tile_X03_Y00_lo[1],Tile_X03_Y00_lo[1],Tile_X03_Y00_lo[0],Tile_X03_Y00_lo[0]};
Tile_IOCoreReadyValid Tile_X03_Y00 (
    .clk(clk),
    .clk_out(Tile_X03_Y00_clk_out),
    .config_config_addr(Tile_X03_Y00_config_config_addr),
    .config_config_data(Tile_X03_Y00_config_config_data),
    .config_out_config_addr(Tile_X03_Y00_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y00_config_out_config_data),
    .config_out_read(Tile_X03_Y00_config_out_read),
    .config_out_write(Tile_X03_Y00_config_out_write),
    .config_read(PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[64]),
    .config_write(PipelineRegister_inst7$Register_inst0$reg_P66_inst0_out[65]),
    .f2io_1(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1),
    .f2io_17(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B17),
    .f2io_17_ready(Tile_X03_Y00_f2io_17_ready),
    .f2io_17_valid(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B17_valid),
    .f2io_1_ready(Tile_X03_Y00_f2io_1_ready),
    .f2io_1_valid(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1_valid),
    .flush(PipelineRegister_inst3$Register_inst0$reg_P1_inst0_out),
    .flush_out(Tile_X03_Y00_flush_out),
    .glb2io_1(glb2io_1_X03_Y00),
    .glb2io_17(glb2io_17_X03_Y00),
    .glb2io_17_ready(Tile_X03_Y00_glb2io_17_ready),
    .glb2io_17_valid(glb2io_17_X03_Y00_valid),
    .glb2io_1_ready(Tile_X03_Y00_glb2io_1_ready),
    .glb2io_1_valid(glb2io_1_X03_Y00_valid),
    .hi(Tile_X03_Y00_hi),
    .io2f_1(Tile_X03_Y00_io2f_1),
    .io2f_17(Tile_X03_Y00_io2f_17),
    .io2f_17_ready(Tile_X03_Y00_io2f_17_ready),
    .io2f_17_valid(Tile_X03_Y00_io2f_17_valid),
    .io2f_1_ready(Tile_X03_Y00_io2f_1_ready),
    .io2f_1_valid(Tile_X03_Y00_io2f_1_valid),
    .io2glb_1(Tile_X03_Y00_io2glb_1),
    .io2glb_17(Tile_X03_Y00_io2glb_17),
    .io2glb_17_ready(io2glb_17_X03_Y00_ready),
    .io2glb_17_valid(Tile_X03_Y00_io2glb_17_valid),
    .io2glb_1_ready(io2glb_1_X03_Y00_ready),
    .io2glb_1_valid(Tile_X03_Y00_io2glb_1_valid),
    .lo(Tile_X03_Y00_lo),
    .read_config_data(Tile_X03_Y00_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X03_Y00_reset_out),
    .stall(self_stall_out[3:3]),
    .stall_out(Tile_X03_Y00_stall_out),
    .tile_id(Tile_X03_Y00_tile_id)
);
wire [15:0] Tile_X03_Y01_tile_id;
assign Tile_X03_Y01_tile_id = {Tile_X03_Y01_lo[7],Tile_X03_Y01_lo[7],Tile_X03_Y01_lo[6],Tile_X03_Y01_lo[6],Tile_X03_Y01_lo[5],Tile_X03_Y01_lo[5],Tile_X03_Y01_hi[5],Tile_X03_Y01_hi[4],Tile_X03_Y01_lo[3],Tile_X03_Y01_lo[3],Tile_X03_Y01_lo[2],Tile_X03_Y01_lo[2],Tile_X03_Y01_lo[1],Tile_X03_Y01_lo[1],Tile_X03_Y01_lo[0],Tile_X03_Y01_hi[0]};
Tile_MemCore Tile_X03_Y01 (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B17(const_0_17_out),
    .SB_T0_EAST_SB_IN_B17_ready(Tile_X03_Y01_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T0_EAST_SB_IN_B1_ready(Tile_X03_Y01_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B17(Tile_X03_Y01_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T0_EAST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T0_EAST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B17(Tile_X03_Y00_io2f_17),
    .SB_T0_NORTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_IN_B17_valid(Tile_X03_Y00_io2f_17_valid),
    .SB_T0_NORTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_IN_B1_valid(Tile_X03_Y00_io2f_1_valid),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B17(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_OUT_B17_ready(Tile_X03_Y00_f2io_17_ready),
    .SB_T0_NORTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_OUT_B1_ready(Tile_X03_Y00_f2io_1_ready),
    .SB_T0_NORTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B17(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B17(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B17(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_WEST_SB_IN_B17_ready(Tile_X03_Y01_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_IN_B17_valid(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_IN_B1_ready(Tile_X03_Y01_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_IN_B1_valid(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B17(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_WEST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B17(const_0_17_out),
    .SB_T1_EAST_SB_IN_B17_ready(Tile_X03_Y01_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T1_EAST_SB_IN_B1_ready(Tile_X03_Y01_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B17(Tile_X03_Y01_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T1_EAST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T1_EAST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B17(Tile_X03_Y00_io2f_17),
    .SB_T1_NORTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_IN_B17_valid(Tile_X03_Y00_io2f_17_valid),
    .SB_T1_NORTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_IN_B1_valid(Tile_X03_Y00_io2f_1_valid),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B17(Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T1_NORTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T1_NORTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B17(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B17(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B17(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_WEST_SB_IN_B17_ready(Tile_X03_Y01_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_IN_B17_valid(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_IN_B1_ready(Tile_X03_Y01_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_IN_B1_valid(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B17(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_WEST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B17(const_0_17_out),
    .SB_T2_EAST_SB_IN_B17_ready(Tile_X03_Y01_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T2_EAST_SB_IN_B1_ready(Tile_X03_Y01_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B17(Tile_X03_Y01_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T2_EAST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T2_EAST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B17(Tile_X03_Y00_io2f_17),
    .SB_T2_NORTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_IN_B17_valid(Tile_X03_Y00_io2f_17_valid),
    .SB_T2_NORTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_IN_B1_valid(Tile_X03_Y00_io2f_1_valid),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B17(Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T2_NORTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T2_NORTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B17(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B17(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B17(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_WEST_SB_IN_B17_ready(Tile_X03_Y01_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_IN_B17_valid(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_IN_B1_ready(Tile_X03_Y01_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_IN_B1_valid(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B17(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_WEST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B17(const_0_17_out),
    .SB_T3_EAST_SB_IN_B17_ready(Tile_X03_Y01_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T3_EAST_SB_IN_B1_ready(Tile_X03_Y01_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B17(Tile_X03_Y01_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T3_EAST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T3_EAST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B17(Tile_X03_Y00_io2f_17),
    .SB_T3_NORTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_IN_B17_valid(Tile_X03_Y00_io2f_17_valid),
    .SB_T3_NORTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_IN_B1_valid(Tile_X03_Y00_io2f_1_valid),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B17(Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T3_NORTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T3_NORTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B17(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B17(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B17(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_WEST_SB_IN_B17_ready(Tile_X03_Y01_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_IN_B17_valid(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_IN_B1_ready(Tile_X03_Y01_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_IN_B1_valid(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B17(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_WEST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B17(const_0_17_out),
    .SB_T4_EAST_SB_IN_B17_ready(Tile_X03_Y01_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T4_EAST_SB_IN_B1_ready(Tile_X03_Y01_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B17(Tile_X03_Y01_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T4_EAST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T4_EAST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B17(Tile_X03_Y00_io2f_17),
    .SB_T4_NORTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_IN_B17_valid(Tile_X03_Y00_io2f_17_valid),
    .SB_T4_NORTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_IN_B1_valid(Tile_X03_Y00_io2f_1_valid),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B17(Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T4_NORTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T4_NORTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B17(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_IN_B17_ready(Tile_X03_Y01_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_IN_B1_ready(Tile_X03_Y01_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B17(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B17(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_WEST_SB_IN_B17_ready(Tile_X03_Y01_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_IN_B17_valid(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_IN_B1_ready(Tile_X03_Y01_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_IN_B1_valid(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B17(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_WEST_SB_OUT_B17_ready(Tile_X02_Y01_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_OUT_B17_valid(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_OUT_B1_ready(Tile_X02_Y01_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_OUT_B1_valid(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B1_valid),
    .clk(Tile_X02_Y01_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y01_clk_out),
    .config_config_addr(Tile_X03_Y00_config_out_config_addr),
    .config_config_data(Tile_X03_Y00_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y01_config_out_config_data),
    .config_out_read(Tile_X03_Y01_config_out_read),
    .config_out_write(Tile_X03_Y01_config_out_write),
    .config_read(Tile_X03_Y00_config_out_read),
    .config_write(Tile_X03_Y00_config_out_write),
    .flush(Tile_X03_Y00_flush_out),
    .flush_out(Tile_X03_Y01_flush_out),
    .hi(Tile_X03_Y01_hi),
    .lo(Tile_X03_Y01_lo),
    .read_config_data(Tile_X03_Y01_read_config_data),
    .read_config_data_in(Tile_X03_Y00_read_config_data),
    .reset(Tile_X03_Y00_reset_out),
    .reset_out(Tile_X03_Y01_reset_out),
    .stall(Tile_X03_Y00_stall_out),
    .stall_out(Tile_X03_Y01_stall_out),
    .tile_id(Tile_X03_Y01_tile_id)
);
wire [15:0] Tile_X03_Y02_tile_id;
assign Tile_X03_Y02_tile_id = {Tile_X03_Y02_lo[7],Tile_X03_Y02_lo[7],Tile_X03_Y02_lo[6],Tile_X03_Y02_lo[6],Tile_X03_Y02_lo[5],Tile_X03_Y02_lo[5],Tile_X03_Y02_hi[5],Tile_X03_Y02_hi[4],Tile_X03_Y02_lo[3],Tile_X03_Y02_lo[3],Tile_X03_Y02_lo[2],Tile_X03_Y02_lo[2],Tile_X03_Y02_lo[1],Tile_X03_Y02_lo[1],Tile_X03_Y02_hi[1],Tile_X03_Y02_lo[0]};
Tile_MemCore Tile_X03_Y02 (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B17(const_0_17_out),
    .SB_T0_EAST_SB_IN_B17_ready(Tile_X03_Y02_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T0_EAST_SB_IN_B1_ready(Tile_X03_Y02_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B17(Tile_X03_Y02_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T0_EAST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T0_EAST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B17(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_IN_B17_valid(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_IN_B1_valid(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B17(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_OUT_B17_ready(Tile_X03_Y01_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_OUT_B1_ready(Tile_X03_Y01_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B17(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B17(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B17(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_WEST_SB_IN_B17_ready(Tile_X03_Y02_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_IN_B17_valid(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_IN_B1_ready(Tile_X03_Y02_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_IN_B1_valid(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B17(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_WEST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B17(const_0_17_out),
    .SB_T1_EAST_SB_IN_B17_ready(Tile_X03_Y02_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T1_EAST_SB_IN_B1_ready(Tile_X03_Y02_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B17(Tile_X03_Y02_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T1_EAST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T1_EAST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B17(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_IN_B17_valid(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_IN_B1_valid(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B17(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_OUT_B17_ready(Tile_X03_Y01_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_OUT_B1_ready(Tile_X03_Y01_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B17(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B17(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B17(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_WEST_SB_IN_B17_ready(Tile_X03_Y02_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_IN_B17_valid(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_IN_B1_ready(Tile_X03_Y02_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_IN_B1_valid(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B17(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_WEST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B17(const_0_17_out),
    .SB_T2_EAST_SB_IN_B17_ready(Tile_X03_Y02_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T2_EAST_SB_IN_B1_ready(Tile_X03_Y02_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B17(Tile_X03_Y02_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T2_EAST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T2_EAST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B17(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_IN_B17_valid(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_IN_B1_valid(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B17(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_OUT_B17_ready(Tile_X03_Y01_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_OUT_B1_ready(Tile_X03_Y01_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B17(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B17(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B17(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_WEST_SB_IN_B17_ready(Tile_X03_Y02_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_IN_B17_valid(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_IN_B1_ready(Tile_X03_Y02_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_IN_B1_valid(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B17(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_WEST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B17(const_0_17_out),
    .SB_T3_EAST_SB_IN_B17_ready(Tile_X03_Y02_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T3_EAST_SB_IN_B1_ready(Tile_X03_Y02_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B17(Tile_X03_Y02_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T3_EAST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T3_EAST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B17(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_IN_B17_valid(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_IN_B1_valid(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B17(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_OUT_B17_ready(Tile_X03_Y01_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_OUT_B1_ready(Tile_X03_Y01_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B17(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B17(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B17(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_WEST_SB_IN_B17_ready(Tile_X03_Y02_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_IN_B17_valid(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_IN_B1_ready(Tile_X03_Y02_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_IN_B1_valid(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B17(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_WEST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B17(const_0_17_out),
    .SB_T4_EAST_SB_IN_B17_ready(Tile_X03_Y02_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T4_EAST_SB_IN_B1_ready(Tile_X03_Y02_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B17(Tile_X03_Y02_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T4_EAST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T4_EAST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B17(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_IN_B17_valid(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_IN_B1_valid(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B17(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_OUT_B17_ready(Tile_X03_Y01_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_OUT_B1_ready(Tile_X03_Y01_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B17(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_IN_B17_ready(Tile_X03_Y02_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_IN_B1_ready(Tile_X03_Y02_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B17(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B17(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_WEST_SB_IN_B17_ready(Tile_X03_Y02_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_IN_B17_valid(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_IN_B1_ready(Tile_X03_Y02_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_IN_B1_valid(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B17(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_WEST_SB_OUT_B17_ready(Tile_X02_Y02_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_OUT_B17_valid(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_OUT_B1_ready(Tile_X02_Y02_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_OUT_B1_valid(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B1_valid),
    .clk(Tile_X02_Y02_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y02_clk_out),
    .config_config_addr(Tile_X03_Y01_config_out_config_addr),
    .config_config_data(Tile_X03_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y02_config_out_config_data),
    .config_out_read(Tile_X03_Y02_config_out_read),
    .config_out_write(Tile_X03_Y02_config_out_write),
    .config_read(Tile_X03_Y01_config_out_read),
    .config_write(Tile_X03_Y01_config_out_write),
    .flush(Tile_X03_Y01_flush_out),
    .flush_out(Tile_X03_Y02_flush_out),
    .hi(Tile_X03_Y02_hi),
    .lo(Tile_X03_Y02_lo),
    .read_config_data(Tile_X03_Y02_read_config_data),
    .read_config_data_in(Tile_X03_Y01_read_config_data),
    .reset(Tile_X03_Y01_reset_out),
    .reset_out(Tile_X03_Y02_reset_out),
    .stall(Tile_X03_Y01_stall_out),
    .stall_out(Tile_X03_Y02_stall_out),
    .tile_id(Tile_X03_Y02_tile_id)
);
wire [15:0] Tile_X03_Y03_tile_id;
assign Tile_X03_Y03_tile_id = {Tile_X03_Y03_lo[7],Tile_X03_Y03_lo[7],Tile_X03_Y03_lo[6],Tile_X03_Y03_lo[6],Tile_X03_Y03_lo[5],Tile_X03_Y03_lo[5],Tile_X03_Y03_hi[5],Tile_X03_Y03_hi[4],Tile_X03_Y03_lo[3],Tile_X03_Y03_lo[3],Tile_X03_Y03_lo[2],Tile_X03_Y03_lo[2],Tile_X03_Y03_lo[1],Tile_X03_Y03_lo[1],Tile_X03_Y03_hi[1],Tile_X03_Y03_hi[0]};
Tile_MemCore Tile_X03_Y03 (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B17(const_0_17_out),
    .SB_T0_EAST_SB_IN_B17_ready(Tile_X03_Y03_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T0_EAST_SB_IN_B1_ready(Tile_X03_Y03_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B17(Tile_X03_Y03_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T0_EAST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T0_EAST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B17(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B17(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B17(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_IN_B17_valid(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_IN_B1_valid(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B17(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_OUT_B17_ready(Tile_X03_Y04_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_OUT_B1_ready(Tile_X03_Y04_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B17(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_WEST_SB_IN_B17_ready(Tile_X03_Y03_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_IN_B17_valid(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_IN_B1_ready(Tile_X03_Y03_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_IN_B1_valid(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B17(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_WEST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B17(const_0_17_out),
    .SB_T1_EAST_SB_IN_B17_ready(Tile_X03_Y03_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T1_EAST_SB_IN_B1_ready(Tile_X03_Y03_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B17(Tile_X03_Y03_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T1_EAST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T1_EAST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B17(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B17(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B17(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_IN_B17_valid(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_IN_B1_valid(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B17(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_OUT_B17_ready(Tile_X03_Y04_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_OUT_B1_ready(Tile_X03_Y04_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B17(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_WEST_SB_IN_B17_ready(Tile_X03_Y03_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_IN_B17_valid(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_IN_B1_ready(Tile_X03_Y03_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_IN_B1_valid(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B17(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_WEST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B17(const_0_17_out),
    .SB_T2_EAST_SB_IN_B17_ready(Tile_X03_Y03_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T2_EAST_SB_IN_B1_ready(Tile_X03_Y03_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B17(Tile_X03_Y03_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T2_EAST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T2_EAST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B17(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B17(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B17(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_IN_B17_valid(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_IN_B1_valid(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B17(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_OUT_B17_ready(Tile_X03_Y04_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_OUT_B1_ready(Tile_X03_Y04_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B17(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_WEST_SB_IN_B17_ready(Tile_X03_Y03_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_IN_B17_valid(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_IN_B1_ready(Tile_X03_Y03_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_IN_B1_valid(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B17(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_WEST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B17(const_0_17_out),
    .SB_T3_EAST_SB_IN_B17_ready(Tile_X03_Y03_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T3_EAST_SB_IN_B1_ready(Tile_X03_Y03_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B17(Tile_X03_Y03_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T3_EAST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T3_EAST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B17(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B17(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B17(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_IN_B17_valid(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_IN_B1_valid(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B17(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_OUT_B17_ready(Tile_X03_Y04_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_OUT_B1_ready(Tile_X03_Y04_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B17(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_WEST_SB_IN_B17_ready(Tile_X03_Y03_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_IN_B17_valid(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_IN_B1_ready(Tile_X03_Y03_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_IN_B1_valid(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B17(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_WEST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B17(const_0_17_out),
    .SB_T4_EAST_SB_IN_B17_ready(Tile_X03_Y03_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T4_EAST_SB_IN_B1_ready(Tile_X03_Y03_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B17(Tile_X03_Y03_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T4_EAST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T4_EAST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B17(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_IN_B17_valid(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_IN_B1_valid(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B17(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_OUT_B17_ready(Tile_X03_Y02_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_OUT_B1_ready(Tile_X03_Y02_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B17(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_IN_B17_ready(Tile_X03_Y03_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_IN_B17_valid(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_IN_B1_ready(Tile_X03_Y03_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_IN_B1_valid(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B17(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_OUT_B17_ready(Tile_X03_Y04_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_OUT_B1_ready(Tile_X03_Y04_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B17(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_WEST_SB_IN_B17_ready(Tile_X03_Y03_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_IN_B17_valid(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_IN_B1_ready(Tile_X03_Y03_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_IN_B1_valid(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B17(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_WEST_SB_OUT_B17_ready(Tile_X02_Y03_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_OUT_B17_valid(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_OUT_B1_ready(Tile_X02_Y03_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_OUT_B1_valid(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B1_valid),
    .clk(Tile_X02_Y03_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y03_clk_out),
    .config_config_addr(Tile_X03_Y02_config_out_config_addr),
    .config_config_data(Tile_X03_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y03_config_out_config_data),
    .config_out_read(Tile_X03_Y03_config_out_read),
    .config_out_write(Tile_X03_Y03_config_out_write),
    .config_read(Tile_X03_Y02_config_out_read),
    .config_write(Tile_X03_Y02_config_out_write),
    .flush(Tile_X03_Y02_flush_out),
    .flush_out(Tile_X03_Y03_flush_out),
    .hi(Tile_X03_Y03_hi),
    .lo(Tile_X03_Y03_lo),
    .read_config_data(Tile_X03_Y03_read_config_data),
    .read_config_data_in(Tile_X03_Y02_read_config_data),
    .reset(Tile_X03_Y02_reset_out),
    .reset_out(Tile_X03_Y03_reset_out),
    .stall(Tile_X03_Y02_stall_out),
    .stall_out(Tile_X03_Y03_stall_out),
    .tile_id(Tile_X03_Y03_tile_id)
);
wire [15:0] Tile_X03_Y04_tile_id;
assign Tile_X03_Y04_tile_id = {Tile_X03_Y04_lo[7],Tile_X03_Y04_lo[7],Tile_X03_Y04_lo[6],Tile_X03_Y04_lo[6],Tile_X03_Y04_lo[5],Tile_X03_Y04_lo[5],Tile_X03_Y04_hi[5],Tile_X03_Y04_hi[4],Tile_X03_Y04_lo[3],Tile_X03_Y04_lo[3],Tile_X03_Y04_lo[2],Tile_X03_Y04_lo[2],Tile_X03_Y04_lo[1],Tile_X03_Y04_hi[1],Tile_X03_Y04_lo[0],Tile_X03_Y04_lo[0]};
Tile_MemCore Tile_X03_Y04 (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B17(const_0_17_out),
    .SB_T0_EAST_SB_IN_B17_ready(Tile_X03_Y04_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T0_EAST_SB_IN_B1_ready(Tile_X03_Y04_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B17(Tile_X03_Y04_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T0_EAST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T0_EAST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B17(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T0_NORTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T0_NORTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B17(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B17),
    .SB_T0_NORTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_NORTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B17_valid),
    .SB_T0_NORTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_NORTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1_valid),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T0_SOUTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T0_SOUTH_SB_IN_B17_ready),
    .SB_T0_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T0_SOUTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T0_SOUTH_SB_IN_B1_ready),
    .SB_T0_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B17(Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B17),
    .SB_T0_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T0_SOUTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B17_valid),
    .SB_T0_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T0_SOUTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B17(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B17),
    .SB_T0_WEST_SB_IN_B17_ready(Tile_X03_Y04_SB_T0_WEST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_IN_B17_valid(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_IN_B1_ready(Tile_X03_Y04_SB_T0_WEST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_IN_B1_valid(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1_valid),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B17(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B17),
    .SB_T0_WEST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T0_EAST_SB_IN_B17_ready),
    .SB_T0_WEST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B17_valid),
    .SB_T0_WEST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T0_EAST_SB_IN_B1_ready),
    .SB_T0_WEST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1_valid),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B17(const_0_17_out),
    .SB_T1_EAST_SB_IN_B17_ready(Tile_X03_Y04_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T1_EAST_SB_IN_B1_ready(Tile_X03_Y04_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B17(Tile_X03_Y04_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T1_EAST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T1_EAST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B17(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T1_NORTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T1_NORTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B17(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B17),
    .SB_T1_NORTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_NORTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B17_valid),
    .SB_T1_NORTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_NORTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1_valid),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T1_SOUTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T1_SOUTH_SB_IN_B17_ready),
    .SB_T1_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T1_SOUTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T1_SOUTH_SB_IN_B1_ready),
    .SB_T1_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B17(Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B17),
    .SB_T1_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T1_SOUTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B17_valid),
    .SB_T1_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T1_SOUTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B17(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B17),
    .SB_T1_WEST_SB_IN_B17_ready(Tile_X03_Y04_SB_T1_WEST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_IN_B17_valid(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_IN_B1_ready(Tile_X03_Y04_SB_T1_WEST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_IN_B1_valid(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1_valid),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B17(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B17),
    .SB_T1_WEST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T1_EAST_SB_IN_B17_ready),
    .SB_T1_WEST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B17_valid),
    .SB_T1_WEST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T1_EAST_SB_IN_B1_ready),
    .SB_T1_WEST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1_valid),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B17(const_0_17_out),
    .SB_T2_EAST_SB_IN_B17_ready(Tile_X03_Y04_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T2_EAST_SB_IN_B1_ready(Tile_X03_Y04_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B17(Tile_X03_Y04_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T2_EAST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T2_EAST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B17(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T2_NORTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T2_NORTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B17(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B17),
    .SB_T2_NORTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_NORTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B17_valid),
    .SB_T2_NORTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_NORTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1_valid),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T2_SOUTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T2_SOUTH_SB_IN_B17_ready),
    .SB_T2_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T2_SOUTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T2_SOUTH_SB_IN_B1_ready),
    .SB_T2_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B17(Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B17),
    .SB_T2_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T2_SOUTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B17_valid),
    .SB_T2_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T2_SOUTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B17(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B17),
    .SB_T2_WEST_SB_IN_B17_ready(Tile_X03_Y04_SB_T2_WEST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_IN_B17_valid(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_IN_B1_ready(Tile_X03_Y04_SB_T2_WEST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_IN_B1_valid(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1_valid),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B17(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B17),
    .SB_T2_WEST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T2_EAST_SB_IN_B17_ready),
    .SB_T2_WEST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B17_valid),
    .SB_T2_WEST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T2_EAST_SB_IN_B1_ready),
    .SB_T2_WEST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1_valid),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B17(const_0_17_out),
    .SB_T3_EAST_SB_IN_B17_ready(Tile_X03_Y04_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T3_EAST_SB_IN_B1_ready(Tile_X03_Y04_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B17(Tile_X03_Y04_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T3_EAST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T3_EAST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B17(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T3_NORTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T3_NORTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B17(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B17),
    .SB_T3_NORTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_NORTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B17_valid),
    .SB_T3_NORTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_NORTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B1_valid),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T3_SOUTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T3_SOUTH_SB_IN_B17_ready),
    .SB_T3_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T3_SOUTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T3_SOUTH_SB_IN_B1_ready),
    .SB_T3_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B17(Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B17),
    .SB_T3_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T3_SOUTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B17_valid),
    .SB_T3_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T3_SOUTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B17(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B17),
    .SB_T3_WEST_SB_IN_B17_ready(Tile_X03_Y04_SB_T3_WEST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_IN_B17_valid(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_IN_B1_ready(Tile_X03_Y04_SB_T3_WEST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_IN_B1_valid(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B1_valid),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B17(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B17),
    .SB_T3_WEST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T3_EAST_SB_IN_B17_ready),
    .SB_T3_WEST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B17_valid),
    .SB_T3_WEST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T3_EAST_SB_IN_B1_ready),
    .SB_T3_WEST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B1_valid),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B17(const_0_17_out),
    .SB_T4_EAST_SB_IN_B17_ready(Tile_X03_Y04_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_EAST_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T4_EAST_SB_IN_B1_ready(Tile_X03_Y04_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_EAST_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B17(Tile_X03_Y04_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_EAST_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T4_EAST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_EAST_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T4_EAST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B17(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T4_NORTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_IN_B17_valid(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T4_NORTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_IN_B1_valid(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B17(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B17),
    .SB_T4_NORTH_SB_OUT_B17_ready(Tile_X03_Y03_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_NORTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B17_valid),
    .SB_T4_NORTH_SB_OUT_B1_ready(Tile_X03_Y03_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_NORTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B1_valid),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B17(const_0_17_out),
    .SB_T4_SOUTH_SB_IN_B17_ready(Tile_X03_Y04_SB_T4_SOUTH_SB_IN_B17_ready),
    .SB_T4_SOUTH_SB_IN_B17_valid(bit_const_0_None_out),
    .SB_T4_SOUTH_SB_IN_B1_ready(Tile_X03_Y04_SB_T4_SOUTH_SB_IN_B1_ready),
    .SB_T4_SOUTH_SB_IN_B1_valid(bit_const_0_None_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B17(Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B17),
    .SB_T4_SOUTH_SB_OUT_B17_ready(bit_const_0_None_out),
    .SB_T4_SOUTH_SB_OUT_B17_valid(Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B17_valid),
    .SB_T4_SOUTH_SB_OUT_B1_ready(bit_const_0_None_out),
    .SB_T4_SOUTH_SB_OUT_B1_valid(Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B17(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B17),
    .SB_T4_WEST_SB_IN_B17_ready(Tile_X03_Y04_SB_T4_WEST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_IN_B17_valid(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_IN_B1_ready(Tile_X03_Y04_SB_T4_WEST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_IN_B1_valid(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B1_valid),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B17(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B17),
    .SB_T4_WEST_SB_OUT_B17_ready(Tile_X02_Y04_SB_T4_EAST_SB_IN_B17_ready),
    .SB_T4_WEST_SB_OUT_B17_valid(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B17_valid),
    .SB_T4_WEST_SB_OUT_B1_ready(Tile_X02_Y04_SB_T4_EAST_SB_IN_B1_ready),
    .SB_T4_WEST_SB_OUT_B1_valid(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B1_valid),
    .clk(Tile_X02_Y04_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y04_clk_out),
    .config_config_addr(Tile_X03_Y03_config_out_config_addr),
    .config_config_data(Tile_X03_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y04_config_out_config_data),
    .config_out_read(Tile_X03_Y04_config_out_read),
    .config_out_write(Tile_X03_Y04_config_out_write),
    .config_read(Tile_X03_Y03_config_out_read),
    .config_write(Tile_X03_Y03_config_out_write),
    .flush(Tile_X03_Y03_flush_out),
    .flush_out(Tile_X03_Y04_flush_out),
    .hi(Tile_X03_Y04_hi),
    .lo(Tile_X03_Y04_lo),
    .read_config_data(Tile_X03_Y04_read_config_data),
    .read_config_data_in(Tile_X03_Y03_read_config_data),
    .reset(Tile_X03_Y03_reset_out),
    .reset_out(Tile_X03_Y04_reset_out),
    .stall(Tile_X03_Y03_stall_out),
    .stall_out(Tile_X03_Y04_stall_out),
    .tile_id(Tile_X03_Y04_tile_id)
);
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
coreir_const #(
    .value(1'h0),
    .width(1)
) const_0_1 (
    .out(const_0_1_out)
);
coreir_const #(
    .value(17'h00000),
    .width(17)
) const_0_17 (
    .out(const_0_17_out)
);
coreir_const #(
    .value(32'h00000000),
    .width(32)
) const_0_32 (
    .out(const_0_32_out)
);
coreir_wrap coreir_wrapInClock_inst0 (
    .in(clk),
    .out(coreir_wrapInClock_inst0_out)
);
coreir_wrap coreir_wrapInClock_inst1 (
    .in(clk),
    .out(coreir_wrapInClock_inst1_out)
);
coreir_wrap coreir_wrapInClock_inst2 (
    .in(clk),
    .out(coreir_wrapInClock_inst2_out)
);
Or4x32 read_config_data_or_final (
    .I0(Tile_X00_Y04_read_config_data),
    .I1(Tile_X01_Y04_read_config_data),
    .I2(Tile_X02_Y04_read_config_data),
    .I3(Tile_X03_Y04_read_config_data),
    .O(read_config_data_or_final_O)
);
mantle_wire__typeBit4 self_stall (
    .in(stall),
    .out(self_stall_out)
);
assign glb2io_17_X00_Y00_ready = Tile_X00_Y00_glb2io_17_ready;
assign glb2io_17_X01_Y00_ready = Tile_X01_Y00_glb2io_17_ready;
assign glb2io_17_X02_Y00_ready = Tile_X02_Y00_glb2io_17_ready;
assign glb2io_17_X03_Y00_ready = Tile_X03_Y00_glb2io_17_ready;
assign glb2io_1_X00_Y00_ready = Tile_X00_Y00_glb2io_1_ready;
assign glb2io_1_X01_Y00_ready = Tile_X01_Y00_glb2io_1_ready;
assign glb2io_1_X02_Y00_ready = Tile_X02_Y00_glb2io_1_ready;
assign glb2io_1_X03_Y00_ready = Tile_X03_Y00_glb2io_1_ready;
assign io2glb_17_X00_Y00 = Tile_X00_Y00_io2glb_17;
assign io2glb_17_X00_Y00_valid = Tile_X00_Y00_io2glb_17_valid;
assign io2glb_17_X01_Y00 = Tile_X01_Y00_io2glb_17;
assign io2glb_17_X01_Y00_valid = Tile_X01_Y00_io2glb_17_valid;
assign io2glb_17_X02_Y00 = Tile_X02_Y00_io2glb_17;
assign io2glb_17_X02_Y00_valid = Tile_X02_Y00_io2glb_17_valid;
assign io2glb_17_X03_Y00 = Tile_X03_Y00_io2glb_17;
assign io2glb_17_X03_Y00_valid = Tile_X03_Y00_io2glb_17_valid;
assign io2glb_1_X00_Y00 = Tile_X00_Y00_io2glb_1;
assign io2glb_1_X00_Y00_valid = Tile_X00_Y00_io2glb_1_valid;
assign io2glb_1_X01_Y00 = Tile_X01_Y00_io2glb_1;
assign io2glb_1_X01_Y00_valid = Tile_X01_Y00_io2glb_1_valid;
assign io2glb_1_X02_Y00 = Tile_X02_Y00_io2glb_1;
assign io2glb_1_X02_Y00_valid = Tile_X02_Y00_io2glb_1_valid;
assign io2glb_1_X03_Y00 = Tile_X03_Y00_io2glb_1;
assign io2glb_1_X03_Y00_valid = Tile_X03_Y00_io2glb_1_valid;
assign read_config_data = read_config_data_or_final_O;
endmodule

module Garnet (
    input [12:0] axi4_slave_araddr,
    output axi4_slave_arready,
    input axi4_slave_arvalid,
    input [12:0] axi4_slave_awaddr,
    output axi4_slave_awready,
    input axi4_slave_awvalid,
    input axi4_slave_bready,
    output [1:0] axi4_slave_bresp,
    output axi4_slave_bvalid,
    output [31:0] axi4_slave_rdata,
    input axi4_slave_rready,
    output [1:0] axi4_slave_rresp,
    output axi4_slave_rvalid,
    input [31:0] axi4_slave_wdata,
    output axi4_slave_wready,
    input axi4_slave_wvalid,
    output cgra_running_clk_out,
    input clk_in,
    output interrupt,
    input jtag_tck,
    input jtag_tdi,
    output jtag_tdo,
    input jtag_tms,
    input jtag_trst_n,
    input [18:0] proc_packet_rd_addr,
    output [63:0] proc_packet_rd_data,
    output proc_packet_rd_data_valid,
    input proc_packet_rd_en,
    input [18:0] proc_packet_wr_addr,
    input [63:0] proc_packet_wr_data,
    input proc_packet_wr_en,
    input [7:0] proc_packet_wr_strb,
    input reset_in
);
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_clk_out;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_reset_out;
wire [3:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_stall;
wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_clk_en_master;
wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_clk_en_bank_master;
wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_pcfg_broadcast_stall;
wire [0:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_flush_crossbar_sel;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_en;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_clk_en;
wire [11:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_addr;
wire [31:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_data;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_en;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_clk_en;
wire [11:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_addr;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_en;
wire [18:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_addr;
wire [31:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_data;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_rd_en;
wire [18:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_rd_addr;
wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_strm_g2f_start_pulse;
wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_strm_f2g_start_pulse;
wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_pc_start_pulse;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_read;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_write;
wire [31:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_addr;
wire [31:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_wr_data;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_awready;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_wready;
wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_bresp;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_bvalid;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_arready;
wire [31:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rdata;
wire [1:0] GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rresp;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rvalid;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_interrupt;
wire GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_tdo;
wire Interconnect_inst0_glb2io_17_X00_Y00_ready;
wire Interconnect_inst0_glb2io_17_X01_Y00_ready;
wire Interconnect_inst0_glb2io_17_X02_Y00_ready;
wire Interconnect_inst0_glb2io_17_X03_Y00_ready;
wire Interconnect_inst0_glb2io_1_X00_Y00_ready;
wire Interconnect_inst0_glb2io_1_X01_Y00_ready;
wire Interconnect_inst0_glb2io_1_X02_Y00_ready;
wire Interconnect_inst0_glb2io_1_X03_Y00_ready;
wire [16:0] Interconnect_inst0_io2glb_17_X00_Y00_unq1;
wire Interconnect_inst0_io2glb_17_X00_Y00_valid;
wire [16:0] Interconnect_inst0_io2glb_17_X01_Y00_unq1;
wire Interconnect_inst0_io2glb_17_X01_Y00_valid;
wire [16:0] Interconnect_inst0_io2glb_17_X02_Y00_unq1;
wire Interconnect_inst0_io2glb_17_X02_Y00_valid;
wire [16:0] Interconnect_inst0_io2glb_17_X03_Y00_unq1;
wire Interconnect_inst0_io2glb_17_X03_Y00_valid;
wire [0:0] Interconnect_inst0_io2glb_1_X00_Y00;
wire Interconnect_inst0_io2glb_1_X00_Y00_valid;
wire [0:0] Interconnect_inst0_io2glb_1_X01_Y00;
wire Interconnect_inst0_io2glb_1_X01_Y00_valid;
wire [0:0] Interconnect_inst0_io2glb_1_X02_Y00;
wire Interconnect_inst0_io2glb_1_X02_Y00_valid;
wire [0:0] Interconnect_inst0_io2glb_1_X03_Y00;
wire Interconnect_inst0_io2glb_1_X03_Y00_valid;
wire [31:0] Interconnect_inst0_read_config_data;
wire [16:0] Interconnect_inst0_glb2io_17_X00_Y00_in;
wire [16:0] Interconnect_inst0_glb2io_17_X01_Y00_in;
wire [16:0] Interconnect_inst0_glb2io_17_X02_Y00_in;
wire [16:0] Interconnect_inst0_glb2io_17_X03_Y00_in;
wire [16:0] Interconnect_inst0_io2glb_17_X00_Y00_out;
wire [16:0] Interconnect_inst0_io2glb_17_X01_Y00_out;
wire [16:0] Interconnect_inst0_io2glb_17_X02_Y00_out;
wire [16:0] Interconnect_inst0_io2glb_17_X03_Y00_out;
wire bit_const_0_None_out;
wire bit_const_1_None_out;
wire [0:0] global_buffer_W_inst0_strm_data_g2f_vld_0_1;
wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_0_1;
wire [15:0] global_buffer_W_inst0_strm_data_g2f_1_1;
wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_0_0;
wire [63:0] global_buffer_W_inst0_proc_rd_data;
wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_0_1;
wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_0_0;
wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_1_1;
wire [15:0] global_buffer_W_inst0_strm_data_g2f_1_0;
wire [1:0] global_buffer_W_inst0_strm_g2f_interrupt_pulse;
wire [0:0] global_buffer_W_inst0_strm_ctrl_g2f_1_0;
wire [0:0] global_buffer_W_inst0_strm_data_g2f_vld_1_0;
wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_0_0;
wire [0:0] global_buffer_W_inst0_strm_data_g2f_vld_0_0;
wire [0:0] global_buffer_W_inst0_strm_data_f2g_rdy_0_1;
wire [0:0] global_buffer_W_inst0_strm_data_g2f_vld_1_1;
wire [0:0] global_buffer_W_inst0_strm_data_flush_g2f;
wire [0:0] global_buffer_W_inst0_strm_ctrl_g2f_0_0;
wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_1_0;
wire [0:0] global_buffer_W_inst0_strm_ctrl_g2f_0_1;
wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_1_1;
wire [0:0] global_buffer_W_inst0_strm_data_f2g_rdy_1_0;
wire [0:0] global_buffer_W_inst0_strm_data_f2g_rdy_0_0;
wire [0:0] global_buffer_W_inst0_strm_ctrl_g2f_1_1;
wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_1_1;
wire [0:0] global_buffer_W_inst0_if_sram_cfg_rd_data_valid;
wire [1:0] global_buffer_W_inst0_pcfg_g2f_interrupt_pulse;
wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_1_1;
wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_0_1;
wire [0:0] global_buffer_W_inst0_if_cfg_rd_data_valid;
wire [3:0] global_buffer_W_inst0_cgra_stall;
wire [31:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_1_0;
wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_0_0;
wire [15:0] global_buffer_W_inst0_strm_data_g2f_0_1;
wire [1:0] global_buffer_W_inst0_strm_f2g_interrupt_pulse;
wire [31:0] global_buffer_W_inst0_if_sram_cfg_rd_data;
wire [0:0] global_buffer_W_inst0_proc_rd_data_valid;
wire [31:0] global_buffer_W_inst0_if_cfg_rd_data;
wire [15:0] global_buffer_W_inst0_strm_data_g2f_0_0;
wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_1_0;
wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_1_0;
wire [0:0] global_buffer_W_inst0_strm_data_f2g_rdy_1_1;
wire [0:0] global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_0_1;
global_controller GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0 (
    .clk_in(clk_in),
    .reset_in(reset_in),
    .clk_out(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_clk_out),
    .reset_out(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_reset_out),
    .cgra_stall(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_stall),
    .glb_clk_en_master(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_clk_en_master),
    .glb_clk_en_bank_master(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_clk_en_bank_master),
    .glb_pcfg_broadcast_stall(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_pcfg_broadcast_stall),
    .glb_flush_crossbar_sel(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_flush_crossbar_sel),
    .glb_cfg_wr_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_en),
    .glb_cfg_wr_clk_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_clk_en),
    .glb_cfg_wr_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_addr),
    .glb_cfg_wr_data(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_data),
    .glb_cfg_rd_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_en),
    .glb_cfg_rd_clk_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_clk_en),
    .glb_cfg_rd_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_addr),
    .glb_cfg_rd_data(global_buffer_W_inst0_if_cfg_rd_data),
    .glb_cfg_rd_data_valid(global_buffer_W_inst0_if_cfg_rd_data_valid[0]),
    .sram_cfg_wr_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_en),
    .sram_cfg_wr_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_addr),
    .sram_cfg_wr_data(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_data),
    .sram_cfg_rd_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_rd_en),
    .sram_cfg_rd_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_rd_addr),
    .sram_cfg_rd_data(global_buffer_W_inst0_if_sram_cfg_rd_data),
    .sram_cfg_rd_data_valid(global_buffer_W_inst0_if_sram_cfg_rd_data_valid[0]),
    .strm_g2f_start_pulse(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_strm_g2f_start_pulse),
    .strm_f2g_start_pulse(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_strm_f2g_start_pulse),
    .pc_start_pulse(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_pc_start_pulse),
    .strm_g2f_interrupt_pulse(global_buffer_W_inst0_strm_g2f_interrupt_pulse),
    .strm_f2g_interrupt_pulse(global_buffer_W_inst0_strm_f2g_interrupt_pulse),
    .pcfg_g2f_interrupt_pulse(global_buffer_W_inst0_pcfg_g2f_interrupt_pulse),
    .cgra_cfg_read(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_read),
    .cgra_cfg_write(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_write),
    .cgra_cfg_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_addr),
    .cgra_cfg_wr_data(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_wr_data),
    .cgra_cfg_rd_data(Interconnect_inst0_read_config_data),
    .axi_awaddr(axi4_slave_awaddr),
    .axi_awvalid(axi4_slave_awvalid),
    .axi_awready(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_awready),
    .axi_wdata(axi4_slave_wdata),
    .axi_wvalid(axi4_slave_wvalid),
    .axi_wready(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_wready),
    .axi_bready(axi4_slave_bready),
    .axi_bresp(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_bresp),
    .axi_bvalid(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_bvalid),
    .axi_araddr(axi4_slave_araddr),
    .axi_arvalid(axi4_slave_arvalid),
    .axi_arready(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_arready),
    .axi_rdata(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rdata),
    .axi_rresp(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rresp),
    .axi_rvalid(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rvalid),
    .axi_rready(axi4_slave_rready),
    .interrupt(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_interrupt),
    .tck(jtag_tck),
    .tdi(jtag_tdi),
    .tms(jtag_tms),
    .trst_n(jtag_trst_n),
    .tdo(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_tdo)
);
Interconnect Interconnect_inst0 (
    .clk(clk_in),
    .config_0_config_addr(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_0_0),
    .config_0_config_data(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_0_0),
    .config_0_read(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_0_0),
    .config_0_write(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_0_0),
    .config_1_config_addr(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_0_1),
    .config_1_config_data(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_0_1),
    .config_1_read(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_0_1),
    .config_1_write(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_0_1),
    .config_2_config_addr(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_1_0),
    .config_2_config_data(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_1_0),
    .config_2_read(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_1_0),
    .config_2_write(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_1_0),
    .config_3_config_addr(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_1_1),
    .config_3_config_data(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_1_1),
    .config_3_read(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_1_1),
    .config_3_write(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_1_1),
    .flush(global_buffer_W_inst0_strm_data_flush_g2f),
    .glb2io_17_X00_Y00(Interconnect_inst0_glb2io_17_X00_Y00_in),
    .glb2io_17_X00_Y00_ready(Interconnect_inst0_glb2io_17_X00_Y00_ready),
    .glb2io_17_X00_Y00_valid(global_buffer_W_inst0_strm_data_g2f_vld_0_0[0]),
    .glb2io_17_X01_Y00(Interconnect_inst0_glb2io_17_X01_Y00_in),
    .glb2io_17_X01_Y00_ready(Interconnect_inst0_glb2io_17_X01_Y00_ready),
    .glb2io_17_X01_Y00_valid(global_buffer_W_inst0_strm_data_g2f_vld_0_1[0]),
    .glb2io_17_X02_Y00(Interconnect_inst0_glb2io_17_X02_Y00_in),
    .glb2io_17_X02_Y00_ready(Interconnect_inst0_glb2io_17_X02_Y00_ready),
    .glb2io_17_X02_Y00_valid(global_buffer_W_inst0_strm_data_g2f_vld_1_0[0]),
    .glb2io_17_X03_Y00(Interconnect_inst0_glb2io_17_X03_Y00_in),
    .glb2io_17_X03_Y00_ready(Interconnect_inst0_glb2io_17_X03_Y00_ready),
    .glb2io_17_X03_Y00_valid(global_buffer_W_inst0_strm_data_g2f_vld_1_1[0]),
    .glb2io_1_X00_Y00(global_buffer_W_inst0_strm_ctrl_g2f_0_0),
    .glb2io_1_X00_Y00_ready(Interconnect_inst0_glb2io_1_X00_Y00_ready),
    .glb2io_1_X00_Y00_valid(bit_const_1_None_out),
    .glb2io_1_X01_Y00(global_buffer_W_inst0_strm_ctrl_g2f_0_1),
    .glb2io_1_X01_Y00_ready(Interconnect_inst0_glb2io_1_X01_Y00_ready),
    .glb2io_1_X01_Y00_valid(bit_const_1_None_out),
    .glb2io_1_X02_Y00(global_buffer_W_inst0_strm_ctrl_g2f_1_0),
    .glb2io_1_X02_Y00_ready(Interconnect_inst0_glb2io_1_X02_Y00_ready),
    .glb2io_1_X02_Y00_valid(bit_const_1_None_out),
    .glb2io_1_X03_Y00(global_buffer_W_inst0_strm_ctrl_g2f_1_1),
    .glb2io_1_X03_Y00_ready(Interconnect_inst0_glb2io_1_X03_Y00_ready),
    .glb2io_1_X03_Y00_valid(bit_const_1_None_out),
    .io2glb_17_X00_Y00(Interconnect_inst0_io2glb_17_X00_Y00_unq1),
    .io2glb_17_X00_Y00_ready(global_buffer_W_inst0_strm_data_f2g_rdy_0_0[0]),
    .io2glb_17_X00_Y00_valid(Interconnect_inst0_io2glb_17_X00_Y00_valid),
    .io2glb_17_X01_Y00(Interconnect_inst0_io2glb_17_X01_Y00_unq1),
    .io2glb_17_X01_Y00_ready(global_buffer_W_inst0_strm_data_f2g_rdy_0_1[0]),
    .io2glb_17_X01_Y00_valid(Interconnect_inst0_io2glb_17_X01_Y00_valid),
    .io2glb_17_X02_Y00(Interconnect_inst0_io2glb_17_X02_Y00_unq1),
    .io2glb_17_X02_Y00_ready(global_buffer_W_inst0_strm_data_f2g_rdy_1_0[0]),
    .io2glb_17_X02_Y00_valid(Interconnect_inst0_io2glb_17_X02_Y00_valid),
    .io2glb_17_X03_Y00(Interconnect_inst0_io2glb_17_X03_Y00_unq1),
    .io2glb_17_X03_Y00_ready(global_buffer_W_inst0_strm_data_f2g_rdy_1_1[0]),
    .io2glb_17_X03_Y00_valid(Interconnect_inst0_io2glb_17_X03_Y00_valid),
    .io2glb_1_X00_Y00(Interconnect_inst0_io2glb_1_X00_Y00),
    .io2glb_1_X00_Y00_ready(bit_const_1_None_out),
    .io2glb_1_X00_Y00_valid(Interconnect_inst0_io2glb_1_X00_Y00_valid),
    .io2glb_1_X01_Y00(Interconnect_inst0_io2glb_1_X01_Y00),
    .io2glb_1_X01_Y00_ready(bit_const_1_None_out),
    .io2glb_1_X01_Y00_valid(Interconnect_inst0_io2glb_1_X01_Y00_valid),
    .io2glb_1_X02_Y00(Interconnect_inst0_io2glb_1_X02_Y00),
    .io2glb_1_X02_Y00_ready(bit_const_1_None_out),
    .io2glb_1_X02_Y00_valid(Interconnect_inst0_io2glb_1_X02_Y00_valid),
    .io2glb_1_X03_Y00(Interconnect_inst0_io2glb_1_X03_Y00),
    .io2glb_1_X03_Y00_ready(bit_const_1_None_out),
    .io2glb_1_X03_Y00_valid(Interconnect_inst0_io2glb_1_X03_Y00_valid),
    .read_config_data(Interconnect_inst0_read_config_data),
    .reset(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_reset_out),
    .stall(global_buffer_W_inst0_cgra_stall)
);
wire [16:0] Interconnect_inst0_glb2io_17_X00_Y00_out;
assign Interconnect_inst0_glb2io_17_X00_Y00_out = {bit_const_0_None_out,global_buffer_W_inst0_strm_data_g2f_0_0};
mantle_wire__typeBitIn17 Interconnect_inst0_glb2io_17_X00_Y00 (
    .in(Interconnect_inst0_glb2io_17_X00_Y00_in),
    .out(Interconnect_inst0_glb2io_17_X00_Y00_out)
);
wire [16:0] Interconnect_inst0_glb2io_17_X01_Y00_out;
assign Interconnect_inst0_glb2io_17_X01_Y00_out = {bit_const_0_None_out,global_buffer_W_inst0_strm_data_g2f_0_1};
mantle_wire__typeBitIn17 Interconnect_inst0_glb2io_17_X01_Y00 (
    .in(Interconnect_inst0_glb2io_17_X01_Y00_in),
    .out(Interconnect_inst0_glb2io_17_X01_Y00_out)
);
wire [16:0] Interconnect_inst0_glb2io_17_X02_Y00_out;
assign Interconnect_inst0_glb2io_17_X02_Y00_out = {bit_const_0_None_out,global_buffer_W_inst0_strm_data_g2f_1_0};
mantle_wire__typeBitIn17 Interconnect_inst0_glb2io_17_X02_Y00 (
    .in(Interconnect_inst0_glb2io_17_X02_Y00_in),
    .out(Interconnect_inst0_glb2io_17_X02_Y00_out)
);
wire [16:0] Interconnect_inst0_glb2io_17_X03_Y00_out;
assign Interconnect_inst0_glb2io_17_X03_Y00_out = {bit_const_0_None_out,global_buffer_W_inst0_strm_data_g2f_1_1};
mantle_wire__typeBitIn17 Interconnect_inst0_glb2io_17_X03_Y00 (
    .in(Interconnect_inst0_glb2io_17_X03_Y00_in),
    .out(Interconnect_inst0_glb2io_17_X03_Y00_out)
);
mantle_wire__typeBit17 Interconnect_inst0_io2glb_17_X00_Y00 (
    .in(Interconnect_inst0_io2glb_17_X00_Y00_unq1),
    .out(Interconnect_inst0_io2glb_17_X00_Y00_out)
);
mantle_wire__typeBit17 Interconnect_inst0_io2glb_17_X01_Y00 (
    .in(Interconnect_inst0_io2glb_17_X01_Y00_unq1),
    .out(Interconnect_inst0_io2glb_17_X01_Y00_out)
);
mantle_wire__typeBit17 Interconnect_inst0_io2glb_17_X02_Y00 (
    .in(Interconnect_inst0_io2glb_17_X02_Y00_unq1),
    .out(Interconnect_inst0_io2glb_17_X02_Y00_out)
);
mantle_wire__typeBit17 Interconnect_inst0_io2glb_17_X03_Y00 (
    .in(Interconnect_inst0_io2glb_17_X03_Y00_unq1),
    .out(Interconnect_inst0_io2glb_17_X03_Y00_out)
);
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
corebit_const #(
    .value(1'b1)
) bit_const_1_None (
    .out(bit_const_1_None_out)
);
global_buffer_W global_buffer_W_inst0 (
    .strm_data_g2f_vld_0_1(global_buffer_W_inst0_strm_data_g2f_vld_0_1),
    .cgra_cfg_g2f_cfg_rd_en_0_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_0_1),
    .reset(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_reset_out),
    .proc_rd_addr(proc_packet_rd_addr),
    .strm_data_g2f_1_1(global_buffer_W_inst0_strm_data_g2f_1_1),
    .proc_wr_strb(proc_packet_wr_strb),
    .if_cfg_wr_data(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_data),
    .strm_data_f2g_vld_1_0(Interconnect_inst0_io2glb_17_X02_Y00_valid),
    .clk(clk_in),
    .cgra_cfg_g2f_cfg_addr_0_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_0_0),
    .if_cfg_wr_clk_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_clk_en),
    .strm_data_f2g_1_0(Interconnect_inst0_io2glb_17_X02_Y00_out[15:0]),
    .proc_wr_addr(proc_packet_wr_addr),
    .strm_data_f2g_vld_0_0(Interconnect_inst0_io2glb_17_X00_Y00_valid),
    .proc_rd_data(global_buffer_W_inst0_proc_rd_data),
    .cgra_cfg_g2f_cfg_addr_0_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_0_1),
    .cgra_cfg_g2f_cfg_data_0_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_0_0),
    .strm_ctrl_f2g_0_1(Interconnect_inst0_io2glb_1_X01_Y00),
    .strm_data_f2g_1_1(Interconnect_inst0_io2glb_17_X03_Y00_out[15:0]),
    .cgra_cfg_g2f_cfg_rd_en_1_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_1_1),
    .strm_data_f2g_0_1(Interconnect_inst0_io2glb_17_X01_Y00_out[15:0]),
    .cgra_stall_in(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_stall),
    .cgra_cfg_jtag_gc2glb_rd_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_read),
    .strm_data_g2f_1_0(global_buffer_W_inst0_strm_data_g2f_1_0),
    .strm_g2f_interrupt_pulse(global_buffer_W_inst0_strm_g2f_interrupt_pulse),
    .if_cfg_rd_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_addr),
    .strm_ctrl_g2f_1_0(global_buffer_W_inst0_strm_ctrl_g2f_1_0),
    .strm_data_g2f_vld_1_0(global_buffer_W_inst0_strm_data_g2f_vld_1_0),
    .strm_data_f2g_0_0(Interconnect_inst0_io2glb_17_X00_Y00_out[15:0]),
    .cgra_cfg_g2f_cfg_wr_en_0_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_0_0),
    .strm_data_g2f_vld_0_0(global_buffer_W_inst0_strm_data_g2f_vld_0_0),
    .flush_crossbar_sel(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_flush_crossbar_sel),
    .cgra_cfg_jtag_gc2glb_wr_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_write),
    .strm_data_f2g_rdy_0_1(global_buffer_W_inst0_strm_data_f2g_rdy_0_1),
    .strm_data_g2f_vld_1_1(global_buffer_W_inst0_strm_data_g2f_vld_1_1),
    .pcfg_broadcast_stall(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_pcfg_broadcast_stall),
    .strm_data_flush_g2f(global_buffer_W_inst0_strm_data_flush_g2f),
    .strm_ctrl_g2f_0_0(global_buffer_W_inst0_strm_ctrl_g2f_0_0),
    .pcfg_start_pulse(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_pc_start_pulse),
    .strm_f2g_start_pulse(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_strm_f2g_start_pulse),
    .cgra_cfg_g2f_cfg_data_1_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_1_0),
    .strm_ctrl_g2f_0_1(global_buffer_W_inst0_strm_ctrl_g2f_0_1),
    .cgra_cfg_g2f_cfg_addr_1_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_1_1),
    .strm_data_f2g_rdy_1_0(global_buffer_W_inst0_strm_data_f2g_rdy_1_0),
    .strm_data_f2g_rdy_0_0(global_buffer_W_inst0_strm_data_f2g_rdy_0_0),
    .cgra_cfg_jtag_gc2glb_data(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_wr_data),
    .strm_ctrl_f2g_1_0(Interconnect_inst0_io2glb_1_X02_Y00),
    .strm_ctrl_g2f_1_1(global_buffer_W_inst0_strm_ctrl_g2f_1_1),
    .if_cfg_wr_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_en),
    .if_cfg_wr_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_wr_addr),
    .if_sram_cfg_rd_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_rd_en),
    .strm_data_g2f_rdy_0_0(Interconnect_inst0_glb2io_17_X00_Y00_ready),
    .cgra_cfg_g2f_cfg_wr_en_1_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_1_1),
    .strm_data_f2g_vld_1_1(Interconnect_inst0_io2glb_17_X03_Y00_valid),
    .if_sram_cfg_rd_data_valid(global_buffer_W_inst0_if_sram_cfg_rd_data_valid),
    .proc_wr_data(proc_packet_wr_data),
    .pcfg_g2f_interrupt_pulse(global_buffer_W_inst0_pcfg_g2f_interrupt_pulse),
    .cgra_cfg_g2f_cfg_data_1_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_1_1),
    .strm_data_f2g_vld_0_1(Interconnect_inst0_io2glb_17_X01_Y00_valid),
    .strm_g2f_start_pulse(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_strm_g2f_start_pulse),
    .strm_data_g2f_rdy_1_1(Interconnect_inst0_glb2io_17_X03_Y00_ready),
    .cgra_cfg_g2f_cfg_data_0_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_data_0_1),
    .proc_rd_en(proc_packet_rd_en),
    .if_cfg_rd_data_valid(global_buffer_W_inst0_if_cfg_rd_data_valid),
    .cgra_stall(global_buffer_W_inst0_cgra_stall),
    .strm_data_g2f_rdy_0_1(Interconnect_inst0_glb2io_17_X01_Y00_ready),
    .strm_ctrl_f2g_1_1(Interconnect_inst0_io2glb_1_X03_Y00),
    .strm_data_g2f_rdy_1_0(Interconnect_inst0_glb2io_17_X02_Y00_ready),
    .if_sram_cfg_rd_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_rd_addr),
    .cgra_cfg_g2f_cfg_addr_1_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_addr_1_0),
    .cgra_cfg_g2f_cfg_rd_en_0_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_0_0),
    .proc_wr_en(proc_packet_wr_en),
    .strm_data_g2f_0_1(global_buffer_W_inst0_strm_data_g2f_0_1),
    .glb_clk_en_master(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_clk_en_master),
    .strm_f2g_interrupt_pulse(global_buffer_W_inst0_strm_f2g_interrupt_pulse),
    .if_sram_cfg_wr_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_addr),
    .if_sram_cfg_rd_data(global_buffer_W_inst0_if_sram_cfg_rd_data),
    .if_sram_cfg_wr_data(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_data),
    .proc_rd_data_valid(global_buffer_W_inst0_proc_rd_data_valid),
    .if_cfg_rd_data(global_buffer_W_inst0_if_cfg_rd_data),
    .strm_ctrl_f2g_0_0(Interconnect_inst0_io2glb_1_X00_Y00),
    .glb_clk_en_bank_master(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_clk_en_bank_master),
    .if_cfg_rd_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_en),
    .strm_data_g2f_0_0(global_buffer_W_inst0_strm_data_g2f_0_0),
    .if_sram_cfg_wr_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_sram_cfg_wr_en),
    .cgra_cfg_g2f_cfg_rd_en_1_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_rd_en_1_0),
    .cgra_cfg_g2f_cfg_wr_en_1_0(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_1_0),
    .strm_data_f2g_rdy_1_1(global_buffer_W_inst0_strm_data_f2g_rdy_1_1),
    .cgra_cfg_jtag_gc2glb_addr(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_cgra_cfg_addr),
    .cgra_cfg_g2f_cfg_wr_en_0_1(global_buffer_W_inst0_cgra_cfg_g2f_cfg_wr_en_0_1),
    .if_cfg_rd_clk_en(GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_glb_cfg_rd_clk_en)
);
assign axi4_slave_arready = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_arready;
assign axi4_slave_awready = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_awready;
assign axi4_slave_bresp = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_bresp;
assign axi4_slave_bvalid = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_bvalid;
assign axi4_slave_rdata = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rdata;
assign axi4_slave_rresp = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rresp;
assign axi4_slave_rvalid = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_rvalid;
assign axi4_slave_wready = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_axi_wready;
assign cgra_running_clk_out = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_clk_out;
assign interrupt = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_interrupt;
assign jtag_tdo = GlobalController_cfg_32_32_axi_13_32_inst0$global_controller_inst0_tdo;
assign proc_packet_rd_data = global_buffer_W_inst0_proc_rd_data;
assign proc_packet_rd_data_valid = global_buffer_W_inst0_proc_rd_data_valid[0];
endmodule

module AN_CELL ( 
input logic  A1, 
input logic  A2, 
output logic  Z); 

`ifdef TSMC16
AN2D0BWP16P90 inst(.A1(A1), .A2(A2), .Z(Z));
`elsif GF12
SC7P5T_AN2X0P5_SSC14R inst(.A(A1), .B(A2), .Z(Z));
`else
assign Z = (A1 & A2); 
`endif

endmodule  
module AO_CELL ( 
input logic  A1,
input logic  A2, 
input logic  B1, 
input logic  B2, 
output logic  Z);  

`ifdef TSMC16
AO22D0BWP16P90 inst(.A1(A1), .A2(A2), .B1(B1), .B2(B2), .Z(Z));
`elsif GF12
SC7P5T_AO22X0P5_SSC14R inst(.A1(A1), .A2(A2), .B1(B1), .B2(B2), .Z(Z));
`else
assign Z = ((A1 & A2) | (B1 & B2)); 
`endif

endmodule 
module PEGEN_coreir_xor #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 ^ in1;
endmodule

module PEGEN_coreir_ule #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = in0 <= in1;
endmodule

module PEGEN_coreir_uge #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = in0 >= in1;
endmodule

module PEGEN_coreir_sle #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = $signed(in0) <= $signed(in1);
endmodule

module PEGEN_coreir_shl #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 << in1;
endmodule

module PEGEN_coreir_sge #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = $signed(in0) >= $signed(in1);
endmodule

module PEGEN_coreir_reg_arst #(
    parameter width = 1,
    parameter arst_posedge = 1,
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input arst,
    input [width-1:0] in,
    output [width-1:0] out
);
  reg [width-1:0] outReg;
  wire real_rst;
  assign real_rst = arst_posedge ? arst : ~arst;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk, posedge real_rst) begin
    if (real_rst) outReg <= init;
    else outReg <= in;
  end
  assign out = outReg;
endmodule

module PEGEN_coreir_or #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 | in1;
endmodule

module PEGEN_coreir_not #(
    parameter width = 1
) (
    input [width-1:0] in,
    output [width-1:0] out
);
  assign out = ~in;
endmodule

module PEGEN_coreir_neg #(
    parameter width = 1
) (
    input [width-1:0] in,
    output [width-1:0] out
);
  assign out = -in;
endmodule

module PEGEN_coreir_mux #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    input sel,
    output [width-1:0] out
);
  assign out = sel ? in1 : in0;
endmodule

module PEGEN_coreir_mul #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 * in1;
endmodule

module PEGEN_coreir_lshr #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 >> in1;
endmodule

module PEGEN_coreir_eq #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = in0 == in1;
endmodule

module PEGEN_coreir_const #(
    parameter width = 1,
    parameter value = 1
) (
    output [width-1:0] out
);
  assign out = value;
endmodule

module PEGEN_coreir_ashr #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = $signed(in0) >>> in1;
endmodule

module PEGEN_coreir_and #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 & in1;
endmodule

module PEGEN_coreir_add #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 + in1;
endmodule

module PEGEN_corebit_xor (
    input in0,
    input in1,
    output out
);
  assign out = in0 ^ in1;
endmodule

module PEGEN_corebit_or (
    input in0,
    input in1,
    output out
);
  assign out = in0 | in1;
endmodule

module PEGEN_corebit_not (
    input in,
    output out
);
  assign out = ~in;
endmodule

module PEGEN_corebit_const #(
    parameter value = 1
) (
    output out
);
  assign out = value;
endmodule

module PEGEN_corebit_and (
    input in0,
    input in1,
    output out
);
  assign out = in0 & in1;
endmodule

module PEGEN_commonlib_muxn__N2__width5 (
    input [4:0] in_data [1:0],
    input [0:0] in_sel,
    output [4:0] out
);
wire [4:0] _join_out;
PEGEN_coreir_mux #(
    .width(5)
) _join (
    .in0(in_data[0]),
    .in1(in_data[1]),
    .sel(in_sel[0]),
    .out(_join_out)
);
assign out = _join_out;
endmodule

module PEGEN_commonlib_muxn__N2__width32 (
    input [31:0] in_data [1:0],
    input [0:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
PEGEN_coreir_mux #(
    .width(32)
) _join (
    .in0(in_data[0]),
    .in1(in_data[1]),
    .sel(in_sel[0]),
    .out(_join_out)
);
assign out = _join_out;
endmodule

module PEGEN_commonlib_muxn__N2__width16 (
    input [15:0] in_data [1:0],
    input [0:0] in_sel,
    output [15:0] out
);
wire [15:0] _join_out;
PEGEN_coreir_mux #(
    .width(16)
) _join (
    .in0(in_data[0]),
    .in1(in_data[1]),
    .sel(in_sel[0]),
    .out(_join_out)
);
assign out = _join_out;
endmodule

module PEGEN_commonlib_muxn__N2__width1 (
    input [0:0] in_data [1:0],
    input [0:0] in_sel,
    output [0:0] out
);
wire [0:0] _join_out;
PEGEN_coreir_mux #(
    .width(1)
) _join (
    .in0(in_data[0]),
    .in1(in_data[1]),
    .sel(in_sel[0]),
    .out(_join_out)
);
assign out = _join_out;
endmodule

module PEGEN_Mux2xUInt32 (
    input [31:0] I0,
    input [31:0] I1,
    input S,
    output [31:0] O
);
wire [31:0] coreir_commonlib_mux2x32_inst0_out;
wire [31:0] coreir_commonlib_mux2x32_inst0_in_data [1:0];
assign coreir_commonlib_mux2x32_inst0_in_data[1] = I1;
assign coreir_commonlib_mux2x32_inst0_in_data[0] = I0;
PEGEN_commonlib_muxn__N2__width32 coreir_commonlib_mux2x32_inst0 (
    .in_data(coreir_commonlib_mux2x32_inst0_in_data),
    .in_sel(S),
    .out(coreir_commonlib_mux2x32_inst0_out)
);
assign O = coreir_commonlib_mux2x32_inst0_out;
endmodule

module PEGEN_Mux2xUInt16 (
    input [15:0] I0,
    input [15:0] I1,
    input S,
    output [15:0] O
);
wire [15:0] coreir_commonlib_mux2x16_inst0_out;
wire [15:0] coreir_commonlib_mux2x16_inst0_in_data [1:0];
assign coreir_commonlib_mux2x16_inst0_in_data[1] = I1;
assign coreir_commonlib_mux2x16_inst0_in_data[0] = I0;
PEGEN_commonlib_muxn__N2__width16 coreir_commonlib_mux2x16_inst0 (
    .in_data(coreir_commonlib_mux2x16_inst0_in_data),
    .in_sel(S),
    .out(coreir_commonlib_mux2x16_inst0_out)
);
assign O = coreir_commonlib_mux2x16_inst0_out;
endmodule

module PEGEN_Mux2xMagmaADTALU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3 (
    input [4:0] I0,
    input [4:0] I1,
    input S,
    output [4:0] O
);
wire [4:0] coreir_commonlib_mux2x5_inst0_out;
wire [4:0] coreir_commonlib_mux2x5_inst0_in_data [1:0];
assign coreir_commonlib_mux2x5_inst0_in_data[1] = I1;
assign coreir_commonlib_mux2x5_inst0_in_data[0] = I0;
PEGEN_commonlib_muxn__N2__width5 coreir_commonlib_mux2x5_inst0 (
    .in_data(coreir_commonlib_mux2x5_inst0_in_data),
    .in_sel(S),
    .out(coreir_commonlib_mux2x5_inst0_out)
);
assign O = coreir_commonlib_mux2x5_inst0_out;
endmodule

module PEGEN_Mux2xBits16 (
    input [15:0] I0,
    input [15:0] I1,
    input S,
    output [15:0] O
);
wire [15:0] coreir_commonlib_mux2x16_inst0_out;
wire [15:0] coreir_commonlib_mux2x16_inst0_in_data [1:0];
assign coreir_commonlib_mux2x16_inst0_in_data[1] = I1;
assign coreir_commonlib_mux2x16_inst0_in_data[0] = I0;
PEGEN_commonlib_muxn__N2__width16 coreir_commonlib_mux2x16_inst0 (
    .in_data(coreir_commonlib_mux2x16_inst0_in_data),
    .in_sel(S),
    .out(coreir_commonlib_mux2x16_inst0_out)
);
assign O = coreir_commonlib_mux2x16_inst0_out;
endmodule

module PEGEN_Register (
    input [15:0] value,
    output [15:0] O,
    input en,
    input CLK,
    input ASYNCRESET
);
wire [15:0] enable_mux_O;
wire [15:0] reg_PR16_inst0_out;
PEGEN_Mux2xBits16 enable_mux (
    .I0(reg_PR16_inst0_out),
    .I1(value),
    .S(en),
    .O(enable_mux_O)
);
PEGEN_coreir_reg_arst #(
    .arst_posedge(1'b1),
    .clk_posedge(1'b1),
    .init(16'h0000),
    .width(16)
) reg_PR16_inst0 (
    .clk(CLK),
    .arst(ASYNCRESET),
    .in(enable_mux_O),
    .out(reg_PR16_inst0_out)
);
assign O = reg_PR16_inst0_out;
endmodule

module PEGEN_Mux2xBit (
    input I0,
    input I1,
    input S,
    output O
);
wire [0:0] coreir_commonlib_mux2x1_inst0_out;
wire [0:0] coreir_commonlib_mux2x1_inst0_in_data [1:0];
assign coreir_commonlib_mux2x1_inst0_in_data[1] = I1;
assign coreir_commonlib_mux2x1_inst0_in_data[0] = I0;
PEGEN_commonlib_muxn__N2__width1 coreir_commonlib_mux2x1_inst0 (
    .in_data(coreir_commonlib_mux2x1_inst0_in_data),
    .in_sel(S),
    .out(coreir_commonlib_mux2x1_inst0_out)
);
assign O = coreir_commonlib_mux2x1_inst0_out[0];
endmodule

module PEGEN_Register_unq1 (
    input value,
    output O,
    input en,
    input CLK,
    input ASYNCRESET
);
wire enable_mux_O;
wire [0:0] reg_PR1_inst0_out;
PEGEN_Mux2xBit enable_mux (
    .I0(reg_PR1_inst0_out[0]),
    .I1(value),
    .S(en),
    .O(enable_mux_O)
);
PEGEN_coreir_reg_arst #(
    .arst_posedge(1'b1),
    .clk_posedge(1'b1),
    .init(1'h0),
    .width(1)
) reg_PR1_inst0 (
    .clk(CLK),
    .arst(ASYNCRESET),
    .in(enable_mux_O),
    .out(reg_PR1_inst0_out)
);
assign O = reg_PR1_inst0_out[0];
endmodule

module PEGEN_RegisterMode_unq1 (
    input [1:0] mode,
    input const_,
    input value,
    input clk_en,
    output O0,
    output O1,
    input CLK,
    input ASYNCRESET
);
wire Mux2xBit_inst0_O;
wire Mux2xBit_inst1_O;
wire Mux2xBit_inst2_O;
wire Mux2xBit_inst3_O;
wire Mux2xBit_inst4_O;
wire Mux2xBit_inst5_O;
wire Register_inst0_O;
wire bit_const_0_None_out;
wire [1:0] const_0_2_out;
wire [1:0] const_2_2_out;
wire [1:0] const_3_2_out;
wire magma_Bits_2_eq_inst0_out;
wire magma_Bits_2_eq_inst1_out;
wire magma_Bits_2_eq_inst2_out;
PEGEN_Mux2xBit Mux2xBit_inst0 (
    .I0(value),
    .I1(value),
    .S(magma_Bits_2_eq_inst0_out),
    .O(Mux2xBit_inst0_O)
);
PEGEN_Mux2xBit Mux2xBit_inst1 (
    .I0(bit_const_0_None_out),
    .I1(clk_en),
    .S(magma_Bits_2_eq_inst0_out),
    .O(Mux2xBit_inst1_O)
);
PEGEN_Mux2xBit Mux2xBit_inst2 (
    .I0(Register_inst0_O),
    .I1(value),
    .S(magma_Bits_2_eq_inst2_out),
    .O(Mux2xBit_inst2_O)
);
PEGEN_Mux2xBit Mux2xBit_inst3 (
    .I0(Register_inst0_O),
    .I1(Register_inst0_O),
    .S(magma_Bits_2_eq_inst2_out),
    .O(Mux2xBit_inst3_O)
);
PEGEN_Mux2xBit Mux2xBit_inst4 (
    .I0(Mux2xBit_inst2_O),
    .I1(const_),
    .S(magma_Bits_2_eq_inst1_out),
    .O(Mux2xBit_inst4_O)
);
PEGEN_Mux2xBit Mux2xBit_inst5 (
    .I0(Mux2xBit_inst3_O),
    .I1(Register_inst0_O),
    .S(magma_Bits_2_eq_inst1_out),
    .O(Mux2xBit_inst5_O)
);
PEGEN_Register_unq1 Register_inst0 (
    .value(Mux2xBit_inst0_O),
    .O(Register_inst0_O),
    .en(Mux2xBit_inst1_O),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
PEGEN_corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
PEGEN_coreir_const #(
    .value(2'h0),
    .width(2)
) const_0_2 (
    .out(const_0_2_out)
);
PEGEN_coreir_const #(
    .value(2'h2),
    .width(2)
) const_2_2 (
    .out(const_2_2_out)
);
PEGEN_coreir_const #(
    .value(2'h3),
    .width(2)
) const_3_2 (
    .out(const_3_2_out)
);
PEGEN_coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst0 (
    .in0(mode),
    .in1(const_3_2_out),
    .out(magma_Bits_2_eq_inst0_out)
);
PEGEN_coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst1 (
    .in0(mode),
    .in1(const_0_2_out),
    .out(magma_Bits_2_eq_inst1_out)
);
PEGEN_coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst2 (
    .in0(mode),
    .in1(const_2_2_out),
    .out(magma_Bits_2_eq_inst2_out)
);
assign O0 = Mux2xBit_inst4_O;
assign O1 = Mux2xBit_inst5_O;
endmodule

module PEGEN_RegisterMode (
    input [1:0] mode,
    input [15:0] const_,
    input [15:0] value,
    input clk_en,
    output [15:0] O0,
    output [15:0] O1,
    input CLK,
    input ASYNCRESET
);
wire Mux2xBit_inst0_O;
wire [15:0] Mux2xBits16_inst0_O;
wire [15:0] Mux2xBits16_inst1_O;
wire [15:0] Mux2xBits16_inst2_O;
wire [15:0] Mux2xBits16_inst3_O;
wire [15:0] Mux2xBits16_inst4_O;
wire [15:0] Register_inst0_O;
wire bit_const_0_None_out;
wire [1:0] const_0_2_out;
wire [1:0] const_2_2_out;
wire [1:0] const_3_2_out;
wire magma_Bits_2_eq_inst0_out;
wire magma_Bits_2_eq_inst1_out;
wire magma_Bits_2_eq_inst2_out;
PEGEN_Mux2xBit Mux2xBit_inst0 (
    .I0(bit_const_0_None_out),
    .I1(clk_en),
    .S(magma_Bits_2_eq_inst0_out),
    .O(Mux2xBit_inst0_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst0 (
    .I0(value),
    .I1(value),
    .S(magma_Bits_2_eq_inst0_out),
    .O(Mux2xBits16_inst0_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst1 (
    .I0(Register_inst0_O),
    .I1(value),
    .S(magma_Bits_2_eq_inst2_out),
    .O(Mux2xBits16_inst1_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst2 (
    .I0(Register_inst0_O),
    .I1(Register_inst0_O),
    .S(magma_Bits_2_eq_inst2_out),
    .O(Mux2xBits16_inst2_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst3 (
    .I0(Mux2xBits16_inst1_O),
    .I1(const_),
    .S(magma_Bits_2_eq_inst1_out),
    .O(Mux2xBits16_inst3_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst4 (
    .I0(Mux2xBits16_inst2_O),
    .I1(Register_inst0_O),
    .S(magma_Bits_2_eq_inst1_out),
    .O(Mux2xBits16_inst4_O)
);
PEGEN_Register Register_inst0 (
    .value(Mux2xBits16_inst0_O),
    .O(Register_inst0_O),
    .en(Mux2xBit_inst0_O),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
PEGEN_corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
PEGEN_coreir_const #(
    .value(2'h0),
    .width(2)
) const_0_2 (
    .out(const_0_2_out)
);
PEGEN_coreir_const #(
    .value(2'h2),
    .width(2)
) const_2_2 (
    .out(const_2_2_out)
);
PEGEN_coreir_const #(
    .value(2'h3),
    .width(2)
) const_3_2 (
    .out(const_3_2_out)
);
PEGEN_coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst0 (
    .in0(mode),
    .in1(const_3_2_out),
    .out(magma_Bits_2_eq_inst0_out)
);
PEGEN_coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst1 (
    .in0(mode),
    .in1(const_0_2_out),
    .out(magma_Bits_2_eq_inst1_out)
);
PEGEN_coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst2 (
    .in0(mode),
    .in1(const_2_2_out),
    .out(magma_Bits_2_eq_inst2_out)
);
assign O0 = Mux2xBits16_inst3_O;
assign O1 = Mux2xBits16_inst4_O;
endmodule

module PEGEN_LUT (
    input [7:0] lut,
    input bit0,
    input bit1,
    input bit2,
    output O,
    input CLK,
    input ASYNCRESET
);
wire bit_const_0_None_out;
wire [7:0] const_1_8_out;
wire [7:0] magma_Bits_8_and_inst0_out;
wire [7:0] magma_Bits_8_lshr_inst0_out;
PEGEN_corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
PEGEN_coreir_const #(
    .value(8'h01),
    .width(8)
) const_1_8 (
    .out(const_1_8_out)
);
PEGEN_coreir_and #(
    .width(8)
) magma_Bits_8_and_inst0 (
    .in0(magma_Bits_8_lshr_inst0_out),
    .in1(const_1_8_out),
    .out(magma_Bits_8_and_inst0_out)
);
wire [7:0] magma_Bits_8_lshr_inst0_in1;
assign magma_Bits_8_lshr_inst0_in1 = {bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit2,bit1,bit0};
PEGEN_coreir_lshr #(
    .width(8)
) magma_Bits_8_lshr_inst0 (
    .in0(lut),
    .in1(magma_Bits_8_lshr_inst0_in1),
    .out(magma_Bits_8_lshr_inst0_out)
);
assign O = magma_Bits_8_and_inst0_out[0];
endmodule

module PEGEN_Cond (
    input [4:0] code,
    input alu,
    input lut,
    input Z,
    input N,
    input C,
    input V,
    output O,
    input CLK,
    input ASYNCRESET
);
wire Mux2xBit_inst0_O;
wire Mux2xBit_inst1_O;
wire Mux2xBit_inst10_O;
wire Mux2xBit_inst11_O;
wire Mux2xBit_inst12_O;
wire Mux2xBit_inst13_O;
wire Mux2xBit_inst14_O;
wire Mux2xBit_inst15_O;
wire Mux2xBit_inst16_O;
wire Mux2xBit_inst17_O;
wire Mux2xBit_inst18_O;
wire Mux2xBit_inst2_O;
wire Mux2xBit_inst3_O;
wire Mux2xBit_inst4_O;
wire Mux2xBit_inst5_O;
wire Mux2xBit_inst6_O;
wire Mux2xBit_inst7_O;
wire Mux2xBit_inst8_O;
wire Mux2xBit_inst9_O;
wire [4:0] const_0_5_out;
wire [4:0] const_10_5_out;
wire [4:0] const_11_5_out;
wire [4:0] const_12_5_out;
wire [4:0] const_13_5_out;
wire [4:0] const_14_5_out;
wire [4:0] const_15_5_out;
wire [4:0] const_16_5_out;
wire [4:0] const_17_5_out;
wire [4:0] const_18_5_out;
wire [4:0] const_1_5_out;
wire [4:0] const_2_5_out;
wire [4:0] const_3_5_out;
wire [4:0] const_4_5_out;
wire [4:0] const_5_5_out;
wire [4:0] const_6_5_out;
wire [4:0] const_7_5_out;
wire [4:0] const_8_5_out;
wire [4:0] const_9_5_out;
wire magma_Bit_and_inst0_out;
wire magma_Bit_and_inst1_out;
wire magma_Bit_and_inst2_out;
wire magma_Bit_and_inst3_out;
wire magma_Bit_not_inst0_out;
wire magma_Bit_not_inst1_out;
wire magma_Bit_not_inst10_out;
wire magma_Bit_not_inst11_out;
wire magma_Bit_not_inst12_out;
wire magma_Bit_not_inst2_out;
wire magma_Bit_not_inst3_out;
wire magma_Bit_not_inst4_out;
wire magma_Bit_not_inst5_out;
wire magma_Bit_not_inst6_out;
wire magma_Bit_not_inst7_out;
wire magma_Bit_not_inst8_out;
wire magma_Bit_not_inst9_out;
wire magma_Bit_or_inst0_out;
wire magma_Bit_or_inst1_out;
wire magma_Bit_or_inst2_out;
wire magma_Bit_or_inst3_out;
wire magma_Bit_or_inst4_out;
wire magma_Bit_or_inst5_out;
wire magma_Bit_xor_inst0_out;
wire magma_Bit_xor_inst1_out;
wire magma_Bit_xor_inst2_out;
wire magma_Bit_xor_inst3_out;
wire magma_Bits_5_eq_inst0_out;
wire magma_Bits_5_eq_inst1_out;
wire magma_Bits_5_eq_inst10_out;
wire magma_Bits_5_eq_inst11_out;
wire magma_Bits_5_eq_inst12_out;
wire magma_Bits_5_eq_inst13_out;
wire magma_Bits_5_eq_inst14_out;
wire magma_Bits_5_eq_inst15_out;
wire magma_Bits_5_eq_inst16_out;
wire magma_Bits_5_eq_inst17_out;
wire magma_Bits_5_eq_inst18_out;
wire magma_Bits_5_eq_inst19_out;
wire magma_Bits_5_eq_inst2_out;
wire magma_Bits_5_eq_inst20_out;
wire magma_Bits_5_eq_inst3_out;
wire magma_Bits_5_eq_inst4_out;
wire magma_Bits_5_eq_inst5_out;
wire magma_Bits_5_eq_inst6_out;
wire magma_Bits_5_eq_inst7_out;
wire magma_Bits_5_eq_inst8_out;
wire magma_Bits_5_eq_inst9_out;
PEGEN_Mux2xBit Mux2xBit_inst0 (
    .I0(magma_Bit_and_inst3_out),
    .I1(magma_Bit_or_inst5_out),
    .S(magma_Bits_5_eq_inst20_out),
    .O(Mux2xBit_inst0_O)
);
PEGEN_Mux2xBit Mux2xBit_inst1 (
    .I0(Mux2xBit_inst0_O),
    .I1(magma_Bit_and_inst2_out),
    .S(magma_Bits_5_eq_inst19_out),
    .O(Mux2xBit_inst1_O)
);
PEGEN_Mux2xBit Mux2xBit_inst10 (
    .I0(Mux2xBit_inst9_O),
    .I1(magma_Bit_and_inst0_out),
    .S(magma_Bits_5_eq_inst10_out),
    .O(Mux2xBit_inst10_O)
);
PEGEN_Mux2xBit Mux2xBit_inst11 (
    .I0(Mux2xBit_inst10_O),
    .I1(magma_Bit_not_inst3_out),
    .S(magma_Bits_5_eq_inst9_out),
    .O(Mux2xBit_inst11_O)
);
PEGEN_Mux2xBit Mux2xBit_inst12 (
    .I0(Mux2xBit_inst11_O),
    .I1(V),
    .S(magma_Bits_5_eq_inst8_out),
    .O(Mux2xBit_inst12_O)
);
PEGEN_Mux2xBit Mux2xBit_inst13 (
    .I0(Mux2xBit_inst12_O),
    .I1(magma_Bit_not_inst2_out),
    .S(magma_Bits_5_eq_inst7_out),
    .O(Mux2xBit_inst13_O)
);
PEGEN_Mux2xBit Mux2xBit_inst14 (
    .I0(Mux2xBit_inst13_O),
    .I1(N),
    .S(magma_Bits_5_eq_inst6_out),
    .O(Mux2xBit_inst14_O)
);
PEGEN_Mux2xBit Mux2xBit_inst15 (
    .I0(Mux2xBit_inst14_O),
    .I1(magma_Bit_not_inst1_out),
    .S(magma_Bit_or_inst1_out),
    .O(Mux2xBit_inst15_O)
);
PEGEN_Mux2xBit Mux2xBit_inst16 (
    .I0(Mux2xBit_inst15_O),
    .I1(C),
    .S(magma_Bit_or_inst0_out),
    .O(Mux2xBit_inst16_O)
);
PEGEN_Mux2xBit Mux2xBit_inst17 (
    .I0(Mux2xBit_inst16_O),
    .I1(magma_Bit_not_inst0_out),
    .S(magma_Bits_5_eq_inst1_out),
    .O(Mux2xBit_inst17_O)
);
PEGEN_Mux2xBit Mux2xBit_inst18 (
    .I0(Mux2xBit_inst17_O),
    .I1(Z),
    .S(magma_Bits_5_eq_inst0_out),
    .O(Mux2xBit_inst18_O)
);
PEGEN_Mux2xBit Mux2xBit_inst2 (
    .I0(Mux2xBit_inst1_O),
    .I1(magma_Bit_or_inst4_out),
    .S(magma_Bits_5_eq_inst18_out),
    .O(Mux2xBit_inst2_O)
);
PEGEN_Mux2xBit Mux2xBit_inst3 (
    .I0(Mux2xBit_inst2_O),
    .I1(lut),
    .S(magma_Bits_5_eq_inst17_out),
    .O(Mux2xBit_inst3_O)
);
PEGEN_Mux2xBit Mux2xBit_inst4 (
    .I0(Mux2xBit_inst3_O),
    .I1(alu),
    .S(magma_Bits_5_eq_inst16_out),
    .O(Mux2xBit_inst4_O)
);
PEGEN_Mux2xBit Mux2xBit_inst5 (
    .I0(Mux2xBit_inst4_O),
    .I1(magma_Bit_or_inst3_out),
    .S(magma_Bits_5_eq_inst15_out),
    .O(Mux2xBit_inst5_O)
);
PEGEN_Mux2xBit Mux2xBit_inst6 (
    .I0(Mux2xBit_inst5_O),
    .I1(magma_Bit_and_inst1_out),
    .S(magma_Bits_5_eq_inst14_out),
    .O(Mux2xBit_inst6_O)
);
PEGEN_Mux2xBit Mux2xBit_inst7 (
    .I0(Mux2xBit_inst6_O),
    .I1(magma_Bit_xor_inst1_out),
    .S(magma_Bits_5_eq_inst13_out),
    .O(Mux2xBit_inst7_O)
);
PEGEN_Mux2xBit Mux2xBit_inst8 (
    .I0(Mux2xBit_inst7_O),
    .I1(magma_Bit_not_inst6_out),
    .S(magma_Bits_5_eq_inst12_out),
    .O(Mux2xBit_inst8_O)
);
PEGEN_Mux2xBit Mux2xBit_inst9 (
    .I0(Mux2xBit_inst8_O),
    .I1(magma_Bit_or_inst2_out),
    .S(magma_Bits_5_eq_inst11_out),
    .O(Mux2xBit_inst9_O)
);
PEGEN_coreir_const #(
    .value(5'h00),
    .width(5)
) const_0_5 (
    .out(const_0_5_out)
);
PEGEN_coreir_const #(
    .value(5'h0a),
    .width(5)
) const_10_5 (
    .out(const_10_5_out)
);
PEGEN_coreir_const #(
    .value(5'h0b),
    .width(5)
) const_11_5 (
    .out(const_11_5_out)
);
PEGEN_coreir_const #(
    .value(5'h0c),
    .width(5)
) const_12_5 (
    .out(const_12_5_out)
);
PEGEN_coreir_const #(
    .value(5'h0d),
    .width(5)
) const_13_5 (
    .out(const_13_5_out)
);
PEGEN_coreir_const #(
    .value(5'h0e),
    .width(5)
) const_14_5 (
    .out(const_14_5_out)
);
PEGEN_coreir_const #(
    .value(5'h0f),
    .width(5)
) const_15_5 (
    .out(const_15_5_out)
);
PEGEN_coreir_const #(
    .value(5'h10),
    .width(5)
) const_16_5 (
    .out(const_16_5_out)
);
PEGEN_coreir_const #(
    .value(5'h11),
    .width(5)
) const_17_5 (
    .out(const_17_5_out)
);
PEGEN_coreir_const #(
    .value(5'h12),
    .width(5)
) const_18_5 (
    .out(const_18_5_out)
);
PEGEN_coreir_const #(
    .value(5'h01),
    .width(5)
) const_1_5 (
    .out(const_1_5_out)
);
PEGEN_coreir_const #(
    .value(5'h02),
    .width(5)
) const_2_5 (
    .out(const_2_5_out)
);
PEGEN_coreir_const #(
    .value(5'h03),
    .width(5)
) const_3_5 (
    .out(const_3_5_out)
);
PEGEN_coreir_const #(
    .value(5'h04),
    .width(5)
) const_4_5 (
    .out(const_4_5_out)
);
PEGEN_coreir_const #(
    .value(5'h05),
    .width(5)
) const_5_5 (
    .out(const_5_5_out)
);
PEGEN_coreir_const #(
    .value(5'h06),
    .width(5)
) const_6_5 (
    .out(const_6_5_out)
);
PEGEN_coreir_const #(
    .value(5'h07),
    .width(5)
) const_7_5 (
    .out(const_7_5_out)
);
PEGEN_coreir_const #(
    .value(5'h08),
    .width(5)
) const_8_5 (
    .out(const_8_5_out)
);
PEGEN_coreir_const #(
    .value(5'h09),
    .width(5)
) const_9_5 (
    .out(const_9_5_out)
);
PEGEN_corebit_and magma_Bit_and_inst0 (
    .in0(C),
    .in1(magma_Bit_not_inst4_out),
    .out(magma_Bit_and_inst0_out)
);
PEGEN_corebit_and magma_Bit_and_inst1 (
    .in0(magma_Bit_not_inst7_out),
    .in1(magma_Bit_not_inst8_out),
    .out(magma_Bit_and_inst1_out)
);
PEGEN_corebit_and magma_Bit_and_inst2 (
    .in0(magma_Bit_not_inst10_out),
    .in1(magma_Bit_not_inst11_out),
    .out(magma_Bit_and_inst2_out)
);
PEGEN_corebit_and magma_Bit_and_inst3 (
    .in0(N),
    .in1(magma_Bit_not_inst12_out),
    .out(magma_Bit_and_inst3_out)
);
PEGEN_corebit_not magma_Bit_not_inst0 (
    .in(Z),
    .out(magma_Bit_not_inst0_out)
);
PEGEN_corebit_not magma_Bit_not_inst1 (
    .in(C),
    .out(magma_Bit_not_inst1_out)
);
PEGEN_corebit_not magma_Bit_not_inst10 (
    .in(N),
    .out(magma_Bit_not_inst10_out)
);
PEGEN_corebit_not magma_Bit_not_inst11 (
    .in(Z),
    .out(magma_Bit_not_inst11_out)
);
PEGEN_corebit_not magma_Bit_not_inst12 (
    .in(Z),
    .out(magma_Bit_not_inst12_out)
);
PEGEN_corebit_not magma_Bit_not_inst2 (
    .in(N),
    .out(magma_Bit_not_inst2_out)
);
PEGEN_corebit_not magma_Bit_not_inst3 (
    .in(V),
    .out(magma_Bit_not_inst3_out)
);
PEGEN_corebit_not magma_Bit_not_inst4 (
    .in(Z),
    .out(magma_Bit_not_inst4_out)
);
PEGEN_corebit_not magma_Bit_not_inst5 (
    .in(C),
    .out(magma_Bit_not_inst5_out)
);
PEGEN_corebit_not magma_Bit_not_inst6 (
    .in(magma_Bit_xor_inst0_out),
    .out(magma_Bit_not_inst6_out)
);
PEGEN_corebit_not magma_Bit_not_inst7 (
    .in(Z),
    .out(magma_Bit_not_inst7_out)
);
PEGEN_corebit_not magma_Bit_not_inst8 (
    .in(magma_Bit_xor_inst2_out),
    .out(magma_Bit_not_inst8_out)
);
PEGEN_corebit_not magma_Bit_not_inst9 (
    .in(N),
    .out(magma_Bit_not_inst9_out)
);
PEGEN_corebit_or magma_Bit_or_inst0 (
    .in0(magma_Bits_5_eq_inst2_out),
    .in1(magma_Bits_5_eq_inst3_out),
    .out(magma_Bit_or_inst0_out)
);
PEGEN_corebit_or magma_Bit_or_inst1 (
    .in0(magma_Bits_5_eq_inst4_out),
    .in1(magma_Bits_5_eq_inst5_out),
    .out(magma_Bit_or_inst1_out)
);
PEGEN_corebit_or magma_Bit_or_inst2 (
    .in0(magma_Bit_not_inst5_out),
    .in1(Z),
    .out(magma_Bit_or_inst2_out)
);
PEGEN_corebit_or magma_Bit_or_inst3 (
    .in0(Z),
    .in1(magma_Bit_xor_inst3_out),
    .out(magma_Bit_or_inst3_out)
);
PEGEN_corebit_or magma_Bit_or_inst4 (
    .in0(magma_Bit_not_inst9_out),
    .in1(Z),
    .out(magma_Bit_or_inst4_out)
);
PEGEN_corebit_or magma_Bit_or_inst5 (
    .in0(N),
    .in1(Z),
    .out(magma_Bit_or_inst5_out)
);
PEGEN_corebit_xor magma_Bit_xor_inst0 (
    .in0(N),
    .in1(V),
    .out(magma_Bit_xor_inst0_out)
);
PEGEN_corebit_xor magma_Bit_xor_inst1 (
    .in0(N),
    .in1(V),
    .out(magma_Bit_xor_inst1_out)
);
PEGEN_corebit_xor magma_Bit_xor_inst2 (
    .in0(N),
    .in1(V),
    .out(magma_Bit_xor_inst2_out)
);
PEGEN_corebit_xor magma_Bit_xor_inst3 (
    .in0(N),
    .in1(V),
    .out(magma_Bit_xor_inst3_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst0 (
    .in0(code),
    .in1(const_0_5_out),
    .out(magma_Bits_5_eq_inst0_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst1 (
    .in0(code),
    .in1(const_1_5_out),
    .out(magma_Bits_5_eq_inst1_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst10 (
    .in0(code),
    .in1(const_8_5_out),
    .out(magma_Bits_5_eq_inst10_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst11 (
    .in0(code),
    .in1(const_9_5_out),
    .out(magma_Bits_5_eq_inst11_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst12 (
    .in0(code),
    .in1(const_10_5_out),
    .out(magma_Bits_5_eq_inst12_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst13 (
    .in0(code),
    .in1(const_11_5_out),
    .out(magma_Bits_5_eq_inst13_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst14 (
    .in0(code),
    .in1(const_12_5_out),
    .out(magma_Bits_5_eq_inst14_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst15 (
    .in0(code),
    .in1(const_13_5_out),
    .out(magma_Bits_5_eq_inst15_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst16 (
    .in0(code),
    .in1(const_15_5_out),
    .out(magma_Bits_5_eq_inst16_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst17 (
    .in0(code),
    .in1(const_14_5_out),
    .out(magma_Bits_5_eq_inst17_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst18 (
    .in0(code),
    .in1(const_16_5_out),
    .out(magma_Bits_5_eq_inst18_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst19 (
    .in0(code),
    .in1(const_17_5_out),
    .out(magma_Bits_5_eq_inst19_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst2 (
    .in0(code),
    .in1(const_2_5_out),
    .out(magma_Bits_5_eq_inst2_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst20 (
    .in0(code),
    .in1(const_18_5_out),
    .out(magma_Bits_5_eq_inst20_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst3 (
    .in0(code),
    .in1(const_2_5_out),
    .out(magma_Bits_5_eq_inst3_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst4 (
    .in0(code),
    .in1(const_3_5_out),
    .out(magma_Bits_5_eq_inst4_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst5 (
    .in0(code),
    .in1(const_3_5_out),
    .out(magma_Bits_5_eq_inst5_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst6 (
    .in0(code),
    .in1(const_4_5_out),
    .out(magma_Bits_5_eq_inst6_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst7 (
    .in0(code),
    .in1(const_5_5_out),
    .out(magma_Bits_5_eq_inst7_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst8 (
    .in0(code),
    .in1(const_6_5_out),
    .out(magma_Bits_5_eq_inst8_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst9 (
    .in0(code),
    .in1(const_7_5_out),
    .out(magma_Bits_5_eq_inst9_out)
);
assign O = Mux2xBit_inst18_O;
endmodule

module PEGEN_ALU (
    input [4:0] alu,
    input [0:0] signed_,
    input [15:0] a,
    input [15:0] b,
    input [15:0] c,
    input d,
    output [15:0] res,
    output res_p,
    output Z,
    output N,
    output C,
    output V,
    input CLK,
    input ASYNCRESET
);
wire Mux2xBit_inst0_O;
wire Mux2xBit_inst1_O;
wire Mux2xBit_inst10_O;
wire Mux2xBit_inst11_O;
wire Mux2xBit_inst12_O;
wire Mux2xBit_inst13_O;
wire Mux2xBit_inst14_O;
wire Mux2xBit_inst15_O;
wire Mux2xBit_inst16_O;
wire Mux2xBit_inst17_O;
wire Mux2xBit_inst18_O;
wire Mux2xBit_inst19_O;
wire Mux2xBit_inst2_O;
wire Mux2xBit_inst20_O;
wire Mux2xBit_inst21_O;
wire Mux2xBit_inst22_O;
wire Mux2xBit_inst23_O;
wire Mux2xBit_inst3_O;
wire Mux2xBit_inst4_O;
wire Mux2xBit_inst5_O;
wire Mux2xBit_inst6_O;
wire Mux2xBit_inst7_O;
wire Mux2xBit_inst8_O;
wire Mux2xBit_inst9_O;
wire [15:0] Mux2xBits16_inst0_O;
wire [15:0] Mux2xBits16_inst1_O;
wire [15:0] Mux2xBits16_inst10_O;
wire [15:0] Mux2xBits16_inst11_O;
wire [15:0] Mux2xBits16_inst12_O;
wire [15:0] Mux2xBits16_inst13_O;
wire [15:0] Mux2xBits16_inst14_O;
wire [15:0] Mux2xBits16_inst15_O;
wire [15:0] Mux2xBits16_inst16_O;
wire [15:0] Mux2xBits16_inst17_O;
wire [15:0] Mux2xBits16_inst18_O;
wire [15:0] Mux2xBits16_inst19_O;
wire [15:0] Mux2xBits16_inst2_O;
wire [15:0] Mux2xBits16_inst20_O;
wire [15:0] Mux2xBits16_inst21_O;
wire [15:0] Mux2xBits16_inst3_O;
wire [15:0] Mux2xBits16_inst4_O;
wire [15:0] Mux2xBits16_inst5_O;
wire [15:0] Mux2xBits16_inst6_O;
wire [15:0] Mux2xBits16_inst7_O;
wire [15:0] Mux2xBits16_inst8_O;
wire [15:0] Mux2xBits16_inst9_O;
wire [15:0] Mux2xUInt16_inst0_O;
wire [31:0] Mux2xUInt32_inst0_O;
wire [31:0] Mux2xUInt32_inst1_O;
wire bit_const_0_None_out;
wire bit_const_1_None_out;
wire [15:0] const_0_16_out;
wire [4:0] const_0_5_out;
wire [4:0] const_10_5_out;
wire [4:0] const_11_5_out;
wire [4:0] const_12_5_out;
wire [4:0] const_13_5_out;
wire [4:0] const_14_5_out;
wire [4:0] const_15_5_out;
wire [4:0] const_16_5_out;
wire [4:0] const_17_5_out;
wire [4:0] const_18_5_out;
wire [4:0] const_19_5_out;
wire [0:0] const_1_1_out;
wire [4:0] const_1_5_out;
wire [4:0] const_2_5_out;
wire [4:0] const_3_5_out;
wire [4:0] const_4_5_out;
wire [4:0] const_5_5_out;
wire [4:0] const_6_5_out;
wire [4:0] const_7_5_out;
wire [4:0] const_8_5_out;
wire [4:0] const_9_5_out;
wire magma_Bit_and_inst0_out;
wire magma_Bit_and_inst1_out;
wire magma_Bit_and_inst2_out;
wire magma_Bit_and_inst3_out;
wire magma_Bit_not_inst0_out;
wire magma_Bit_not_inst1_out;
wire magma_Bit_not_inst2_out;
wire magma_Bit_or_inst0_out;
wire magma_Bit_or_inst1_out;
wire magma_Bit_or_inst10_out;
wire magma_Bit_or_inst11_out;
wire magma_Bit_or_inst12_out;
wire magma_Bit_or_inst13_out;
wire magma_Bit_or_inst2_out;
wire magma_Bit_or_inst3_out;
wire magma_Bit_or_inst4_out;
wire magma_Bit_or_inst5_out;
wire magma_Bit_or_inst6_out;
wire magma_Bit_or_inst7_out;
wire magma_Bit_or_inst8_out;
wire magma_Bit_or_inst9_out;
wire [15:0] magma_Bits_16_and_inst0_out;
wire [15:0] magma_Bits_16_not_inst0_out;
wire [15:0] magma_Bits_16_not_inst1_out;
wire [15:0] magma_Bits_16_or_inst0_out;
wire [15:0] magma_Bits_16_shl_inst0_out;
wire [15:0] magma_Bits_16_xor_inst0_out;
wire magma_Bits_1_eq_inst0_out;
wire magma_Bits_1_eq_inst1_out;
wire magma_Bits_1_eq_inst2_out;
wire magma_Bits_1_eq_inst3_out;
wire magma_Bits_5_eq_inst0_out;
wire magma_Bits_5_eq_inst1_out;
wire magma_Bits_5_eq_inst10_out;
wire magma_Bits_5_eq_inst11_out;
wire magma_Bits_5_eq_inst12_out;
wire magma_Bits_5_eq_inst13_out;
wire magma_Bits_5_eq_inst14_out;
wire magma_Bits_5_eq_inst15_out;
wire magma_Bits_5_eq_inst16_out;
wire magma_Bits_5_eq_inst17_out;
wire magma_Bits_5_eq_inst18_out;
wire magma_Bits_5_eq_inst19_out;
wire magma_Bits_5_eq_inst2_out;
wire magma_Bits_5_eq_inst20_out;
wire magma_Bits_5_eq_inst21_out;
wire magma_Bits_5_eq_inst22_out;
wire magma_Bits_5_eq_inst23_out;
wire magma_Bits_5_eq_inst24_out;
wire magma_Bits_5_eq_inst25_out;
wire magma_Bits_5_eq_inst26_out;
wire magma_Bits_5_eq_inst27_out;
wire magma_Bits_5_eq_inst28_out;
wire magma_Bits_5_eq_inst29_out;
wire magma_Bits_5_eq_inst3_out;
wire magma_Bits_5_eq_inst30_out;
wire magma_Bits_5_eq_inst4_out;
wire magma_Bits_5_eq_inst5_out;
wire magma_Bits_5_eq_inst6_out;
wire magma_Bits_5_eq_inst7_out;
wire magma_Bits_5_eq_inst8_out;
wire magma_Bits_5_eq_inst9_out;
wire [15:0] magma_SInt_16_ashr_inst0_out;
wire magma_SInt_16_eq_inst0_out;
wire [15:0] magma_SInt_16_neg_inst0_out;
wire magma_SInt_16_sge_inst0_out;
wire magma_SInt_16_sle_inst0_out;
wire magma_SInt_16_sle_inst1_out;
wire [15:0] magma_UInt_16_lshr_inst0_out;
wire magma_UInt_16_uge_inst0_out;
wire magma_UInt_16_ule_inst0_out;
wire [16:0] magma_UInt_17_add_inst0_out;
wire [16:0] magma_UInt_17_add_inst1_out;
wire [16:0] magma_UInt_17_add_inst2_out;
wire [16:0] magma_UInt_17_add_inst3_out;
wire [31:0] magma_UInt_32_mul_inst0_out;
PEGEN_Mux2xBit Mux2xBit_inst0 (
    .I0(magma_UInt_16_ule_inst0_out),
    .I1(magma_SInt_16_sle_inst0_out),
    .S(magma_Bits_1_eq_inst1_out),
    .O(Mux2xBit_inst0_O)
);
PEGEN_Mux2xBit Mux2xBit_inst1 (
    .I0(magma_UInt_16_uge_inst0_out),
    .I1(magma_SInt_16_sge_inst0_out),
    .S(magma_Bits_1_eq_inst2_out),
    .O(Mux2xBit_inst1_O)
);
PEGEN_Mux2xBit Mux2xBit_inst10 (
    .I0(Mux2xBit_inst9_O),
    .I1(bit_const_0_None_out),
    .S(magma_Bits_5_eq_inst18_out),
    .O(Mux2xBit_inst10_O)
);
PEGEN_Mux2xBit Mux2xBit_inst11 (
    .I0(Mux2xBit_inst10_O),
    .I1(a[15]),
    .S(magma_Bits_5_eq_inst17_out),
    .O(Mux2xBit_inst11_O)
);
PEGEN_Mux2xBit Mux2xBit_inst12 (
    .I0(bit_const_0_None_out),
    .I1(bit_const_0_None_out),
    .S(magma_Bits_5_eq_inst16_out),
    .O(Mux2xBit_inst12_O)
);
PEGEN_Mux2xBit Mux2xBit_inst13 (
    .I0(bit_const_0_None_out),
    .I1(bit_const_0_None_out),
    .S(magma_Bits_5_eq_inst16_out),
    .O(Mux2xBit_inst13_O)
);
PEGEN_Mux2xBit Mux2xBit_inst14 (
    .I0(Mux2xBit_inst11_O),
    .I1(bit_const_0_None_out),
    .S(magma_Bits_5_eq_inst16_out),
    .O(Mux2xBit_inst14_O)
);
PEGEN_Mux2xBit Mux2xBit_inst15 (
    .I0(Mux2xBit_inst12_O),
    .I1(bit_const_0_None_out),
    .S(magma_Bits_5_eq_inst15_out),
    .O(Mux2xBit_inst15_O)
);
PEGEN_Mux2xBit Mux2xBit_inst16 (
    .I0(Mux2xBit_inst13_O),
    .I1(bit_const_0_None_out),
    .S(magma_Bits_5_eq_inst15_out),
    .O(Mux2xBit_inst16_O)
);
PEGEN_Mux2xBit Mux2xBit_inst17 (
    .I0(Mux2xBit_inst14_O),
    .I1(bit_const_0_None_out),
    .S(magma_Bits_5_eq_inst15_out),
    .O(Mux2xBit_inst17_O)
);
PEGEN_Mux2xBit Mux2xBit_inst18 (
    .I0(Mux2xBit_inst15_O),
    .I1(bit_const_0_None_out),
    .S(magma_Bits_5_eq_inst14_out),
    .O(Mux2xBit_inst18_O)
);
PEGEN_Mux2xBit Mux2xBit_inst19 (
    .I0(Mux2xBit_inst16_O),
    .I1(bit_const_0_None_out),
    .S(magma_Bits_5_eq_inst14_out),
    .O(Mux2xBit_inst19_O)
);
PEGEN_Mux2xBit Mux2xBit_inst2 (
    .I0(bit_const_0_None_out),
    .I1(bit_const_1_None_out),
    .S(magma_Bit_or_inst6_out),
    .O(Mux2xBit_inst2_O)
);
PEGEN_Mux2xBit Mux2xBit_inst20 (
    .I0(Mux2xBit_inst17_O),
    .I1(bit_const_0_None_out),
    .S(magma_Bits_5_eq_inst14_out),
    .O(Mux2xBit_inst20_O)
);
PEGEN_Mux2xBit Mux2xBit_inst21 (
    .I0(Mux2xBit_inst18_O),
    .I1(magma_UInt_17_add_inst1_out[16]),
    .S(magma_Bit_or_inst7_out),
    .O(Mux2xBit_inst21_O)
);
PEGEN_Mux2xBit Mux2xBit_inst22 (
    .I0(Mux2xBit_inst19_O),
    .I1(magma_Bit_or_inst8_out),
    .S(magma_Bit_or_inst7_out),
    .O(Mux2xBit_inst22_O)
);
PEGEN_Mux2xBit Mux2xBit_inst23 (
    .I0(Mux2xBit_inst20_O),
    .I1(magma_UInt_17_add_inst1_out[16]),
    .S(magma_Bit_or_inst7_out),
    .O(Mux2xBit_inst23_O)
);
PEGEN_Mux2xBit Mux2xBit_inst3 (
    .I0(bit_const_0_None_out),
    .I1(bit_const_0_None_out),
    .S(magma_Bits_5_eq_inst30_out),
    .O(Mux2xBit_inst3_O)
);
PEGEN_Mux2xBit Mux2xBit_inst4 (
    .I0(Mux2xBit_inst3_O),
    .I1(bit_const_0_None_out),
    .S(magma_Bit_or_inst13_out),
    .O(Mux2xBit_inst4_O)
);
PEGEN_Mux2xBit Mux2xBit_inst5 (
    .I0(Mux2xBit_inst4_O),
    .I1(bit_const_0_None_out),
    .S(magma_Bits_5_eq_inst23_out),
    .O(Mux2xBit_inst5_O)
);
PEGEN_Mux2xBit Mux2xBit_inst6 (
    .I0(Mux2xBit_inst5_O),
    .I1(bit_const_0_None_out),
    .S(magma_Bits_5_eq_inst22_out),
    .O(Mux2xBit_inst6_O)
);
PEGEN_Mux2xBit Mux2xBit_inst7 (
    .I0(Mux2xBit_inst6_O),
    .I1(bit_const_0_None_out),
    .S(magma_Bits_5_eq_inst21_out),
    .O(Mux2xBit_inst7_O)
);
PEGEN_Mux2xBit Mux2xBit_inst8 (
    .I0(Mux2xBit_inst7_O),
    .I1(bit_const_0_None_out),
    .S(magma_Bits_5_eq_inst20_out),
    .O(Mux2xBit_inst8_O)
);
PEGEN_Mux2xBit Mux2xBit_inst9 (
    .I0(Mux2xBit_inst8_O),
    .I1(bit_const_0_None_out),
    .S(magma_Bits_5_eq_inst19_out),
    .O(Mux2xBit_inst9_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst0 (
    .I0(b),
    .I1(a),
    .S(Mux2xBit_inst0_O),
    .O(Mux2xBits16_inst0_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst1 (
    .I0(b),
    .I1(Mux2xBits16_inst0_O),
    .S(magma_Bits_5_eq_inst0_out),
    .O(Mux2xBits16_inst1_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst10 (
    .I0(Mux2xBits16_inst9_O),
    .I1(magma_UInt_17_add_inst3_out[15:0]),
    .S(magma_Bit_or_inst13_out),
    .O(Mux2xBits16_inst10_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst11 (
    .I0(Mux2xBits16_inst10_O),
    .I1(magma_Bits_16_shl_inst0_out),
    .S(magma_Bits_5_eq_inst23_out),
    .O(Mux2xBits16_inst11_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst12 (
    .I0(Mux2xBits16_inst11_O),
    .I1(Mux2xBits16_inst4_O),
    .S(magma_Bits_5_eq_inst22_out),
    .O(Mux2xBits16_inst12_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst13 (
    .I0(Mux2xBits16_inst12_O),
    .I1(magma_Bits_16_xor_inst0_out),
    .S(magma_Bits_5_eq_inst21_out),
    .O(Mux2xBits16_inst13_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst14 (
    .I0(Mux2xBits16_inst13_O),
    .I1(magma_Bits_16_or_inst0_out),
    .S(magma_Bits_5_eq_inst20_out),
    .O(Mux2xBits16_inst14_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst15 (
    .I0(Mux2xBits16_inst14_O),
    .I1(magma_Bits_16_and_inst0_out),
    .S(magma_Bits_5_eq_inst19_out),
    .O(Mux2xBits16_inst15_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst16 (
    .I0(Mux2xBits16_inst15_O),
    .I1(Mux2xBits16_inst8_O),
    .S(magma_Bits_5_eq_inst18_out),
    .O(Mux2xBits16_inst16_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst17 (
    .I0(Mux2xBits16_inst16_O),
    .I1(Mux2xBits16_inst7_O),
    .S(magma_Bits_5_eq_inst17_out),
    .O(Mux2xBits16_inst17_O)
);
wire [15:0] Mux2xBits16_inst18_I1;
assign Mux2xBits16_inst18_I1 = {magma_UInt_32_mul_inst0_out[31],magma_UInt_32_mul_inst0_out[30],magma_UInt_32_mul_inst0_out[29],magma_UInt_32_mul_inst0_out[28],magma_UInt_32_mul_inst0_out[27],magma_UInt_32_mul_inst0_out[26],magma_UInt_32_mul_inst0_out[25],magma_UInt_32_mul_inst0_out[24],magma_UInt_32_mul_inst0_out[23],magma_UInt_32_mul_inst0_out[22],magma_UInt_32_mul_inst0_out[21],magma_UInt_32_mul_inst0_out[20],magma_UInt_32_mul_inst0_out[19],magma_UInt_32_mul_inst0_out[18],magma_UInt_32_mul_inst0_out[17],magma_UInt_32_mul_inst0_out[16]};
PEGEN_Mux2xBits16 Mux2xBits16_inst18 (
    .I0(Mux2xBits16_inst17_O),
    .I1(Mux2xBits16_inst18_I1),
    .S(magma_Bits_5_eq_inst16_out),
    .O(Mux2xBits16_inst18_O)
);
wire [15:0] Mux2xBits16_inst19_I1;
assign Mux2xBits16_inst19_I1 = {magma_UInt_32_mul_inst0_out[23],magma_UInt_32_mul_inst0_out[22],magma_UInt_32_mul_inst0_out[21],magma_UInt_32_mul_inst0_out[20],magma_UInt_32_mul_inst0_out[19],magma_UInt_32_mul_inst0_out[18],magma_UInt_32_mul_inst0_out[17],magma_UInt_32_mul_inst0_out[16],magma_UInt_32_mul_inst0_out[15],magma_UInt_32_mul_inst0_out[14],magma_UInt_32_mul_inst0_out[13],magma_UInt_32_mul_inst0_out[12],magma_UInt_32_mul_inst0_out[11],magma_UInt_32_mul_inst0_out[10],magma_UInt_32_mul_inst0_out[9],magma_UInt_32_mul_inst0_out[8]};
PEGEN_Mux2xBits16 Mux2xBits16_inst19 (
    .I0(Mux2xBits16_inst18_O),
    .I1(Mux2xBits16_inst19_I1),
    .S(magma_Bits_5_eq_inst15_out),
    .O(Mux2xBits16_inst19_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst2 (
    .I0(c),
    .I1(Mux2xBits16_inst1_O),
    .S(Mux2xBit_inst1_O),
    .O(Mux2xBits16_inst2_O)
);
wire [15:0] Mux2xBits16_inst20_I1;
assign Mux2xBits16_inst20_I1 = {magma_UInt_32_mul_inst0_out[15],magma_UInt_32_mul_inst0_out[14],magma_UInt_32_mul_inst0_out[13],magma_UInt_32_mul_inst0_out[12],magma_UInt_32_mul_inst0_out[11],magma_UInt_32_mul_inst0_out[10],magma_UInt_32_mul_inst0_out[9],magma_UInt_32_mul_inst0_out[8],magma_UInt_32_mul_inst0_out[7],magma_UInt_32_mul_inst0_out[6],magma_UInt_32_mul_inst0_out[5],magma_UInt_32_mul_inst0_out[4],magma_UInt_32_mul_inst0_out[3],magma_UInt_32_mul_inst0_out[2],magma_UInt_32_mul_inst0_out[1],magma_UInt_32_mul_inst0_out[0]};
PEGEN_Mux2xBits16 Mux2xBits16_inst20 (
    .I0(Mux2xBits16_inst19_O),
    .I1(Mux2xBits16_inst20_I1),
    .S(magma_Bits_5_eq_inst14_out),
    .O(Mux2xBits16_inst20_O)
);
wire [15:0] Mux2xBits16_inst21_I1;
assign Mux2xBits16_inst21_I1 = {magma_UInt_17_add_inst1_out[15],magma_UInt_17_add_inst1_out[14],magma_UInt_17_add_inst1_out[13],magma_UInt_17_add_inst1_out[12],magma_UInt_17_add_inst1_out[11],magma_UInt_17_add_inst1_out[10],magma_UInt_17_add_inst1_out[9],magma_UInt_17_add_inst1_out[8],magma_UInt_17_add_inst1_out[7],magma_UInt_17_add_inst1_out[6],magma_UInt_17_add_inst1_out[5],magma_UInt_17_add_inst1_out[4],magma_UInt_17_add_inst1_out[3],magma_UInt_17_add_inst1_out[2],magma_UInt_17_add_inst1_out[1],magma_UInt_17_add_inst1_out[0]};
PEGEN_Mux2xBits16 Mux2xBits16_inst21 (
    .I0(Mux2xBits16_inst20_O),
    .I1(Mux2xBits16_inst21_I1),
    .S(magma_Bit_or_inst7_out),
    .O(Mux2xBits16_inst21_O)
);
wire [15:0] Mux2xBits16_inst3_I1;
assign Mux2xBits16_inst3_I1 = {magma_UInt_32_mul_inst0_out[15],magma_UInt_32_mul_inst0_out[14],magma_UInt_32_mul_inst0_out[13],magma_UInt_32_mul_inst0_out[12],magma_UInt_32_mul_inst0_out[11],magma_UInt_32_mul_inst0_out[10],magma_UInt_32_mul_inst0_out[9],magma_UInt_32_mul_inst0_out[8],magma_UInt_32_mul_inst0_out[7],magma_UInt_32_mul_inst0_out[6],magma_UInt_32_mul_inst0_out[5],magma_UInt_32_mul_inst0_out[4],magma_UInt_32_mul_inst0_out[3],magma_UInt_32_mul_inst0_out[2],magma_UInt_32_mul_inst0_out[1],magma_UInt_32_mul_inst0_out[0]};
PEGEN_Mux2xBits16 Mux2xBits16_inst3 (
    .I0(a),
    .I1(Mux2xBits16_inst3_I1),
    .S(magma_Bits_5_eq_inst1_out),
    .O(Mux2xBits16_inst3_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst4 (
    .I0(magma_UInt_16_lshr_inst0_out),
    .I1(magma_SInt_16_ashr_inst0_out),
    .S(magma_Bits_1_eq_inst3_out),
    .O(Mux2xBits16_inst4_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst5 (
    .I0(b),
    .I1(magma_Bits_16_not_inst0_out),
    .S(magma_Bit_or_inst1_out),
    .O(Mux2xBits16_inst5_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst6 (
    .I0(c),
    .I1(magma_Bits_16_not_inst1_out),
    .S(magma_Bit_or_inst6_out),
    .O(Mux2xBits16_inst6_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst7 (
    .I0(magma_SInt_16_neg_inst0_out),
    .I1(a),
    .S(magma_SInt_16_sle_inst1_out),
    .O(Mux2xBits16_inst7_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst8 (
    .I0(Mux2xBits16_inst5_O),
    .I1(a),
    .S(d),
    .O(Mux2xBits16_inst8_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst9 (
    .I0(Mux2xBits16_inst4_O),
    .I1(Mux2xBits16_inst2_O),
    .S(magma_Bits_5_eq_inst30_out),
    .O(Mux2xBits16_inst9_O)
);
wire [15:0] Mux2xUInt16_inst0_I0;
assign Mux2xUInt16_inst0_I0 = {magma_UInt_32_mul_inst0_out[15],magma_UInt_32_mul_inst0_out[14],magma_UInt_32_mul_inst0_out[13],magma_UInt_32_mul_inst0_out[12],magma_UInt_32_mul_inst0_out[11],magma_UInt_32_mul_inst0_out[10],magma_UInt_32_mul_inst0_out[9],magma_UInt_32_mul_inst0_out[8],magma_UInt_32_mul_inst0_out[7],magma_UInt_32_mul_inst0_out[6],magma_UInt_32_mul_inst0_out[5],magma_UInt_32_mul_inst0_out[4],magma_UInt_32_mul_inst0_out[3],magma_UInt_32_mul_inst0_out[2],magma_UInt_32_mul_inst0_out[1],magma_UInt_32_mul_inst0_out[0]};
wire [15:0] Mux2xUInt16_inst0_I1;
assign Mux2xUInt16_inst0_I1 = {magma_UInt_17_add_inst1_out[15],magma_UInt_17_add_inst1_out[14],magma_UInt_17_add_inst1_out[13],magma_UInt_17_add_inst1_out[12],magma_UInt_17_add_inst1_out[11],magma_UInt_17_add_inst1_out[10],magma_UInt_17_add_inst1_out[9],magma_UInt_17_add_inst1_out[8],magma_UInt_17_add_inst1_out[7],magma_UInt_17_add_inst1_out[6],magma_UInt_17_add_inst1_out[5],magma_UInt_17_add_inst1_out[4],magma_UInt_17_add_inst1_out[3],magma_UInt_17_add_inst1_out[2],magma_UInt_17_add_inst1_out[1],magma_UInt_17_add_inst1_out[0]};
PEGEN_Mux2xUInt16 Mux2xUInt16_inst0 (
    .I0(Mux2xUInt16_inst0_I0),
    .I1(Mux2xUInt16_inst0_I1),
    .S(magma_Bit_or_inst4_out),
    .O(Mux2xUInt16_inst0_O)
);
wire [31:0] Mux2xUInt32_inst0_I0;
assign Mux2xUInt32_inst0_I0 = {bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,a};
wire [31:0] Mux2xUInt32_inst0_I1;
assign Mux2xUInt32_inst0_I1 = {a[15],a[15],a[15],a[15],a[15],a[15],a[15],a[15],a[15],a[15],a[15],a[15],a[15],a[15],a[15],a[15],a};
PEGEN_Mux2xUInt32 Mux2xUInt32_inst0 (
    .I0(Mux2xUInt32_inst0_I0),
    .I1(Mux2xUInt32_inst0_I1),
    .S(magma_Bits_1_eq_inst0_out),
    .O(Mux2xUInt32_inst0_O)
);
wire [31:0] Mux2xUInt32_inst1_I0;
assign Mux2xUInt32_inst1_I0 = {bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,b};
wire [31:0] Mux2xUInt32_inst1_I1;
assign Mux2xUInt32_inst1_I1 = {b[15],b[15],b[15],b[15],b[15],b[15],b[15],b[15],b[15],b[15],b[15],b[15],b[15],b[15],b[15],b[15],b};
PEGEN_Mux2xUInt32 Mux2xUInt32_inst1 (
    .I0(Mux2xUInt32_inst1_I0),
    .I1(Mux2xUInt32_inst1_I1),
    .S(magma_Bits_1_eq_inst0_out),
    .O(Mux2xUInt32_inst1_O)
);
PEGEN_corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
PEGEN_corebit_const #(
    .value(1'b1)
) bit_const_1_None (
    .out(bit_const_1_None_out)
);
PEGEN_coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
PEGEN_coreir_const #(
    .value(5'h00),
    .width(5)
) const_0_5 (
    .out(const_0_5_out)
);
PEGEN_coreir_const #(
    .value(5'h0a),
    .width(5)
) const_10_5 (
    .out(const_10_5_out)
);
PEGEN_coreir_const #(
    .value(5'h0b),
    .width(5)
) const_11_5 (
    .out(const_11_5_out)
);
PEGEN_coreir_const #(
    .value(5'h0c),
    .width(5)
) const_12_5 (
    .out(const_12_5_out)
);
PEGEN_coreir_const #(
    .value(5'h0d),
    .width(5)
) const_13_5 (
    .out(const_13_5_out)
);
PEGEN_coreir_const #(
    .value(5'h0e),
    .width(5)
) const_14_5 (
    .out(const_14_5_out)
);
PEGEN_coreir_const #(
    .value(5'h0f),
    .width(5)
) const_15_5 (
    .out(const_15_5_out)
);
PEGEN_coreir_const #(
    .value(5'h10),
    .width(5)
) const_16_5 (
    .out(const_16_5_out)
);
PEGEN_coreir_const #(
    .value(5'h11),
    .width(5)
) const_17_5 (
    .out(const_17_5_out)
);
PEGEN_coreir_const #(
    .value(5'h12),
    .width(5)
) const_18_5 (
    .out(const_18_5_out)
);
PEGEN_coreir_const #(
    .value(5'h13),
    .width(5)
) const_19_5 (
    .out(const_19_5_out)
);
PEGEN_coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
PEGEN_coreir_const #(
    .value(5'h01),
    .width(5)
) const_1_5 (
    .out(const_1_5_out)
);
PEGEN_coreir_const #(
    .value(5'h02),
    .width(5)
) const_2_5 (
    .out(const_2_5_out)
);
PEGEN_coreir_const #(
    .value(5'h03),
    .width(5)
) const_3_5 (
    .out(const_3_5_out)
);
PEGEN_coreir_const #(
    .value(5'h04),
    .width(5)
) const_4_5 (
    .out(const_4_5_out)
);
PEGEN_coreir_const #(
    .value(5'h05),
    .width(5)
) const_5_5 (
    .out(const_5_5_out)
);
PEGEN_coreir_const #(
    .value(5'h06),
    .width(5)
) const_6_5 (
    .out(const_6_5_out)
);
PEGEN_coreir_const #(
    .value(5'h07),
    .width(5)
) const_7_5 (
    .out(const_7_5_out)
);
PEGEN_coreir_const #(
    .value(5'h08),
    .width(5)
) const_8_5 (
    .out(const_8_5_out)
);
PEGEN_coreir_const #(
    .value(5'h09),
    .width(5)
) const_9_5 (
    .out(const_9_5_out)
);
PEGEN_corebit_and magma_Bit_and_inst0 (
    .in0(a[15]),
    .in1(Mux2xBits16_inst5_O[15]),
    .out(magma_Bit_and_inst0_out)
);
PEGEN_corebit_and magma_Bit_and_inst1 (
    .in0(magma_Bit_and_inst0_out),
    .in1(magma_Bit_not_inst0_out),
    .out(magma_Bit_and_inst1_out)
);
PEGEN_corebit_and magma_Bit_and_inst2 (
    .in0(magma_Bit_not_inst1_out),
    .in1(magma_Bit_not_inst2_out),
    .out(magma_Bit_and_inst2_out)
);
PEGEN_corebit_and magma_Bit_and_inst3 (
    .in0(magma_Bit_and_inst2_out),
    .in1(magma_UInt_17_add_inst1_out[15]),
    .out(magma_Bit_and_inst3_out)
);
PEGEN_corebit_not magma_Bit_not_inst0 (
    .in(magma_UInt_17_add_inst1_out[15]),
    .out(magma_Bit_not_inst0_out)
);
PEGEN_corebit_not magma_Bit_not_inst1 (
    .in(a[15]),
    .out(magma_Bit_not_inst1_out)
);
PEGEN_corebit_not magma_Bit_not_inst2 (
    .in(Mux2xBits16_inst5_O[15]),
    .out(magma_Bit_not_inst2_out)
);
PEGEN_corebit_or magma_Bit_or_inst0 (
    .in0(magma_Bits_5_eq_inst2_out),
    .in1(magma_Bits_5_eq_inst3_out),
    .out(magma_Bit_or_inst0_out)
);
PEGEN_corebit_or magma_Bit_or_inst1 (
    .in0(magma_Bit_or_inst0_out),
    .in1(magma_Bits_5_eq_inst4_out),
    .out(magma_Bit_or_inst1_out)
);
PEGEN_corebit_or magma_Bit_or_inst10 (
    .in0(magma_Bit_or_inst9_out),
    .in1(magma_Bits_5_eq_inst26_out),
    .out(magma_Bit_or_inst10_out)
);
PEGEN_corebit_or magma_Bit_or_inst11 (
    .in0(magma_Bit_or_inst10_out),
    .in1(magma_Bits_5_eq_inst27_out),
    .out(magma_Bit_or_inst11_out)
);
PEGEN_corebit_or magma_Bit_or_inst12 (
    .in0(magma_Bit_or_inst11_out),
    .in1(magma_Bits_5_eq_inst28_out),
    .out(magma_Bit_or_inst12_out)
);
PEGEN_corebit_or magma_Bit_or_inst13 (
    .in0(magma_Bit_or_inst12_out),
    .in1(magma_Bits_5_eq_inst29_out),
    .out(magma_Bit_or_inst13_out)
);
PEGEN_corebit_or magma_Bit_or_inst2 (
    .in0(magma_Bits_5_eq_inst5_out),
    .in1(magma_Bits_5_eq_inst6_out),
    .out(magma_Bit_or_inst2_out)
);
PEGEN_corebit_or magma_Bit_or_inst3 (
    .in0(magma_Bit_or_inst2_out),
    .in1(magma_Bits_5_eq_inst7_out),
    .out(magma_Bit_or_inst3_out)
);
PEGEN_corebit_or magma_Bit_or_inst4 (
    .in0(magma_Bit_or_inst3_out),
    .in1(magma_Bits_5_eq_inst8_out),
    .out(magma_Bit_or_inst4_out)
);
PEGEN_corebit_or magma_Bit_or_inst5 (
    .in0(magma_Bits_5_eq_inst9_out),
    .in1(magma_Bits_5_eq_inst10_out),
    .out(magma_Bit_or_inst5_out)
);
PEGEN_corebit_or magma_Bit_or_inst6 (
    .in0(magma_Bit_or_inst5_out),
    .in1(magma_Bits_5_eq_inst11_out),
    .out(magma_Bit_or_inst6_out)
);
PEGEN_corebit_or magma_Bit_or_inst7 (
    .in0(magma_Bits_5_eq_inst12_out),
    .in1(magma_Bits_5_eq_inst13_out),
    .out(magma_Bit_or_inst7_out)
);
PEGEN_corebit_or magma_Bit_or_inst8 (
    .in0(magma_Bit_and_inst1_out),
    .in1(magma_Bit_and_inst3_out),
    .out(magma_Bit_or_inst8_out)
);
PEGEN_corebit_or magma_Bit_or_inst9 (
    .in0(magma_Bits_5_eq_inst24_out),
    .in1(magma_Bits_5_eq_inst25_out),
    .out(magma_Bit_or_inst9_out)
);
PEGEN_coreir_and #(
    .width(16)
) magma_Bits_16_and_inst0 (
    .in0(a),
    .in1(Mux2xBits16_inst5_O),
    .out(magma_Bits_16_and_inst0_out)
);
PEGEN_coreir_not #(
    .width(16)
) magma_Bits_16_not_inst0 (
    .in(b),
    .out(magma_Bits_16_not_inst0_out)
);
PEGEN_coreir_not #(
    .width(16)
) magma_Bits_16_not_inst1 (
    .in(c),
    .out(magma_Bits_16_not_inst1_out)
);
PEGEN_coreir_or #(
    .width(16)
) magma_Bits_16_or_inst0 (
    .in0(a),
    .in1(Mux2xBits16_inst5_O),
    .out(magma_Bits_16_or_inst0_out)
);
PEGEN_coreir_shl #(
    .width(16)
) magma_Bits_16_shl_inst0 (
    .in0(a),
    .in1(Mux2xBits16_inst5_O),
    .out(magma_Bits_16_shl_inst0_out)
);
PEGEN_coreir_xor #(
    .width(16)
) magma_Bits_16_xor_inst0 (
    .in0(a),
    .in1(Mux2xBits16_inst5_O),
    .out(magma_Bits_16_xor_inst0_out)
);
PEGEN_coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst0 (
    .in0(signed_),
    .in1(const_1_1_out),
    .out(magma_Bits_1_eq_inst0_out)
);
PEGEN_coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst1 (
    .in0(signed_),
    .in1(const_1_1_out),
    .out(magma_Bits_1_eq_inst1_out)
);
PEGEN_coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst2 (
    .in0(signed_),
    .in1(const_1_1_out),
    .out(magma_Bits_1_eq_inst2_out)
);
PEGEN_coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst3 (
    .in0(signed_),
    .in1(const_1_1_out),
    .out(magma_Bits_1_eq_inst3_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst0 (
    .in0(alu),
    .in1(const_18_5_out),
    .out(magma_Bits_5_eq_inst0_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst1 (
    .in0(alu),
    .in1(const_19_5_out),
    .out(magma_Bits_5_eq_inst1_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst10 (
    .in0(alu),
    .in1(const_15_5_out),
    .out(magma_Bits_5_eq_inst10_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst11 (
    .in0(alu),
    .in1(const_17_5_out),
    .out(magma_Bits_5_eq_inst11_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst12 (
    .in0(alu),
    .in1(const_0_5_out),
    .out(magma_Bits_5_eq_inst12_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst13 (
    .in0(alu),
    .in1(const_1_5_out),
    .out(magma_Bits_5_eq_inst13_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst14 (
    .in0(alu),
    .in1(const_4_5_out),
    .out(magma_Bits_5_eq_inst14_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst15 (
    .in0(alu),
    .in1(const_5_5_out),
    .out(magma_Bits_5_eq_inst15_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst16 (
    .in0(alu),
    .in1(const_6_5_out),
    .out(magma_Bits_5_eq_inst16_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst17 (
    .in0(alu),
    .in1(const_2_5_out),
    .out(magma_Bits_5_eq_inst17_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst18 (
    .in0(alu),
    .in1(const_3_5_out),
    .out(magma_Bits_5_eq_inst18_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst19 (
    .in0(alu),
    .in1(const_10_5_out),
    .out(magma_Bits_5_eq_inst19_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst2 (
    .in0(alu),
    .in1(const_1_5_out),
    .out(magma_Bits_5_eq_inst2_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst20 (
    .in0(alu),
    .in1(const_9_5_out),
    .out(magma_Bits_5_eq_inst20_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst21 (
    .in0(alu),
    .in1(const_11_5_out),
    .out(magma_Bits_5_eq_inst21_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst22 (
    .in0(alu),
    .in1(const_7_5_out),
    .out(magma_Bits_5_eq_inst22_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst23 (
    .in0(alu),
    .in1(const_8_5_out),
    .out(magma_Bits_5_eq_inst23_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst24 (
    .in0(alu),
    .in1(const_12_5_out),
    .out(magma_Bits_5_eq_inst24_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst25 (
    .in0(alu),
    .in1(const_13_5_out),
    .out(magma_Bits_5_eq_inst25_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst26 (
    .in0(alu),
    .in1(const_14_5_out),
    .out(magma_Bits_5_eq_inst26_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst27 (
    .in0(alu),
    .in1(const_16_5_out),
    .out(magma_Bits_5_eq_inst27_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst28 (
    .in0(alu),
    .in1(const_15_5_out),
    .out(magma_Bits_5_eq_inst28_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst29 (
    .in0(alu),
    .in1(const_17_5_out),
    .out(magma_Bits_5_eq_inst29_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst3 (
    .in0(alu),
    .in1(const_16_5_out),
    .out(magma_Bits_5_eq_inst3_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst30 (
    .in0(alu),
    .in1(const_18_5_out),
    .out(magma_Bits_5_eq_inst30_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst4 (
    .in0(alu),
    .in1(const_17_5_out),
    .out(magma_Bits_5_eq_inst4_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst5 (
    .in0(alu),
    .in1(const_14_5_out),
    .out(magma_Bits_5_eq_inst5_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst6 (
    .in0(alu),
    .in1(const_15_5_out),
    .out(magma_Bits_5_eq_inst6_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst7 (
    .in0(alu),
    .in1(const_16_5_out),
    .out(magma_Bits_5_eq_inst7_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst8 (
    .in0(alu),
    .in1(const_17_5_out),
    .out(magma_Bits_5_eq_inst8_out)
);
PEGEN_coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst9 (
    .in0(alu),
    .in1(const_13_5_out),
    .out(magma_Bits_5_eq_inst9_out)
);
PEGEN_coreir_ashr #(
    .width(16)
) magma_SInt_16_ashr_inst0 (
    .in0(Mux2xBits16_inst3_O),
    .in1(c),
    .out(magma_SInt_16_ashr_inst0_out)
);
PEGEN_coreir_eq #(
    .width(16)
) magma_SInt_16_eq_inst0 (
    .in0(const_0_16_out),
    .in1(Mux2xBits16_inst21_O),
    .out(magma_SInt_16_eq_inst0_out)
);
PEGEN_coreir_neg #(
    .width(16)
) magma_SInt_16_neg_inst0 (
    .in(a),
    .out(magma_SInt_16_neg_inst0_out)
);
PEGEN_coreir_sge #(
    .width(16)
) magma_SInt_16_sge_inst0 (
    .in0(Mux2xBits16_inst1_O),
    .in1(c),
    .out(magma_SInt_16_sge_inst0_out)
);
PEGEN_coreir_sle #(
    .width(16)
) magma_SInt_16_sle_inst0 (
    .in0(a),
    .in1(b),
    .out(magma_SInt_16_sle_inst0_out)
);
PEGEN_coreir_sle #(
    .width(16)
) magma_SInt_16_sle_inst1 (
    .in0(const_0_16_out),
    .in1(a),
    .out(magma_SInt_16_sle_inst1_out)
);
PEGEN_coreir_lshr #(
    .width(16)
) magma_UInt_16_lshr_inst0 (
    .in0(Mux2xBits16_inst3_O),
    .in1(c),
    .out(magma_UInt_16_lshr_inst0_out)
);
PEGEN_coreir_uge #(
    .width(16)
) magma_UInt_16_uge_inst0 (
    .in0(Mux2xBits16_inst1_O),
    .in1(c),
    .out(magma_UInt_16_uge_inst0_out)
);
PEGEN_coreir_ule #(
    .width(16)
) magma_UInt_16_ule_inst0 (
    .in0(a),
    .in1(b),
    .out(magma_UInt_16_ule_inst0_out)
);
wire [16:0] magma_UInt_17_add_inst0_in0;
assign magma_UInt_17_add_inst0_in0 = {bit_const_0_None_out,a};
wire [16:0] magma_UInt_17_add_inst0_in1;
assign magma_UInt_17_add_inst0_in1 = {bit_const_0_None_out,Mux2xBits16_inst5_O};
PEGEN_coreir_add #(
    .width(17)
) magma_UInt_17_add_inst0 (
    .in0(magma_UInt_17_add_inst0_in0),
    .in1(magma_UInt_17_add_inst0_in1),
    .out(magma_UInt_17_add_inst0_out)
);
wire [16:0] magma_UInt_17_add_inst1_in1;
assign magma_UInt_17_add_inst1_in1 = {bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,d};
PEGEN_coreir_add #(
    .width(17)
) magma_UInt_17_add_inst1 (
    .in0(magma_UInt_17_add_inst0_out),
    .in1(magma_UInt_17_add_inst1_in1),
    .out(magma_UInt_17_add_inst1_out)
);
wire [16:0] magma_UInt_17_add_inst2_in0;
assign magma_UInt_17_add_inst2_in0 = {bit_const_0_None_out,Mux2xUInt16_inst0_O};
wire [16:0] magma_UInt_17_add_inst2_in1;
assign magma_UInt_17_add_inst2_in1 = {bit_const_0_None_out,Mux2xBits16_inst6_O};
PEGEN_coreir_add #(
    .width(17)
) magma_UInt_17_add_inst2 (
    .in0(magma_UInt_17_add_inst2_in0),
    .in1(magma_UInt_17_add_inst2_in1),
    .out(magma_UInt_17_add_inst2_out)
);
wire [16:0] magma_UInt_17_add_inst3_in1;
assign magma_UInt_17_add_inst3_in1 = {bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,Mux2xBit_inst2_O};
PEGEN_coreir_add #(
    .width(17)
) magma_UInt_17_add_inst3 (
    .in0(magma_UInt_17_add_inst2_out),
    .in1(magma_UInt_17_add_inst3_in1),
    .out(magma_UInt_17_add_inst3_out)
);
PEGEN_coreir_mul #(
    .width(32)
) magma_UInt_32_mul_inst0 (
    .in0(Mux2xUInt32_inst0_O),
    .in1(Mux2xUInt32_inst1_O),
    .out(magma_UInt_32_mul_inst0_out)
);
assign res = Mux2xBits16_inst21_O;
assign res_p = Mux2xBit_inst23_O;
assign Z = magma_SInt_16_eq_inst0_out;
assign N = Mux2xBits16_inst21_O[15];
assign C = Mux2xBit_inst21_O;
assign V = Mux2xBit_inst22_O;
endmodule

module PEGEN_PE (
    input [83:0] inst,
    input [15:0] data0,
    input [15:0] data1,
    input [15:0] data2,
    input bit0,
    input bit1,
    input bit2,
    input clk_en,
    output [15:0] O0,
    output O1,
    output [15:0] O2,
    output [15:0] O3,
    output [15:0] O4,
    input CLK,
    input ASYNCRESET
);
wire [15:0] ALU_inst0_res;
wire ALU_inst0_res_p;
wire ALU_inst0_Z;
wire ALU_inst0_N;
wire ALU_inst0_C;
wire ALU_inst0_V;
wire Cond_inst0_O;
wire LUT_inst0_O;
wire Mux2xBit_inst0_O;
wire Mux2xBit_inst1_O;
wire Mux2xBit_inst2_O;
wire Mux2xBit_inst3_O;
wire [15:0] Mux2xBits16_inst0_O;
wire [4:0] Mux2xMagmaADTALU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_O;
wire [15:0] RegisterMode_inst0_O0;
wire [15:0] RegisterMode_inst0_O1;
wire [15:0] RegisterMode_inst1_O0;
wire [15:0] RegisterMode_inst1_O1;
wire [15:0] RegisterMode_inst2_O0;
wire [15:0] RegisterMode_inst2_O1;
wire RegisterMode_inst3_O0;
wire RegisterMode_inst3_O1;
wire RegisterMode_inst4_O0;
wire RegisterMode_inst4_O1;
wire RegisterMode_inst5_O0;
wire RegisterMode_inst5_O1;
wire bit_const_0_None_out;
wire [15:0] const_0_16_out;
wire [1:0] const_0_2_out;
wire [4:0] const_0_5_out;
wire magma_Bits_2_eq_inst0_out;
wire magma_Bits_2_eq_inst1_out;
wire magma_Bits_2_eq_inst2_out;
PEGEN_ALU ALU_inst0 (
    .alu(Mux2xMagmaADTALU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_O),
    .signed_(inst[7:7]),
    .a(RegisterMode_inst0_O0),
    .b(RegisterMode_inst1_O0),
    .c(RegisterMode_inst2_O0),
    .d(RegisterMode_inst3_O0),
    .res(ALU_inst0_res),
    .res_p(ALU_inst0_res_p),
    .Z(ALU_inst0_Z),
    .N(ALU_inst0_N),
    .C(ALU_inst0_C),
    .V(ALU_inst0_V),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
PEGEN_Cond Cond_inst0 (
    .code(inst[20:16]),
    .alu(Mux2xBit_inst3_O),
    .lut(LUT_inst0_O),
    .Z(Mux2xBit_inst2_O),
    .N(Mux2xBit_inst0_O),
    .C(ALU_inst0_C),
    .V(Mux2xBit_inst1_O),
    .O(Cond_inst0_O),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
wire [7:0] LUT_inst0_lut;
assign LUT_inst0_lut = {inst[15],inst[14],inst[13],inst[12],inst[11],inst[10],inst[9],inst[8]};
PEGEN_LUT LUT_inst0 (
    .lut(LUT_inst0_lut),
    .bit0(RegisterMode_inst3_O0),
    .bit1(RegisterMode_inst4_O0),
    .bit2(RegisterMode_inst5_O0),
    .O(LUT_inst0_O),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
PEGEN_Mux2xBit Mux2xBit_inst0 (
    .I0(bit_const_0_None_out),
    .I1(ALU_inst0_N),
    .S(magma_Bits_2_eq_inst2_out),
    .O(Mux2xBit_inst0_O)
);
PEGEN_Mux2xBit Mux2xBit_inst1 (
    .I0(bit_const_0_None_out),
    .I1(ALU_inst0_V),
    .S(magma_Bits_2_eq_inst2_out),
    .O(Mux2xBit_inst1_O)
);
PEGEN_Mux2xBit Mux2xBit_inst2 (
    .I0(bit_const_0_None_out),
    .I1(ALU_inst0_Z),
    .S(magma_Bits_2_eq_inst2_out),
    .O(Mux2xBit_inst2_O)
);
PEGEN_Mux2xBit Mux2xBit_inst3 (
    .I0(bit_const_0_None_out),
    .I1(ALU_inst0_res_p),
    .S(magma_Bits_2_eq_inst2_out),
    .O(Mux2xBit_inst3_O)
);
PEGEN_Mux2xBits16 Mux2xBits16_inst0 (
    .I0(const_0_16_out),
    .I1(ALU_inst0_res),
    .S(magma_Bits_2_eq_inst2_out),
    .O(Mux2xBits16_inst0_O)
);
wire [4:0] Mux2xMagmaADTALU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_I1;
assign Mux2xMagmaADTALU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_I1 = {inst[6],inst[5],inst[4],inst[3],inst[2]};
PEGEN_Mux2xMagmaADTALU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3 Mux2xMagmaADTALU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0 (
    .I0(const_0_5_out),
    .I1(Mux2xMagmaADTALU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_I1),
    .S(magma_Bits_2_eq_inst0_out),
    .O(Mux2xMagmaADTALU_t_classpeakassemblerassemblerAssembler_Bits_DirectionUndirected3_inst0_O)
);
wire [15:0] RegisterMode_inst0_const_;
assign RegisterMode_inst0_const_ = {inst[38],inst[37],inst[36],inst[35],inst[34],inst[33],inst[32],inst[31],inst[30],inst[29],inst[28],inst[27],inst[26],inst[25],inst[24],inst[23]};
PEGEN_RegisterMode RegisterMode_inst0 (
    .mode(inst[22:21]),
    .const_(RegisterMode_inst0_const_),
    .value(data0),
    .clk_en(clk_en),
    .O0(RegisterMode_inst0_O0),
    .O1(RegisterMode_inst0_O1),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
wire [15:0] RegisterMode_inst1_const_;
assign RegisterMode_inst1_const_ = {inst[56],inst[55],inst[54],inst[53],inst[52],inst[51],inst[50],inst[49],inst[48],inst[47],inst[46],inst[45],inst[44],inst[43],inst[42],inst[41]};
PEGEN_RegisterMode RegisterMode_inst1 (
    .mode(inst[40:39]),
    .const_(RegisterMode_inst1_const_),
    .value(data1),
    .clk_en(clk_en),
    .O0(RegisterMode_inst1_O0),
    .O1(RegisterMode_inst1_O1),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
wire [15:0] RegisterMode_inst2_const_;
assign RegisterMode_inst2_const_ = {inst[74],inst[73],inst[72],inst[71],inst[70],inst[69],inst[68],inst[67],inst[66],inst[65],inst[64],inst[63],inst[62],inst[61],inst[60],inst[59]};
PEGEN_RegisterMode RegisterMode_inst2 (
    .mode(inst[58:57]),
    .const_(RegisterMode_inst2_const_),
    .value(data2),
    .clk_en(clk_en),
    .O0(RegisterMode_inst2_O0),
    .O1(RegisterMode_inst2_O1),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
PEGEN_RegisterMode_unq1 RegisterMode_inst3 (
    .mode(inst[76:75]),
    .const_(inst[77]),
    .value(bit0),
    .clk_en(clk_en),
    .O0(RegisterMode_inst3_O0),
    .O1(RegisterMode_inst3_O1),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
PEGEN_RegisterMode_unq1 RegisterMode_inst4 (
    .mode(inst[79:78]),
    .const_(inst[80]),
    .value(bit1),
    .clk_en(clk_en),
    .O0(RegisterMode_inst4_O0),
    .O1(RegisterMode_inst4_O1),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
PEGEN_RegisterMode_unq1 RegisterMode_inst5 (
    .mode(inst[82:81]),
    .const_(inst[83]),
    .value(bit2),
    .clk_en(clk_en),
    .O0(RegisterMode_inst5_O0),
    .O1(RegisterMode_inst5_O1),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
PEGEN_corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
PEGEN_coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
PEGEN_coreir_const #(
    .value(2'h0),
    .width(2)
) const_0_2 (
    .out(const_0_2_out)
);
PEGEN_coreir_const #(
    .value(5'h00),
    .width(5)
) const_0_5 (
    .out(const_0_5_out)
);
wire [1:0] magma_Bits_2_eq_inst0_in0;
assign magma_Bits_2_eq_inst0_in0 = {inst[1],inst[0]};
PEGEN_coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst0 (
    .in0(magma_Bits_2_eq_inst0_in0),
    .in1(const_0_2_out),
    .out(magma_Bits_2_eq_inst0_out)
);
wire [1:0] magma_Bits_2_eq_inst1_in0;
assign magma_Bits_2_eq_inst1_in0 = {inst[1],inst[0]};
PEGEN_coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst1 (
    .in0(magma_Bits_2_eq_inst1_in0),
    .in1(const_0_2_out),
    .out(magma_Bits_2_eq_inst1_out)
);
wire [1:0] magma_Bits_2_eq_inst2_in0;
assign magma_Bits_2_eq_inst2_in0 = {inst[1],inst[0]};
PEGEN_coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst2 (
    .in0(magma_Bits_2_eq_inst2_in0),
    .in1(const_0_2_out),
    .out(magma_Bits_2_eq_inst2_out)
);
assign O0 = Mux2xBits16_inst0_O;
assign O1 = Cond_inst0_O;
assign O2 = RegisterMode_inst0_O1;
assign O3 = RegisterMode_inst1_O1;
assign O4 = RegisterMode_inst2_O1;
endmodule

